// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689
`timescale 1ns / 1ps

module out_axis_args #(
    parameter C_NUM_OUTPUT_AXISs = 0,
    parameter [31:0] M_AXIS_OARG_0_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_1_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_2_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_3_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_4_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_5_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_6_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_7_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_8_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_9_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_10_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_11_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_12_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_13_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_14_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_15_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_16_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_17_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_18_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_19_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_20_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_21_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_22_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_23_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_24_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_25_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_26_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_27_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_28_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_29_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_30_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_31_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_32_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_33_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_34_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_35_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_36_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_37_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_38_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_39_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_40_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_41_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_42_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_43_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_44_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_45_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_46_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_47_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_48_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_49_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_50_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_51_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_52_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_53_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_54_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_55_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_56_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_57_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_58_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_59_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_60_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_61_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_62_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_63_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_64_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_65_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_66_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_67_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_68_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_69_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_70_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_71_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_72_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_73_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_74_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_75_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_76_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_77_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_78_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_79_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_80_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_81_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_82_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_83_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_84_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_85_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_86_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_87_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_88_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_89_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_90_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_91_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_92_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_93_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_94_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_95_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_96_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_97_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_98_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_99_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_100_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_101_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_102_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_103_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_104_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_105_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_106_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_107_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_108_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_109_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_110_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_111_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_112_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_113_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_114_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_115_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_116_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_117_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_118_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_119_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_120_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_121_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_122_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_123_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_124_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_125_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_126_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_127_WIDTH = 8,    //width of output axis interface on the accelerator
    parameter [31:0] M_AXIS_OARG_0_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_1_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_2_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_3_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_4_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_5_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_6_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_7_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_8_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_9_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_10_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_11_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_12_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_13_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_14_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_15_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_16_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_17_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_18_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_19_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_20_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_21_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_22_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_23_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_24_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_25_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_26_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_27_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_28_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_29_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_30_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_31_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_32_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_33_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_34_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_35_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_36_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_37_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_38_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_39_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_40_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_41_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_42_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_43_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_44_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_45_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_46_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_47_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_48_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_49_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_50_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_51_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_52_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_53_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_54_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_55_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_56_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_57_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_58_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_59_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_60_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_61_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_62_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_63_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_64_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_65_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_66_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_67_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_68_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_69_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_70_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_71_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_72_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_73_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_74_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_75_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_76_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_77_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_78_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_79_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_80_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_81_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_82_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_83_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_84_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_85_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_86_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_87_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_88_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_89_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_90_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_91_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_92_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_93_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_94_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_95_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_96_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_97_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_98_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_99_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_100_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_101_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_102_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_103_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_104_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_105_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_106_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_107_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_108_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_109_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_110_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_111_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_112_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_113_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_114_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_115_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_116_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_117_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_118_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_119_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_120_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_121_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_122_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_123_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_124_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_125_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_126_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_127_DEPTH = 16,     //depth of FIFO in adapter for output axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_0_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_1_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_2_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_3_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_4_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_5_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_6_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_7_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_8_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_9_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_10_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_11_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_12_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_13_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_14_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_15_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_16_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_17_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_18_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_19_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_20_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_21_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_22_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_23_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_24_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_25_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_26_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_27_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_28_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_29_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_30_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_31_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_32_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_33_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_34_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_35_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_36_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_37_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_38_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_39_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_40_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_41_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_42_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_43_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_44_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_45_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_46_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_47_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_48_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_49_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_50_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_51_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_52_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_53_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_54_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_55_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_56_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_57_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_58_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_59_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_60_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_61_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_62_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_63_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_64_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_65_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_66_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_67_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_68_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_69_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_70_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_71_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_72_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_73_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_74_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_75_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_76_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_77_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_78_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_79_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_80_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_81_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_82_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_83_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_84_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_85_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_86_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_87_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_88_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_89_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_90_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_91_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_92_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_93_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_94_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_95_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_96_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_97_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_98_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_99_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_100_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_101_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_102_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_103_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_104_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_105_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_106_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_107_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_108_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_109_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_110_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_111_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_112_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_113_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_114_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_115_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_116_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_117_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_118_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_119_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_120_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_121_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_122_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_123_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_124_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_125_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_126_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_127_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output axis interface
    parameter [31:0] M_AXIS_OARG_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_0_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_1_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_2_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_3_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_4_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_5_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_6_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_7_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_8_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_9_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_10_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_11_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_12_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_13_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_14_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_15_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_16_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_17_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_18_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_19_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_20_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_21_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_22_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_23_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_24_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_25_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_26_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_27_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_28_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_29_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_30_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_31_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_32_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_33_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_34_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_35_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_36_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_37_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_38_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_39_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_40_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_41_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_42_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_43_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_44_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_45_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_46_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_47_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_48_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_49_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_50_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_51_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_52_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_53_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_54_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_55_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_56_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_57_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_58_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_59_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_60_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_61_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_62_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_63_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_64_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_65_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_66_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_67_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_68_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_69_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_70_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_71_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_72_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_73_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_74_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_75_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_76_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_77_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_78_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_79_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_80_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_81_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_82_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_83_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_84_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_85_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_86_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_87_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_88_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_89_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_90_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_91_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_92_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_93_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_94_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_95_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_96_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_97_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_98_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_99_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_100_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_101_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_102_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_103_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_104_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_105_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_106_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_107_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_108_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_109_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_110_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_111_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_112_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_113_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_114_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_115_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_116_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_117_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_118_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_119_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_120_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_121_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_122_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_123_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_124_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_125_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_126_GEN_TLAST = 0,  //generate TLAST signal
    parameter [31:0] M_AXIS_OARG_127_GEN_TLAST = 0  //generate TLAST signal
 ) (
    input acc_clk,
    input acc_aresetn,
    //control interface
    input out_axis_allow,
    output [C_NUM_OUTPUT_AXISs-1:0] out_axis_ready,
    output [C_NUM_OUTPUT_AXISs-1:0] out_axis_finished,
    //output AXIS to AXI-Stream interface 0
    input m_axis_oarg_0_aclk,
    input m_axis_oarg_0_aresetn,
    output m_axis_oarg_0_tlast,
    output m_axis_oarg_0_tvalid,
    output [M_AXIS_OARG_0_DMWIDTH/8-1:0] m_axis_oarg_0_tkeep,
    output [M_AXIS_OARG_0_DMWIDTH/8-1:0] m_axis_oarg_0_tstrb,
    output [M_AXIS_OARG_0_DMWIDTH-1:0] m_axis_oarg_0_tdata,
    input m_axis_oarg_0_tready,
    input ap_axis_oarg_0_tlast,
    input ap_axis_oarg_0_tvalid,
    input [M_AXIS_OARG_0_WIDTH/8-1:0] ap_axis_oarg_0_tkeep,
    input [M_AXIS_OARG_0_WIDTH/8-1:0] ap_axis_oarg_0_tstrb,
    input [M_AXIS_OARG_0_WIDTH-1:0] ap_axis_oarg_0_tdata,
    output ap_axis_oarg_0_tready,
    //output AXIS to AXI-Stream interface 1
    input m_axis_oarg_1_aclk,
    input m_axis_oarg_1_aresetn,
    output m_axis_oarg_1_tlast,
    output m_axis_oarg_1_tvalid,
    output [M_AXIS_OARG_1_DMWIDTH/8-1:0] m_axis_oarg_1_tkeep,
    output [M_AXIS_OARG_1_DMWIDTH/8-1:0] m_axis_oarg_1_tstrb,
    output [M_AXIS_OARG_1_DMWIDTH-1:0] m_axis_oarg_1_tdata,
    input m_axis_oarg_1_tready,
    input ap_axis_oarg_1_tlast,
    input ap_axis_oarg_1_tvalid,
    input [M_AXIS_OARG_1_WIDTH/8-1:0] ap_axis_oarg_1_tkeep,
    input [M_AXIS_OARG_1_WIDTH/8-1:0] ap_axis_oarg_1_tstrb,
    input [M_AXIS_OARG_1_WIDTH-1:0] ap_axis_oarg_1_tdata,
    output ap_axis_oarg_1_tready,
    //output AXIS to AXI-Stream interface 2
    input m_axis_oarg_2_aclk,
    input m_axis_oarg_2_aresetn,
    output m_axis_oarg_2_tlast,
    output m_axis_oarg_2_tvalid,
    output [M_AXIS_OARG_2_DMWIDTH/8-1:0] m_axis_oarg_2_tkeep,
    output [M_AXIS_OARG_2_DMWIDTH/8-1:0] m_axis_oarg_2_tstrb,
    output [M_AXIS_OARG_2_DMWIDTH-1:0] m_axis_oarg_2_tdata,
    input m_axis_oarg_2_tready,
    input ap_axis_oarg_2_tlast,
    input ap_axis_oarg_2_tvalid,
    input [M_AXIS_OARG_2_WIDTH/8-1:0] ap_axis_oarg_2_tkeep,
    input [M_AXIS_OARG_2_WIDTH/8-1:0] ap_axis_oarg_2_tstrb,
    input [M_AXIS_OARG_2_WIDTH-1:0] ap_axis_oarg_2_tdata,
    output ap_axis_oarg_2_tready,
    //output AXIS to AXI-Stream interface 3
    input m_axis_oarg_3_aclk,
    input m_axis_oarg_3_aresetn,
    output m_axis_oarg_3_tlast,
    output m_axis_oarg_3_tvalid,
    output [M_AXIS_OARG_3_DMWIDTH/8-1:0] m_axis_oarg_3_tkeep,
    output [M_AXIS_OARG_3_DMWIDTH/8-1:0] m_axis_oarg_3_tstrb,
    output [M_AXIS_OARG_3_DMWIDTH-1:0] m_axis_oarg_3_tdata,
    input m_axis_oarg_3_tready,
    input ap_axis_oarg_3_tlast,
    input ap_axis_oarg_3_tvalid,
    input [M_AXIS_OARG_3_WIDTH/8-1:0] ap_axis_oarg_3_tkeep,
    input [M_AXIS_OARG_3_WIDTH/8-1:0] ap_axis_oarg_3_tstrb,
    input [M_AXIS_OARG_3_WIDTH-1:0] ap_axis_oarg_3_tdata,
    output ap_axis_oarg_3_tready,
    //output AXIS to AXI-Stream interface 4
    input m_axis_oarg_4_aclk,
    input m_axis_oarg_4_aresetn,
    output m_axis_oarg_4_tlast,
    output m_axis_oarg_4_tvalid,
    output [M_AXIS_OARG_4_DMWIDTH/8-1:0] m_axis_oarg_4_tkeep,
    output [M_AXIS_OARG_4_DMWIDTH/8-1:0] m_axis_oarg_4_tstrb,
    output [M_AXIS_OARG_4_DMWIDTH-1:0] m_axis_oarg_4_tdata,
    input m_axis_oarg_4_tready,
    input ap_axis_oarg_4_tlast,
    input ap_axis_oarg_4_tvalid,
    input [M_AXIS_OARG_4_WIDTH/8-1:0] ap_axis_oarg_4_tkeep,
    input [M_AXIS_OARG_4_WIDTH/8-1:0] ap_axis_oarg_4_tstrb,
    input [M_AXIS_OARG_4_WIDTH-1:0] ap_axis_oarg_4_tdata,
    output ap_axis_oarg_4_tready,
    //output AXIS to AXI-Stream interface 5
    input m_axis_oarg_5_aclk,
    input m_axis_oarg_5_aresetn,
    output m_axis_oarg_5_tlast,
    output m_axis_oarg_5_tvalid,
    output [M_AXIS_OARG_5_DMWIDTH/8-1:0] m_axis_oarg_5_tkeep,
    output [M_AXIS_OARG_5_DMWIDTH/8-1:0] m_axis_oarg_5_tstrb,
    output [M_AXIS_OARG_5_DMWIDTH-1:0] m_axis_oarg_5_tdata,
    input m_axis_oarg_5_tready,
    input ap_axis_oarg_5_tlast,
    input ap_axis_oarg_5_tvalid,
    input [M_AXIS_OARG_5_WIDTH/8-1:0] ap_axis_oarg_5_tkeep,
    input [M_AXIS_OARG_5_WIDTH/8-1:0] ap_axis_oarg_5_tstrb,
    input [M_AXIS_OARG_5_WIDTH-1:0] ap_axis_oarg_5_tdata,
    output ap_axis_oarg_5_tready,
    //output AXIS to AXI-Stream interface 6
    input m_axis_oarg_6_aclk,
    input m_axis_oarg_6_aresetn,
    output m_axis_oarg_6_tlast,
    output m_axis_oarg_6_tvalid,
    output [M_AXIS_OARG_6_DMWIDTH/8-1:0] m_axis_oarg_6_tkeep,
    output [M_AXIS_OARG_6_DMWIDTH/8-1:0] m_axis_oarg_6_tstrb,
    output [M_AXIS_OARG_6_DMWIDTH-1:0] m_axis_oarg_6_tdata,
    input m_axis_oarg_6_tready,
    input ap_axis_oarg_6_tlast,
    input ap_axis_oarg_6_tvalid,
    input [M_AXIS_OARG_6_WIDTH/8-1:0] ap_axis_oarg_6_tkeep,
    input [M_AXIS_OARG_6_WIDTH/8-1:0] ap_axis_oarg_6_tstrb,
    input [M_AXIS_OARG_6_WIDTH-1:0] ap_axis_oarg_6_tdata,
    output ap_axis_oarg_6_tready,
    //output AXIS to AXI-Stream interface 7
    input m_axis_oarg_7_aclk,
    input m_axis_oarg_7_aresetn,
    output m_axis_oarg_7_tlast,
    output m_axis_oarg_7_tvalid,
    output [M_AXIS_OARG_7_DMWIDTH/8-1:0] m_axis_oarg_7_tkeep,
    output [M_AXIS_OARG_7_DMWIDTH/8-1:0] m_axis_oarg_7_tstrb,
    output [M_AXIS_OARG_7_DMWIDTH-1:0] m_axis_oarg_7_tdata,
    input m_axis_oarg_7_tready,
    input ap_axis_oarg_7_tlast,
    input ap_axis_oarg_7_tvalid,
    input [M_AXIS_OARG_7_WIDTH/8-1:0] ap_axis_oarg_7_tkeep,
    input [M_AXIS_OARG_7_WIDTH/8-1:0] ap_axis_oarg_7_tstrb,
    input [M_AXIS_OARG_7_WIDTH-1:0] ap_axis_oarg_7_tdata,
    output ap_axis_oarg_7_tready,
    //output AXIS to AXI-Stream interface 8
    input m_axis_oarg_8_aclk,
    input m_axis_oarg_8_aresetn,
    output m_axis_oarg_8_tlast,
    output m_axis_oarg_8_tvalid,
    output [M_AXIS_OARG_8_DMWIDTH/8-1:0] m_axis_oarg_8_tkeep,
    output [M_AXIS_OARG_8_DMWIDTH/8-1:0] m_axis_oarg_8_tstrb,
    output [M_AXIS_OARG_8_DMWIDTH-1:0] m_axis_oarg_8_tdata,
    input m_axis_oarg_8_tready,
    input ap_axis_oarg_8_tlast,
    input ap_axis_oarg_8_tvalid,
    input [M_AXIS_OARG_8_WIDTH/8-1:0] ap_axis_oarg_8_tkeep,
    input [M_AXIS_OARG_8_WIDTH/8-1:0] ap_axis_oarg_8_tstrb,
    input [M_AXIS_OARG_8_WIDTH-1:0] ap_axis_oarg_8_tdata,
    output ap_axis_oarg_8_tready,
    //output AXIS to AXI-Stream interface 9
    input m_axis_oarg_9_aclk,
    input m_axis_oarg_9_aresetn,
    output m_axis_oarg_9_tlast,
    output m_axis_oarg_9_tvalid,
    output [M_AXIS_OARG_9_DMWIDTH/8-1:0] m_axis_oarg_9_tkeep,
    output [M_AXIS_OARG_9_DMWIDTH/8-1:0] m_axis_oarg_9_tstrb,
    output [M_AXIS_OARG_9_DMWIDTH-1:0] m_axis_oarg_9_tdata,
    input m_axis_oarg_9_tready,
    input ap_axis_oarg_9_tlast,
    input ap_axis_oarg_9_tvalid,
    input [M_AXIS_OARG_9_WIDTH/8-1:0] ap_axis_oarg_9_tkeep,
    input [M_AXIS_OARG_9_WIDTH/8-1:0] ap_axis_oarg_9_tstrb,
    input [M_AXIS_OARG_9_WIDTH-1:0] ap_axis_oarg_9_tdata,
    output ap_axis_oarg_9_tready,
    //output AXIS to AXI-Stream interface 10
    input m_axis_oarg_10_aclk,
    input m_axis_oarg_10_aresetn,
    output m_axis_oarg_10_tlast,
    output m_axis_oarg_10_tvalid,
    output [M_AXIS_OARG_10_DMWIDTH/8-1:0] m_axis_oarg_10_tkeep,
    output [M_AXIS_OARG_10_DMWIDTH/8-1:0] m_axis_oarg_10_tstrb,
    output [M_AXIS_OARG_10_DMWIDTH-1:0] m_axis_oarg_10_tdata,
    input m_axis_oarg_10_tready,
    input ap_axis_oarg_10_tlast,
    input ap_axis_oarg_10_tvalid,
    input [M_AXIS_OARG_10_WIDTH/8-1:0] ap_axis_oarg_10_tkeep,
    input [M_AXIS_OARG_10_WIDTH/8-1:0] ap_axis_oarg_10_tstrb,
    input [M_AXIS_OARG_10_WIDTH-1:0] ap_axis_oarg_10_tdata,
    output ap_axis_oarg_10_tready,
    //output AXIS to AXI-Stream interface 11
    input m_axis_oarg_11_aclk,
    input m_axis_oarg_11_aresetn,
    output m_axis_oarg_11_tlast,
    output m_axis_oarg_11_tvalid,
    output [M_AXIS_OARG_11_DMWIDTH/8-1:0] m_axis_oarg_11_tkeep,
    output [M_AXIS_OARG_11_DMWIDTH/8-1:0] m_axis_oarg_11_tstrb,
    output [M_AXIS_OARG_11_DMWIDTH-1:0] m_axis_oarg_11_tdata,
    input m_axis_oarg_11_tready,
    input ap_axis_oarg_11_tlast,
    input ap_axis_oarg_11_tvalid,
    input [M_AXIS_OARG_11_WIDTH/8-1:0] ap_axis_oarg_11_tkeep,
    input [M_AXIS_OARG_11_WIDTH/8-1:0] ap_axis_oarg_11_tstrb,
    input [M_AXIS_OARG_11_WIDTH-1:0] ap_axis_oarg_11_tdata,
    output ap_axis_oarg_11_tready,
    //output AXIS to AXI-Stream interface 12
    input m_axis_oarg_12_aclk,
    input m_axis_oarg_12_aresetn,
    output m_axis_oarg_12_tlast,
    output m_axis_oarg_12_tvalid,
    output [M_AXIS_OARG_12_DMWIDTH/8-1:0] m_axis_oarg_12_tkeep,
    output [M_AXIS_OARG_12_DMWIDTH/8-1:0] m_axis_oarg_12_tstrb,
    output [M_AXIS_OARG_12_DMWIDTH-1:0] m_axis_oarg_12_tdata,
    input m_axis_oarg_12_tready,
    input ap_axis_oarg_12_tlast,
    input ap_axis_oarg_12_tvalid,
    input [M_AXIS_OARG_12_WIDTH/8-1:0] ap_axis_oarg_12_tkeep,
    input [M_AXIS_OARG_12_WIDTH/8-1:0] ap_axis_oarg_12_tstrb,
    input [M_AXIS_OARG_12_WIDTH-1:0] ap_axis_oarg_12_tdata,
    output ap_axis_oarg_12_tready,
    //output AXIS to AXI-Stream interface 13
    input m_axis_oarg_13_aclk,
    input m_axis_oarg_13_aresetn,
    output m_axis_oarg_13_tlast,
    output m_axis_oarg_13_tvalid,
    output [M_AXIS_OARG_13_DMWIDTH/8-1:0] m_axis_oarg_13_tkeep,
    output [M_AXIS_OARG_13_DMWIDTH/8-1:0] m_axis_oarg_13_tstrb,
    output [M_AXIS_OARG_13_DMWIDTH-1:0] m_axis_oarg_13_tdata,
    input m_axis_oarg_13_tready,
    input ap_axis_oarg_13_tlast,
    input ap_axis_oarg_13_tvalid,
    input [M_AXIS_OARG_13_WIDTH/8-1:0] ap_axis_oarg_13_tkeep,
    input [M_AXIS_OARG_13_WIDTH/8-1:0] ap_axis_oarg_13_tstrb,
    input [M_AXIS_OARG_13_WIDTH-1:0] ap_axis_oarg_13_tdata,
    output ap_axis_oarg_13_tready,
    //output AXIS to AXI-Stream interface 14
    input m_axis_oarg_14_aclk,
    input m_axis_oarg_14_aresetn,
    output m_axis_oarg_14_tlast,
    output m_axis_oarg_14_tvalid,
    output [M_AXIS_OARG_14_DMWIDTH/8-1:0] m_axis_oarg_14_tkeep,
    output [M_AXIS_OARG_14_DMWIDTH/8-1:0] m_axis_oarg_14_tstrb,
    output [M_AXIS_OARG_14_DMWIDTH-1:0] m_axis_oarg_14_tdata,
    input m_axis_oarg_14_tready,
    input ap_axis_oarg_14_tlast,
    input ap_axis_oarg_14_tvalid,
    input [M_AXIS_OARG_14_WIDTH/8-1:0] ap_axis_oarg_14_tkeep,
    input [M_AXIS_OARG_14_WIDTH/8-1:0] ap_axis_oarg_14_tstrb,
    input [M_AXIS_OARG_14_WIDTH-1:0] ap_axis_oarg_14_tdata,
    output ap_axis_oarg_14_tready,
    //output AXIS to AXI-Stream interface 15
    input m_axis_oarg_15_aclk,
    input m_axis_oarg_15_aresetn,
    output m_axis_oarg_15_tlast,
    output m_axis_oarg_15_tvalid,
    output [M_AXIS_OARG_15_DMWIDTH/8-1:0] m_axis_oarg_15_tkeep,
    output [M_AXIS_OARG_15_DMWIDTH/8-1:0] m_axis_oarg_15_tstrb,
    output [M_AXIS_OARG_15_DMWIDTH-1:0] m_axis_oarg_15_tdata,
    input m_axis_oarg_15_tready,
    input ap_axis_oarg_15_tlast,
    input ap_axis_oarg_15_tvalid,
    input [M_AXIS_OARG_15_WIDTH/8-1:0] ap_axis_oarg_15_tkeep,
    input [M_AXIS_OARG_15_WIDTH/8-1:0] ap_axis_oarg_15_tstrb,
    input [M_AXIS_OARG_15_WIDTH-1:0] ap_axis_oarg_15_tdata,
    output ap_axis_oarg_15_tready,
    //output AXIS to AXI-Stream interface 16
    input m_axis_oarg_16_aclk,
    input m_axis_oarg_16_aresetn,
    output m_axis_oarg_16_tlast,
    output m_axis_oarg_16_tvalid,
    output [M_AXIS_OARG_16_DMWIDTH/8-1:0] m_axis_oarg_16_tkeep,
    output [M_AXIS_OARG_16_DMWIDTH/8-1:0] m_axis_oarg_16_tstrb,
    output [M_AXIS_OARG_16_DMWIDTH-1:0] m_axis_oarg_16_tdata,
    input m_axis_oarg_16_tready,
    input ap_axis_oarg_16_tlast,
    input ap_axis_oarg_16_tvalid,
    input [M_AXIS_OARG_16_WIDTH/8-1:0] ap_axis_oarg_16_tkeep,
    input [M_AXIS_OARG_16_WIDTH/8-1:0] ap_axis_oarg_16_tstrb,
    input [M_AXIS_OARG_16_WIDTH-1:0] ap_axis_oarg_16_tdata,
    output ap_axis_oarg_16_tready,
    //output AXIS to AXI-Stream interface 17
    input m_axis_oarg_17_aclk,
    input m_axis_oarg_17_aresetn,
    output m_axis_oarg_17_tlast,
    output m_axis_oarg_17_tvalid,
    output [M_AXIS_OARG_17_DMWIDTH/8-1:0] m_axis_oarg_17_tkeep,
    output [M_AXIS_OARG_17_DMWIDTH/8-1:0] m_axis_oarg_17_tstrb,
    output [M_AXIS_OARG_17_DMWIDTH-1:0] m_axis_oarg_17_tdata,
    input m_axis_oarg_17_tready,
    input ap_axis_oarg_17_tlast,
    input ap_axis_oarg_17_tvalid,
    input [M_AXIS_OARG_17_WIDTH/8-1:0] ap_axis_oarg_17_tkeep,
    input [M_AXIS_OARG_17_WIDTH/8-1:0] ap_axis_oarg_17_tstrb,
    input [M_AXIS_OARG_17_WIDTH-1:0] ap_axis_oarg_17_tdata,
    output ap_axis_oarg_17_tready,
    //output AXIS to AXI-Stream interface 18
    input m_axis_oarg_18_aclk,
    input m_axis_oarg_18_aresetn,
    output m_axis_oarg_18_tlast,
    output m_axis_oarg_18_tvalid,
    output [M_AXIS_OARG_18_DMWIDTH/8-1:0] m_axis_oarg_18_tkeep,
    output [M_AXIS_OARG_18_DMWIDTH/8-1:0] m_axis_oarg_18_tstrb,
    output [M_AXIS_OARG_18_DMWIDTH-1:0] m_axis_oarg_18_tdata,
    input m_axis_oarg_18_tready,
    input ap_axis_oarg_18_tlast,
    input ap_axis_oarg_18_tvalid,
    input [M_AXIS_OARG_18_WIDTH/8-1:0] ap_axis_oarg_18_tkeep,
    input [M_AXIS_OARG_18_WIDTH/8-1:0] ap_axis_oarg_18_tstrb,
    input [M_AXIS_OARG_18_WIDTH-1:0] ap_axis_oarg_18_tdata,
    output ap_axis_oarg_18_tready,
    //output AXIS to AXI-Stream interface 19
    input m_axis_oarg_19_aclk,
    input m_axis_oarg_19_aresetn,
    output m_axis_oarg_19_tlast,
    output m_axis_oarg_19_tvalid,
    output [M_AXIS_OARG_19_DMWIDTH/8-1:0] m_axis_oarg_19_tkeep,
    output [M_AXIS_OARG_19_DMWIDTH/8-1:0] m_axis_oarg_19_tstrb,
    output [M_AXIS_OARG_19_DMWIDTH-1:0] m_axis_oarg_19_tdata,
    input m_axis_oarg_19_tready,
    input ap_axis_oarg_19_tlast,
    input ap_axis_oarg_19_tvalid,
    input [M_AXIS_OARG_19_WIDTH/8-1:0] ap_axis_oarg_19_tkeep,
    input [M_AXIS_OARG_19_WIDTH/8-1:0] ap_axis_oarg_19_tstrb,
    input [M_AXIS_OARG_19_WIDTH-1:0] ap_axis_oarg_19_tdata,
    output ap_axis_oarg_19_tready,
    //output AXIS to AXI-Stream interface 20
    input m_axis_oarg_20_aclk,
    input m_axis_oarg_20_aresetn,
    output m_axis_oarg_20_tlast,
    output m_axis_oarg_20_tvalid,
    output [M_AXIS_OARG_20_DMWIDTH/8-1:0] m_axis_oarg_20_tkeep,
    output [M_AXIS_OARG_20_DMWIDTH/8-1:0] m_axis_oarg_20_tstrb,
    output [M_AXIS_OARG_20_DMWIDTH-1:0] m_axis_oarg_20_tdata,
    input m_axis_oarg_20_tready,
    input ap_axis_oarg_20_tlast,
    input ap_axis_oarg_20_tvalid,
    input [M_AXIS_OARG_20_WIDTH/8-1:0] ap_axis_oarg_20_tkeep,
    input [M_AXIS_OARG_20_WIDTH/8-1:0] ap_axis_oarg_20_tstrb,
    input [M_AXIS_OARG_20_WIDTH-1:0] ap_axis_oarg_20_tdata,
    output ap_axis_oarg_20_tready,
    //output AXIS to AXI-Stream interface 21
    input m_axis_oarg_21_aclk,
    input m_axis_oarg_21_aresetn,
    output m_axis_oarg_21_tlast,
    output m_axis_oarg_21_tvalid,
    output [M_AXIS_OARG_21_DMWIDTH/8-1:0] m_axis_oarg_21_tkeep,
    output [M_AXIS_OARG_21_DMWIDTH/8-1:0] m_axis_oarg_21_tstrb,
    output [M_AXIS_OARG_21_DMWIDTH-1:0] m_axis_oarg_21_tdata,
    input m_axis_oarg_21_tready,
    input ap_axis_oarg_21_tlast,
    input ap_axis_oarg_21_tvalid,
    input [M_AXIS_OARG_21_WIDTH/8-1:0] ap_axis_oarg_21_tkeep,
    input [M_AXIS_OARG_21_WIDTH/8-1:0] ap_axis_oarg_21_tstrb,
    input [M_AXIS_OARG_21_WIDTH-1:0] ap_axis_oarg_21_tdata,
    output ap_axis_oarg_21_tready,
    //output AXIS to AXI-Stream interface 22
    input m_axis_oarg_22_aclk,
    input m_axis_oarg_22_aresetn,
    output m_axis_oarg_22_tlast,
    output m_axis_oarg_22_tvalid,
    output [M_AXIS_OARG_22_DMWIDTH/8-1:0] m_axis_oarg_22_tkeep,
    output [M_AXIS_OARG_22_DMWIDTH/8-1:0] m_axis_oarg_22_tstrb,
    output [M_AXIS_OARG_22_DMWIDTH-1:0] m_axis_oarg_22_tdata,
    input m_axis_oarg_22_tready,
    input ap_axis_oarg_22_tlast,
    input ap_axis_oarg_22_tvalid,
    input [M_AXIS_OARG_22_WIDTH/8-1:0] ap_axis_oarg_22_tkeep,
    input [M_AXIS_OARG_22_WIDTH/8-1:0] ap_axis_oarg_22_tstrb,
    input [M_AXIS_OARG_22_WIDTH-1:0] ap_axis_oarg_22_tdata,
    output ap_axis_oarg_22_tready,
    //output AXIS to AXI-Stream interface 23
    input m_axis_oarg_23_aclk,
    input m_axis_oarg_23_aresetn,
    output m_axis_oarg_23_tlast,
    output m_axis_oarg_23_tvalid,
    output [M_AXIS_OARG_23_DMWIDTH/8-1:0] m_axis_oarg_23_tkeep,
    output [M_AXIS_OARG_23_DMWIDTH/8-1:0] m_axis_oarg_23_tstrb,
    output [M_AXIS_OARG_23_DMWIDTH-1:0] m_axis_oarg_23_tdata,
    input m_axis_oarg_23_tready,
    input ap_axis_oarg_23_tlast,
    input ap_axis_oarg_23_tvalid,
    input [M_AXIS_OARG_23_WIDTH/8-1:0] ap_axis_oarg_23_tkeep,
    input [M_AXIS_OARG_23_WIDTH/8-1:0] ap_axis_oarg_23_tstrb,
    input [M_AXIS_OARG_23_WIDTH-1:0] ap_axis_oarg_23_tdata,
    output ap_axis_oarg_23_tready,
    //output AXIS to AXI-Stream interface 24
    input m_axis_oarg_24_aclk,
    input m_axis_oarg_24_aresetn,
    output m_axis_oarg_24_tlast,
    output m_axis_oarg_24_tvalid,
    output [M_AXIS_OARG_24_DMWIDTH/8-1:0] m_axis_oarg_24_tkeep,
    output [M_AXIS_OARG_24_DMWIDTH/8-1:0] m_axis_oarg_24_tstrb,
    output [M_AXIS_OARG_24_DMWIDTH-1:0] m_axis_oarg_24_tdata,
    input m_axis_oarg_24_tready,
    input ap_axis_oarg_24_tlast,
    input ap_axis_oarg_24_tvalid,
    input [M_AXIS_OARG_24_WIDTH/8-1:0] ap_axis_oarg_24_tkeep,
    input [M_AXIS_OARG_24_WIDTH/8-1:0] ap_axis_oarg_24_tstrb,
    input [M_AXIS_OARG_24_WIDTH-1:0] ap_axis_oarg_24_tdata,
    output ap_axis_oarg_24_tready,
    //output AXIS to AXI-Stream interface 25
    input m_axis_oarg_25_aclk,
    input m_axis_oarg_25_aresetn,
    output m_axis_oarg_25_tlast,
    output m_axis_oarg_25_tvalid,
    output [M_AXIS_OARG_25_DMWIDTH/8-1:0] m_axis_oarg_25_tkeep,
    output [M_AXIS_OARG_25_DMWIDTH/8-1:0] m_axis_oarg_25_tstrb,
    output [M_AXIS_OARG_25_DMWIDTH-1:0] m_axis_oarg_25_tdata,
    input m_axis_oarg_25_tready,
    input ap_axis_oarg_25_tlast,
    input ap_axis_oarg_25_tvalid,
    input [M_AXIS_OARG_25_WIDTH/8-1:0] ap_axis_oarg_25_tkeep,
    input [M_AXIS_OARG_25_WIDTH/8-1:0] ap_axis_oarg_25_tstrb,
    input [M_AXIS_OARG_25_WIDTH-1:0] ap_axis_oarg_25_tdata,
    output ap_axis_oarg_25_tready,
    //output AXIS to AXI-Stream interface 26
    input m_axis_oarg_26_aclk,
    input m_axis_oarg_26_aresetn,
    output m_axis_oarg_26_tlast,
    output m_axis_oarg_26_tvalid,
    output [M_AXIS_OARG_26_DMWIDTH/8-1:0] m_axis_oarg_26_tkeep,
    output [M_AXIS_OARG_26_DMWIDTH/8-1:0] m_axis_oarg_26_tstrb,
    output [M_AXIS_OARG_26_DMWIDTH-1:0] m_axis_oarg_26_tdata,
    input m_axis_oarg_26_tready,
    input ap_axis_oarg_26_tlast,
    input ap_axis_oarg_26_tvalid,
    input [M_AXIS_OARG_26_WIDTH/8-1:0] ap_axis_oarg_26_tkeep,
    input [M_AXIS_OARG_26_WIDTH/8-1:0] ap_axis_oarg_26_tstrb,
    input [M_AXIS_OARG_26_WIDTH-1:0] ap_axis_oarg_26_tdata,
    output ap_axis_oarg_26_tready,
    //output AXIS to AXI-Stream interface 27
    input m_axis_oarg_27_aclk,
    input m_axis_oarg_27_aresetn,
    output m_axis_oarg_27_tlast,
    output m_axis_oarg_27_tvalid,
    output [M_AXIS_OARG_27_DMWIDTH/8-1:0] m_axis_oarg_27_tkeep,
    output [M_AXIS_OARG_27_DMWIDTH/8-1:0] m_axis_oarg_27_tstrb,
    output [M_AXIS_OARG_27_DMWIDTH-1:0] m_axis_oarg_27_tdata,
    input m_axis_oarg_27_tready,
    input ap_axis_oarg_27_tlast,
    input ap_axis_oarg_27_tvalid,
    input [M_AXIS_OARG_27_WIDTH/8-1:0] ap_axis_oarg_27_tkeep,
    input [M_AXIS_OARG_27_WIDTH/8-1:0] ap_axis_oarg_27_tstrb,
    input [M_AXIS_OARG_27_WIDTH-1:0] ap_axis_oarg_27_tdata,
    output ap_axis_oarg_27_tready,
    //output AXIS to AXI-Stream interface 28
    input m_axis_oarg_28_aclk,
    input m_axis_oarg_28_aresetn,
    output m_axis_oarg_28_tlast,
    output m_axis_oarg_28_tvalid,
    output [M_AXIS_OARG_28_DMWIDTH/8-1:0] m_axis_oarg_28_tkeep,
    output [M_AXIS_OARG_28_DMWIDTH/8-1:0] m_axis_oarg_28_tstrb,
    output [M_AXIS_OARG_28_DMWIDTH-1:0] m_axis_oarg_28_tdata,
    input m_axis_oarg_28_tready,
    input ap_axis_oarg_28_tlast,
    input ap_axis_oarg_28_tvalid,
    input [M_AXIS_OARG_28_WIDTH/8-1:0] ap_axis_oarg_28_tkeep,
    input [M_AXIS_OARG_28_WIDTH/8-1:0] ap_axis_oarg_28_tstrb,
    input [M_AXIS_OARG_28_WIDTH-1:0] ap_axis_oarg_28_tdata,
    output ap_axis_oarg_28_tready,
    //output AXIS to AXI-Stream interface 29
    input m_axis_oarg_29_aclk,
    input m_axis_oarg_29_aresetn,
    output m_axis_oarg_29_tlast,
    output m_axis_oarg_29_tvalid,
    output [M_AXIS_OARG_29_DMWIDTH/8-1:0] m_axis_oarg_29_tkeep,
    output [M_AXIS_OARG_29_DMWIDTH/8-1:0] m_axis_oarg_29_tstrb,
    output [M_AXIS_OARG_29_DMWIDTH-1:0] m_axis_oarg_29_tdata,
    input m_axis_oarg_29_tready,
    input ap_axis_oarg_29_tlast,
    input ap_axis_oarg_29_tvalid,
    input [M_AXIS_OARG_29_WIDTH/8-1:0] ap_axis_oarg_29_tkeep,
    input [M_AXIS_OARG_29_WIDTH/8-1:0] ap_axis_oarg_29_tstrb,
    input [M_AXIS_OARG_29_WIDTH-1:0] ap_axis_oarg_29_tdata,
    output ap_axis_oarg_29_tready,
    //output AXIS to AXI-Stream interface 30
    input m_axis_oarg_30_aclk,
    input m_axis_oarg_30_aresetn,
    output m_axis_oarg_30_tlast,
    output m_axis_oarg_30_tvalid,
    output [M_AXIS_OARG_30_DMWIDTH/8-1:0] m_axis_oarg_30_tkeep,
    output [M_AXIS_OARG_30_DMWIDTH/8-1:0] m_axis_oarg_30_tstrb,
    output [M_AXIS_OARG_30_DMWIDTH-1:0] m_axis_oarg_30_tdata,
    input m_axis_oarg_30_tready,
    input ap_axis_oarg_30_tlast,
    input ap_axis_oarg_30_tvalid,
    input [M_AXIS_OARG_30_WIDTH/8-1:0] ap_axis_oarg_30_tkeep,
    input [M_AXIS_OARG_30_WIDTH/8-1:0] ap_axis_oarg_30_tstrb,
    input [M_AXIS_OARG_30_WIDTH-1:0] ap_axis_oarg_30_tdata,
    output ap_axis_oarg_30_tready,
    //output AXIS to AXI-Stream interface 31
    input m_axis_oarg_31_aclk,
    input m_axis_oarg_31_aresetn,
    output m_axis_oarg_31_tlast,
    output m_axis_oarg_31_tvalid,
    output [M_AXIS_OARG_31_DMWIDTH/8-1:0] m_axis_oarg_31_tkeep,
    output [M_AXIS_OARG_31_DMWIDTH/8-1:0] m_axis_oarg_31_tstrb,
    output [M_AXIS_OARG_31_DMWIDTH-1:0] m_axis_oarg_31_tdata,
    input m_axis_oarg_31_tready,
    input ap_axis_oarg_31_tlast,
    input ap_axis_oarg_31_tvalid,
    input [M_AXIS_OARG_31_WIDTH/8-1:0] ap_axis_oarg_31_tkeep,
    input [M_AXIS_OARG_31_WIDTH/8-1:0] ap_axis_oarg_31_tstrb,
    input [M_AXIS_OARG_31_WIDTH-1:0] ap_axis_oarg_31_tdata,
    output ap_axis_oarg_31_tready,
    //output AXIS to AXI-Stream interface 32
    input m_axis_oarg_32_aclk,
    input m_axis_oarg_32_aresetn,
    output m_axis_oarg_32_tlast,
    output m_axis_oarg_32_tvalid,
    output [M_AXIS_OARG_32_DMWIDTH/8-1:0] m_axis_oarg_32_tkeep,
    output [M_AXIS_OARG_32_DMWIDTH/8-1:0] m_axis_oarg_32_tstrb,
    output [M_AXIS_OARG_32_DMWIDTH-1:0] m_axis_oarg_32_tdata,
    input m_axis_oarg_32_tready,
    input ap_axis_oarg_32_tlast,
    input ap_axis_oarg_32_tvalid,
    input [M_AXIS_OARG_32_WIDTH/8-1:0] ap_axis_oarg_32_tkeep,
    input [M_AXIS_OARG_32_WIDTH/8-1:0] ap_axis_oarg_32_tstrb,
    input [M_AXIS_OARG_32_WIDTH-1:0] ap_axis_oarg_32_tdata,
    output ap_axis_oarg_32_tready,
    //output AXIS to AXI-Stream interface 33
    input m_axis_oarg_33_aclk,
    input m_axis_oarg_33_aresetn,
    output m_axis_oarg_33_tlast,
    output m_axis_oarg_33_tvalid,
    output [M_AXIS_OARG_33_DMWIDTH/8-1:0] m_axis_oarg_33_tkeep,
    output [M_AXIS_OARG_33_DMWIDTH/8-1:0] m_axis_oarg_33_tstrb,
    output [M_AXIS_OARG_33_DMWIDTH-1:0] m_axis_oarg_33_tdata,
    input m_axis_oarg_33_tready,
    input ap_axis_oarg_33_tlast,
    input ap_axis_oarg_33_tvalid,
    input [M_AXIS_OARG_33_WIDTH/8-1:0] ap_axis_oarg_33_tkeep,
    input [M_AXIS_OARG_33_WIDTH/8-1:0] ap_axis_oarg_33_tstrb,
    input [M_AXIS_OARG_33_WIDTH-1:0] ap_axis_oarg_33_tdata,
    output ap_axis_oarg_33_tready,
    //output AXIS to AXI-Stream interface 34
    input m_axis_oarg_34_aclk,
    input m_axis_oarg_34_aresetn,
    output m_axis_oarg_34_tlast,
    output m_axis_oarg_34_tvalid,
    output [M_AXIS_OARG_34_DMWIDTH/8-1:0] m_axis_oarg_34_tkeep,
    output [M_AXIS_OARG_34_DMWIDTH/8-1:0] m_axis_oarg_34_tstrb,
    output [M_AXIS_OARG_34_DMWIDTH-1:0] m_axis_oarg_34_tdata,
    input m_axis_oarg_34_tready,
    input ap_axis_oarg_34_tlast,
    input ap_axis_oarg_34_tvalid,
    input [M_AXIS_OARG_34_WIDTH/8-1:0] ap_axis_oarg_34_tkeep,
    input [M_AXIS_OARG_34_WIDTH/8-1:0] ap_axis_oarg_34_tstrb,
    input [M_AXIS_OARG_34_WIDTH-1:0] ap_axis_oarg_34_tdata,
    output ap_axis_oarg_34_tready,
    //output AXIS to AXI-Stream interface 35
    input m_axis_oarg_35_aclk,
    input m_axis_oarg_35_aresetn,
    output m_axis_oarg_35_tlast,
    output m_axis_oarg_35_tvalid,
    output [M_AXIS_OARG_35_DMWIDTH/8-1:0] m_axis_oarg_35_tkeep,
    output [M_AXIS_OARG_35_DMWIDTH/8-1:0] m_axis_oarg_35_tstrb,
    output [M_AXIS_OARG_35_DMWIDTH-1:0] m_axis_oarg_35_tdata,
    input m_axis_oarg_35_tready,
    input ap_axis_oarg_35_tlast,
    input ap_axis_oarg_35_tvalid,
    input [M_AXIS_OARG_35_WIDTH/8-1:0] ap_axis_oarg_35_tkeep,
    input [M_AXIS_OARG_35_WIDTH/8-1:0] ap_axis_oarg_35_tstrb,
    input [M_AXIS_OARG_35_WIDTH-1:0] ap_axis_oarg_35_tdata,
    output ap_axis_oarg_35_tready,
    //output AXIS to AXI-Stream interface 36
    input m_axis_oarg_36_aclk,
    input m_axis_oarg_36_aresetn,
    output m_axis_oarg_36_tlast,
    output m_axis_oarg_36_tvalid,
    output [M_AXIS_OARG_36_DMWIDTH/8-1:0] m_axis_oarg_36_tkeep,
    output [M_AXIS_OARG_36_DMWIDTH/8-1:0] m_axis_oarg_36_tstrb,
    output [M_AXIS_OARG_36_DMWIDTH-1:0] m_axis_oarg_36_tdata,
    input m_axis_oarg_36_tready,
    input ap_axis_oarg_36_tlast,
    input ap_axis_oarg_36_tvalid,
    input [M_AXIS_OARG_36_WIDTH/8-1:0] ap_axis_oarg_36_tkeep,
    input [M_AXIS_OARG_36_WIDTH/8-1:0] ap_axis_oarg_36_tstrb,
    input [M_AXIS_OARG_36_WIDTH-1:0] ap_axis_oarg_36_tdata,
    output ap_axis_oarg_36_tready,
    //output AXIS to AXI-Stream interface 37
    input m_axis_oarg_37_aclk,
    input m_axis_oarg_37_aresetn,
    output m_axis_oarg_37_tlast,
    output m_axis_oarg_37_tvalid,
    output [M_AXIS_OARG_37_DMWIDTH/8-1:0] m_axis_oarg_37_tkeep,
    output [M_AXIS_OARG_37_DMWIDTH/8-1:0] m_axis_oarg_37_tstrb,
    output [M_AXIS_OARG_37_DMWIDTH-1:0] m_axis_oarg_37_tdata,
    input m_axis_oarg_37_tready,
    input ap_axis_oarg_37_tlast,
    input ap_axis_oarg_37_tvalid,
    input [M_AXIS_OARG_37_WIDTH/8-1:0] ap_axis_oarg_37_tkeep,
    input [M_AXIS_OARG_37_WIDTH/8-1:0] ap_axis_oarg_37_tstrb,
    input [M_AXIS_OARG_37_WIDTH-1:0] ap_axis_oarg_37_tdata,
    output ap_axis_oarg_37_tready,
    //output AXIS to AXI-Stream interface 38
    input m_axis_oarg_38_aclk,
    input m_axis_oarg_38_aresetn,
    output m_axis_oarg_38_tlast,
    output m_axis_oarg_38_tvalid,
    output [M_AXIS_OARG_38_DMWIDTH/8-1:0] m_axis_oarg_38_tkeep,
    output [M_AXIS_OARG_38_DMWIDTH/8-1:0] m_axis_oarg_38_tstrb,
    output [M_AXIS_OARG_38_DMWIDTH-1:0] m_axis_oarg_38_tdata,
    input m_axis_oarg_38_tready,
    input ap_axis_oarg_38_tlast,
    input ap_axis_oarg_38_tvalid,
    input [M_AXIS_OARG_38_WIDTH/8-1:0] ap_axis_oarg_38_tkeep,
    input [M_AXIS_OARG_38_WIDTH/8-1:0] ap_axis_oarg_38_tstrb,
    input [M_AXIS_OARG_38_WIDTH-1:0] ap_axis_oarg_38_tdata,
    output ap_axis_oarg_38_tready,
    //output AXIS to AXI-Stream interface 39
    input m_axis_oarg_39_aclk,
    input m_axis_oarg_39_aresetn,
    output m_axis_oarg_39_tlast,
    output m_axis_oarg_39_tvalid,
    output [M_AXIS_OARG_39_DMWIDTH/8-1:0] m_axis_oarg_39_tkeep,
    output [M_AXIS_OARG_39_DMWIDTH/8-1:0] m_axis_oarg_39_tstrb,
    output [M_AXIS_OARG_39_DMWIDTH-1:0] m_axis_oarg_39_tdata,
    input m_axis_oarg_39_tready,
    input ap_axis_oarg_39_tlast,
    input ap_axis_oarg_39_tvalid,
    input [M_AXIS_OARG_39_WIDTH/8-1:0] ap_axis_oarg_39_tkeep,
    input [M_AXIS_OARG_39_WIDTH/8-1:0] ap_axis_oarg_39_tstrb,
    input [M_AXIS_OARG_39_WIDTH-1:0] ap_axis_oarg_39_tdata,
    output ap_axis_oarg_39_tready,
    //output AXIS to AXI-Stream interface 40
    input m_axis_oarg_40_aclk,
    input m_axis_oarg_40_aresetn,
    output m_axis_oarg_40_tlast,
    output m_axis_oarg_40_tvalid,
    output [M_AXIS_OARG_40_DMWIDTH/8-1:0] m_axis_oarg_40_tkeep,
    output [M_AXIS_OARG_40_DMWIDTH/8-1:0] m_axis_oarg_40_tstrb,
    output [M_AXIS_OARG_40_DMWIDTH-1:0] m_axis_oarg_40_tdata,
    input m_axis_oarg_40_tready,
    input ap_axis_oarg_40_tlast,
    input ap_axis_oarg_40_tvalid,
    input [M_AXIS_OARG_40_WIDTH/8-1:0] ap_axis_oarg_40_tkeep,
    input [M_AXIS_OARG_40_WIDTH/8-1:0] ap_axis_oarg_40_tstrb,
    input [M_AXIS_OARG_40_WIDTH-1:0] ap_axis_oarg_40_tdata,
    output ap_axis_oarg_40_tready,
    //output AXIS to AXI-Stream interface 41
    input m_axis_oarg_41_aclk,
    input m_axis_oarg_41_aresetn,
    output m_axis_oarg_41_tlast,
    output m_axis_oarg_41_tvalid,
    output [M_AXIS_OARG_41_DMWIDTH/8-1:0] m_axis_oarg_41_tkeep,
    output [M_AXIS_OARG_41_DMWIDTH/8-1:0] m_axis_oarg_41_tstrb,
    output [M_AXIS_OARG_41_DMWIDTH-1:0] m_axis_oarg_41_tdata,
    input m_axis_oarg_41_tready,
    input ap_axis_oarg_41_tlast,
    input ap_axis_oarg_41_tvalid,
    input [M_AXIS_OARG_41_WIDTH/8-1:0] ap_axis_oarg_41_tkeep,
    input [M_AXIS_OARG_41_WIDTH/8-1:0] ap_axis_oarg_41_tstrb,
    input [M_AXIS_OARG_41_WIDTH-1:0] ap_axis_oarg_41_tdata,
    output ap_axis_oarg_41_tready,
    //output AXIS to AXI-Stream interface 42
    input m_axis_oarg_42_aclk,
    input m_axis_oarg_42_aresetn,
    output m_axis_oarg_42_tlast,
    output m_axis_oarg_42_tvalid,
    output [M_AXIS_OARG_42_DMWIDTH/8-1:0] m_axis_oarg_42_tkeep,
    output [M_AXIS_OARG_42_DMWIDTH/8-1:0] m_axis_oarg_42_tstrb,
    output [M_AXIS_OARG_42_DMWIDTH-1:0] m_axis_oarg_42_tdata,
    input m_axis_oarg_42_tready,
    input ap_axis_oarg_42_tlast,
    input ap_axis_oarg_42_tvalid,
    input [M_AXIS_OARG_42_WIDTH/8-1:0] ap_axis_oarg_42_tkeep,
    input [M_AXIS_OARG_42_WIDTH/8-1:0] ap_axis_oarg_42_tstrb,
    input [M_AXIS_OARG_42_WIDTH-1:0] ap_axis_oarg_42_tdata,
    output ap_axis_oarg_42_tready,
    //output AXIS to AXI-Stream interface 43
    input m_axis_oarg_43_aclk,
    input m_axis_oarg_43_aresetn,
    output m_axis_oarg_43_tlast,
    output m_axis_oarg_43_tvalid,
    output [M_AXIS_OARG_43_DMWIDTH/8-1:0] m_axis_oarg_43_tkeep,
    output [M_AXIS_OARG_43_DMWIDTH/8-1:0] m_axis_oarg_43_tstrb,
    output [M_AXIS_OARG_43_DMWIDTH-1:0] m_axis_oarg_43_tdata,
    input m_axis_oarg_43_tready,
    input ap_axis_oarg_43_tlast,
    input ap_axis_oarg_43_tvalid,
    input [M_AXIS_OARG_43_WIDTH/8-1:0] ap_axis_oarg_43_tkeep,
    input [M_AXIS_OARG_43_WIDTH/8-1:0] ap_axis_oarg_43_tstrb,
    input [M_AXIS_OARG_43_WIDTH-1:0] ap_axis_oarg_43_tdata,
    output ap_axis_oarg_43_tready,
    //output AXIS to AXI-Stream interface 44
    input m_axis_oarg_44_aclk,
    input m_axis_oarg_44_aresetn,
    output m_axis_oarg_44_tlast,
    output m_axis_oarg_44_tvalid,
    output [M_AXIS_OARG_44_DMWIDTH/8-1:0] m_axis_oarg_44_tkeep,
    output [M_AXIS_OARG_44_DMWIDTH/8-1:0] m_axis_oarg_44_tstrb,
    output [M_AXIS_OARG_44_DMWIDTH-1:0] m_axis_oarg_44_tdata,
    input m_axis_oarg_44_tready,
    input ap_axis_oarg_44_tlast,
    input ap_axis_oarg_44_tvalid,
    input [M_AXIS_OARG_44_WIDTH/8-1:0] ap_axis_oarg_44_tkeep,
    input [M_AXIS_OARG_44_WIDTH/8-1:0] ap_axis_oarg_44_tstrb,
    input [M_AXIS_OARG_44_WIDTH-1:0] ap_axis_oarg_44_tdata,
    output ap_axis_oarg_44_tready,
    //output AXIS to AXI-Stream interface 45
    input m_axis_oarg_45_aclk,
    input m_axis_oarg_45_aresetn,
    output m_axis_oarg_45_tlast,
    output m_axis_oarg_45_tvalid,
    output [M_AXIS_OARG_45_DMWIDTH/8-1:0] m_axis_oarg_45_tkeep,
    output [M_AXIS_OARG_45_DMWIDTH/8-1:0] m_axis_oarg_45_tstrb,
    output [M_AXIS_OARG_45_DMWIDTH-1:0] m_axis_oarg_45_tdata,
    input m_axis_oarg_45_tready,
    input ap_axis_oarg_45_tlast,
    input ap_axis_oarg_45_tvalid,
    input [M_AXIS_OARG_45_WIDTH/8-1:0] ap_axis_oarg_45_tkeep,
    input [M_AXIS_OARG_45_WIDTH/8-1:0] ap_axis_oarg_45_tstrb,
    input [M_AXIS_OARG_45_WIDTH-1:0] ap_axis_oarg_45_tdata,
    output ap_axis_oarg_45_tready,
    //output AXIS to AXI-Stream interface 46
    input m_axis_oarg_46_aclk,
    input m_axis_oarg_46_aresetn,
    output m_axis_oarg_46_tlast,
    output m_axis_oarg_46_tvalid,
    output [M_AXIS_OARG_46_DMWIDTH/8-1:0] m_axis_oarg_46_tkeep,
    output [M_AXIS_OARG_46_DMWIDTH/8-1:0] m_axis_oarg_46_tstrb,
    output [M_AXIS_OARG_46_DMWIDTH-1:0] m_axis_oarg_46_tdata,
    input m_axis_oarg_46_tready,
    input ap_axis_oarg_46_tlast,
    input ap_axis_oarg_46_tvalid,
    input [M_AXIS_OARG_46_WIDTH/8-1:0] ap_axis_oarg_46_tkeep,
    input [M_AXIS_OARG_46_WIDTH/8-1:0] ap_axis_oarg_46_tstrb,
    input [M_AXIS_OARG_46_WIDTH-1:0] ap_axis_oarg_46_tdata,
    output ap_axis_oarg_46_tready,
    //output AXIS to AXI-Stream interface 47
    input m_axis_oarg_47_aclk,
    input m_axis_oarg_47_aresetn,
    output m_axis_oarg_47_tlast,
    output m_axis_oarg_47_tvalid,
    output [M_AXIS_OARG_47_DMWIDTH/8-1:0] m_axis_oarg_47_tkeep,
    output [M_AXIS_OARG_47_DMWIDTH/8-1:0] m_axis_oarg_47_tstrb,
    output [M_AXIS_OARG_47_DMWIDTH-1:0] m_axis_oarg_47_tdata,
    input m_axis_oarg_47_tready,
    input ap_axis_oarg_47_tlast,
    input ap_axis_oarg_47_tvalid,
    input [M_AXIS_OARG_47_WIDTH/8-1:0] ap_axis_oarg_47_tkeep,
    input [M_AXIS_OARG_47_WIDTH/8-1:0] ap_axis_oarg_47_tstrb,
    input [M_AXIS_OARG_47_WIDTH-1:0] ap_axis_oarg_47_tdata,
    output ap_axis_oarg_47_tready,
    //output AXIS to AXI-Stream interface 48
    input m_axis_oarg_48_aclk,
    input m_axis_oarg_48_aresetn,
    output m_axis_oarg_48_tlast,
    output m_axis_oarg_48_tvalid,
    output [M_AXIS_OARG_48_DMWIDTH/8-1:0] m_axis_oarg_48_tkeep,
    output [M_AXIS_OARG_48_DMWIDTH/8-1:0] m_axis_oarg_48_tstrb,
    output [M_AXIS_OARG_48_DMWIDTH-1:0] m_axis_oarg_48_tdata,
    input m_axis_oarg_48_tready,
    input ap_axis_oarg_48_tlast,
    input ap_axis_oarg_48_tvalid,
    input [M_AXIS_OARG_48_WIDTH/8-1:0] ap_axis_oarg_48_tkeep,
    input [M_AXIS_OARG_48_WIDTH/8-1:0] ap_axis_oarg_48_tstrb,
    input [M_AXIS_OARG_48_WIDTH-1:0] ap_axis_oarg_48_tdata,
    output ap_axis_oarg_48_tready,
    //output AXIS to AXI-Stream interface 49
    input m_axis_oarg_49_aclk,
    input m_axis_oarg_49_aresetn,
    output m_axis_oarg_49_tlast,
    output m_axis_oarg_49_tvalid,
    output [M_AXIS_OARG_49_DMWIDTH/8-1:0] m_axis_oarg_49_tkeep,
    output [M_AXIS_OARG_49_DMWIDTH/8-1:0] m_axis_oarg_49_tstrb,
    output [M_AXIS_OARG_49_DMWIDTH-1:0] m_axis_oarg_49_tdata,
    input m_axis_oarg_49_tready,
    input ap_axis_oarg_49_tlast,
    input ap_axis_oarg_49_tvalid,
    input [M_AXIS_OARG_49_WIDTH/8-1:0] ap_axis_oarg_49_tkeep,
    input [M_AXIS_OARG_49_WIDTH/8-1:0] ap_axis_oarg_49_tstrb,
    input [M_AXIS_OARG_49_WIDTH-1:0] ap_axis_oarg_49_tdata,
    output ap_axis_oarg_49_tready,
    //output AXIS to AXI-Stream interface 50
    input m_axis_oarg_50_aclk,
    input m_axis_oarg_50_aresetn,
    output m_axis_oarg_50_tlast,
    output m_axis_oarg_50_tvalid,
    output [M_AXIS_OARG_50_DMWIDTH/8-1:0] m_axis_oarg_50_tkeep,
    output [M_AXIS_OARG_50_DMWIDTH/8-1:0] m_axis_oarg_50_tstrb,
    output [M_AXIS_OARG_50_DMWIDTH-1:0] m_axis_oarg_50_tdata,
    input m_axis_oarg_50_tready,
    input ap_axis_oarg_50_tlast,
    input ap_axis_oarg_50_tvalid,
    input [M_AXIS_OARG_50_WIDTH/8-1:0] ap_axis_oarg_50_tkeep,
    input [M_AXIS_OARG_50_WIDTH/8-1:0] ap_axis_oarg_50_tstrb,
    input [M_AXIS_OARG_50_WIDTH-1:0] ap_axis_oarg_50_tdata,
    output ap_axis_oarg_50_tready,
    //output AXIS to AXI-Stream interface 51
    input m_axis_oarg_51_aclk,
    input m_axis_oarg_51_aresetn,
    output m_axis_oarg_51_tlast,
    output m_axis_oarg_51_tvalid,
    output [M_AXIS_OARG_51_DMWIDTH/8-1:0] m_axis_oarg_51_tkeep,
    output [M_AXIS_OARG_51_DMWIDTH/8-1:0] m_axis_oarg_51_tstrb,
    output [M_AXIS_OARG_51_DMWIDTH-1:0] m_axis_oarg_51_tdata,
    input m_axis_oarg_51_tready,
    input ap_axis_oarg_51_tlast,
    input ap_axis_oarg_51_tvalid,
    input [M_AXIS_OARG_51_WIDTH/8-1:0] ap_axis_oarg_51_tkeep,
    input [M_AXIS_OARG_51_WIDTH/8-1:0] ap_axis_oarg_51_tstrb,
    input [M_AXIS_OARG_51_WIDTH-1:0] ap_axis_oarg_51_tdata,
    output ap_axis_oarg_51_tready,
    //output AXIS to AXI-Stream interface 52
    input m_axis_oarg_52_aclk,
    input m_axis_oarg_52_aresetn,
    output m_axis_oarg_52_tlast,
    output m_axis_oarg_52_tvalid,
    output [M_AXIS_OARG_52_DMWIDTH/8-1:0] m_axis_oarg_52_tkeep,
    output [M_AXIS_OARG_52_DMWIDTH/8-1:0] m_axis_oarg_52_tstrb,
    output [M_AXIS_OARG_52_DMWIDTH-1:0] m_axis_oarg_52_tdata,
    input m_axis_oarg_52_tready,
    input ap_axis_oarg_52_tlast,
    input ap_axis_oarg_52_tvalid,
    input [M_AXIS_OARG_52_WIDTH/8-1:0] ap_axis_oarg_52_tkeep,
    input [M_AXIS_OARG_52_WIDTH/8-1:0] ap_axis_oarg_52_tstrb,
    input [M_AXIS_OARG_52_WIDTH-1:0] ap_axis_oarg_52_tdata,
    output ap_axis_oarg_52_tready,
    //output AXIS to AXI-Stream interface 53
    input m_axis_oarg_53_aclk,
    input m_axis_oarg_53_aresetn,
    output m_axis_oarg_53_tlast,
    output m_axis_oarg_53_tvalid,
    output [M_AXIS_OARG_53_DMWIDTH/8-1:0] m_axis_oarg_53_tkeep,
    output [M_AXIS_OARG_53_DMWIDTH/8-1:0] m_axis_oarg_53_tstrb,
    output [M_AXIS_OARG_53_DMWIDTH-1:0] m_axis_oarg_53_tdata,
    input m_axis_oarg_53_tready,
    input ap_axis_oarg_53_tlast,
    input ap_axis_oarg_53_tvalid,
    input [M_AXIS_OARG_53_WIDTH/8-1:0] ap_axis_oarg_53_tkeep,
    input [M_AXIS_OARG_53_WIDTH/8-1:0] ap_axis_oarg_53_tstrb,
    input [M_AXIS_OARG_53_WIDTH-1:0] ap_axis_oarg_53_tdata,
    output ap_axis_oarg_53_tready,
    //output AXIS to AXI-Stream interface 54
    input m_axis_oarg_54_aclk,
    input m_axis_oarg_54_aresetn,
    output m_axis_oarg_54_tlast,
    output m_axis_oarg_54_tvalid,
    output [M_AXIS_OARG_54_DMWIDTH/8-1:0] m_axis_oarg_54_tkeep,
    output [M_AXIS_OARG_54_DMWIDTH/8-1:0] m_axis_oarg_54_tstrb,
    output [M_AXIS_OARG_54_DMWIDTH-1:0] m_axis_oarg_54_tdata,
    input m_axis_oarg_54_tready,
    input ap_axis_oarg_54_tlast,
    input ap_axis_oarg_54_tvalid,
    input [M_AXIS_OARG_54_WIDTH/8-1:0] ap_axis_oarg_54_tkeep,
    input [M_AXIS_OARG_54_WIDTH/8-1:0] ap_axis_oarg_54_tstrb,
    input [M_AXIS_OARG_54_WIDTH-1:0] ap_axis_oarg_54_tdata,
    output ap_axis_oarg_54_tready,
    //output AXIS to AXI-Stream interface 55
    input m_axis_oarg_55_aclk,
    input m_axis_oarg_55_aresetn,
    output m_axis_oarg_55_tlast,
    output m_axis_oarg_55_tvalid,
    output [M_AXIS_OARG_55_DMWIDTH/8-1:0] m_axis_oarg_55_tkeep,
    output [M_AXIS_OARG_55_DMWIDTH/8-1:0] m_axis_oarg_55_tstrb,
    output [M_AXIS_OARG_55_DMWIDTH-1:0] m_axis_oarg_55_tdata,
    input m_axis_oarg_55_tready,
    input ap_axis_oarg_55_tlast,
    input ap_axis_oarg_55_tvalid,
    input [M_AXIS_OARG_55_WIDTH/8-1:0] ap_axis_oarg_55_tkeep,
    input [M_AXIS_OARG_55_WIDTH/8-1:0] ap_axis_oarg_55_tstrb,
    input [M_AXIS_OARG_55_WIDTH-1:0] ap_axis_oarg_55_tdata,
    output ap_axis_oarg_55_tready,
    //output AXIS to AXI-Stream interface 56
    input m_axis_oarg_56_aclk,
    input m_axis_oarg_56_aresetn,
    output m_axis_oarg_56_tlast,
    output m_axis_oarg_56_tvalid,
    output [M_AXIS_OARG_56_DMWIDTH/8-1:0] m_axis_oarg_56_tkeep,
    output [M_AXIS_OARG_56_DMWIDTH/8-1:0] m_axis_oarg_56_tstrb,
    output [M_AXIS_OARG_56_DMWIDTH-1:0] m_axis_oarg_56_tdata,
    input m_axis_oarg_56_tready,
    input ap_axis_oarg_56_tlast,
    input ap_axis_oarg_56_tvalid,
    input [M_AXIS_OARG_56_WIDTH/8-1:0] ap_axis_oarg_56_tkeep,
    input [M_AXIS_OARG_56_WIDTH/8-1:0] ap_axis_oarg_56_tstrb,
    input [M_AXIS_OARG_56_WIDTH-1:0] ap_axis_oarg_56_tdata,
    output ap_axis_oarg_56_tready,
    //output AXIS to AXI-Stream interface 57
    input m_axis_oarg_57_aclk,
    input m_axis_oarg_57_aresetn,
    output m_axis_oarg_57_tlast,
    output m_axis_oarg_57_tvalid,
    output [M_AXIS_OARG_57_DMWIDTH/8-1:0] m_axis_oarg_57_tkeep,
    output [M_AXIS_OARG_57_DMWIDTH/8-1:0] m_axis_oarg_57_tstrb,
    output [M_AXIS_OARG_57_DMWIDTH-1:0] m_axis_oarg_57_tdata,
    input m_axis_oarg_57_tready,
    input ap_axis_oarg_57_tlast,
    input ap_axis_oarg_57_tvalid,
    input [M_AXIS_OARG_57_WIDTH/8-1:0] ap_axis_oarg_57_tkeep,
    input [M_AXIS_OARG_57_WIDTH/8-1:0] ap_axis_oarg_57_tstrb,
    input [M_AXIS_OARG_57_WIDTH-1:0] ap_axis_oarg_57_tdata,
    output ap_axis_oarg_57_tready,
    //output AXIS to AXI-Stream interface 58
    input m_axis_oarg_58_aclk,
    input m_axis_oarg_58_aresetn,
    output m_axis_oarg_58_tlast,
    output m_axis_oarg_58_tvalid,
    output [M_AXIS_OARG_58_DMWIDTH/8-1:0] m_axis_oarg_58_tkeep,
    output [M_AXIS_OARG_58_DMWIDTH/8-1:0] m_axis_oarg_58_tstrb,
    output [M_AXIS_OARG_58_DMWIDTH-1:0] m_axis_oarg_58_tdata,
    input m_axis_oarg_58_tready,
    input ap_axis_oarg_58_tlast,
    input ap_axis_oarg_58_tvalid,
    input [M_AXIS_OARG_58_WIDTH/8-1:0] ap_axis_oarg_58_tkeep,
    input [M_AXIS_OARG_58_WIDTH/8-1:0] ap_axis_oarg_58_tstrb,
    input [M_AXIS_OARG_58_WIDTH-1:0] ap_axis_oarg_58_tdata,
    output ap_axis_oarg_58_tready,
    //output AXIS to AXI-Stream interface 59
    input m_axis_oarg_59_aclk,
    input m_axis_oarg_59_aresetn,
    output m_axis_oarg_59_tlast,
    output m_axis_oarg_59_tvalid,
    output [M_AXIS_OARG_59_DMWIDTH/8-1:0] m_axis_oarg_59_tkeep,
    output [M_AXIS_OARG_59_DMWIDTH/8-1:0] m_axis_oarg_59_tstrb,
    output [M_AXIS_OARG_59_DMWIDTH-1:0] m_axis_oarg_59_tdata,
    input m_axis_oarg_59_tready,
    input ap_axis_oarg_59_tlast,
    input ap_axis_oarg_59_tvalid,
    input [M_AXIS_OARG_59_WIDTH/8-1:0] ap_axis_oarg_59_tkeep,
    input [M_AXIS_OARG_59_WIDTH/8-1:0] ap_axis_oarg_59_tstrb,
    input [M_AXIS_OARG_59_WIDTH-1:0] ap_axis_oarg_59_tdata,
    output ap_axis_oarg_59_tready,
    //output AXIS to AXI-Stream interface 60
    input m_axis_oarg_60_aclk,
    input m_axis_oarg_60_aresetn,
    output m_axis_oarg_60_tlast,
    output m_axis_oarg_60_tvalid,
    output [M_AXIS_OARG_60_DMWIDTH/8-1:0] m_axis_oarg_60_tkeep,
    output [M_AXIS_OARG_60_DMWIDTH/8-1:0] m_axis_oarg_60_tstrb,
    output [M_AXIS_OARG_60_DMWIDTH-1:0] m_axis_oarg_60_tdata,
    input m_axis_oarg_60_tready,
    input ap_axis_oarg_60_tlast,
    input ap_axis_oarg_60_tvalid,
    input [M_AXIS_OARG_60_WIDTH/8-1:0] ap_axis_oarg_60_tkeep,
    input [M_AXIS_OARG_60_WIDTH/8-1:0] ap_axis_oarg_60_tstrb,
    input [M_AXIS_OARG_60_WIDTH-1:0] ap_axis_oarg_60_tdata,
    output ap_axis_oarg_60_tready,
    //output AXIS to AXI-Stream interface 61
    input m_axis_oarg_61_aclk,
    input m_axis_oarg_61_aresetn,
    output m_axis_oarg_61_tlast,
    output m_axis_oarg_61_tvalid,
    output [M_AXIS_OARG_61_DMWIDTH/8-1:0] m_axis_oarg_61_tkeep,
    output [M_AXIS_OARG_61_DMWIDTH/8-1:0] m_axis_oarg_61_tstrb,
    output [M_AXIS_OARG_61_DMWIDTH-1:0] m_axis_oarg_61_tdata,
    input m_axis_oarg_61_tready,
    input ap_axis_oarg_61_tlast,
    input ap_axis_oarg_61_tvalid,
    input [M_AXIS_OARG_61_WIDTH/8-1:0] ap_axis_oarg_61_tkeep,
    input [M_AXIS_OARG_61_WIDTH/8-1:0] ap_axis_oarg_61_tstrb,
    input [M_AXIS_OARG_61_WIDTH-1:0] ap_axis_oarg_61_tdata,
    output ap_axis_oarg_61_tready,
    //output AXIS to AXI-Stream interface 62
    input m_axis_oarg_62_aclk,
    input m_axis_oarg_62_aresetn,
    output m_axis_oarg_62_tlast,
    output m_axis_oarg_62_tvalid,
    output [M_AXIS_OARG_62_DMWIDTH/8-1:0] m_axis_oarg_62_tkeep,
    output [M_AXIS_OARG_62_DMWIDTH/8-1:0] m_axis_oarg_62_tstrb,
    output [M_AXIS_OARG_62_DMWIDTH-1:0] m_axis_oarg_62_tdata,
    input m_axis_oarg_62_tready,
    input ap_axis_oarg_62_tlast,
    input ap_axis_oarg_62_tvalid,
    input [M_AXIS_OARG_62_WIDTH/8-1:0] ap_axis_oarg_62_tkeep,
    input [M_AXIS_OARG_62_WIDTH/8-1:0] ap_axis_oarg_62_tstrb,
    input [M_AXIS_OARG_62_WIDTH-1:0] ap_axis_oarg_62_tdata,
    output ap_axis_oarg_62_tready,
    //output AXIS to AXI-Stream interface 63
    input m_axis_oarg_63_aclk,
    input m_axis_oarg_63_aresetn,
    output m_axis_oarg_63_tlast,
    output m_axis_oarg_63_tvalid,
    output [M_AXIS_OARG_63_DMWIDTH/8-1:0] m_axis_oarg_63_tkeep,
    output [M_AXIS_OARG_63_DMWIDTH/8-1:0] m_axis_oarg_63_tstrb,
    output [M_AXIS_OARG_63_DMWIDTH-1:0] m_axis_oarg_63_tdata,
    input m_axis_oarg_63_tready,
    input ap_axis_oarg_63_tlast,
    input ap_axis_oarg_63_tvalid,
    input [M_AXIS_OARG_63_WIDTH/8-1:0] ap_axis_oarg_63_tkeep,
    input [M_AXIS_OARG_63_WIDTH/8-1:0] ap_axis_oarg_63_tstrb,
    input [M_AXIS_OARG_63_WIDTH-1:0] ap_axis_oarg_63_tdata,
    output ap_axis_oarg_63_tready,
    //output AXIS to AXI-Stream interface 64
    input m_axis_oarg_64_aclk,
    input m_axis_oarg_64_aresetn,
    output m_axis_oarg_64_tlast,
    output m_axis_oarg_64_tvalid,
    output [M_AXIS_OARG_64_DMWIDTH/8-1:0] m_axis_oarg_64_tkeep,
    output [M_AXIS_OARG_64_DMWIDTH/8-1:0] m_axis_oarg_64_tstrb,
    output [M_AXIS_OARG_64_DMWIDTH-1:0] m_axis_oarg_64_tdata,
    input m_axis_oarg_64_tready,
    input ap_axis_oarg_64_tlast,
    input ap_axis_oarg_64_tvalid,
    input [M_AXIS_OARG_64_WIDTH/8-1:0] ap_axis_oarg_64_tkeep,
    input [M_AXIS_OARG_64_WIDTH/8-1:0] ap_axis_oarg_64_tstrb,
    input [M_AXIS_OARG_64_WIDTH-1:0] ap_axis_oarg_64_tdata,
    output ap_axis_oarg_64_tready,
    //output AXIS to AXI-Stream interface 65
    input m_axis_oarg_65_aclk,
    input m_axis_oarg_65_aresetn,
    output m_axis_oarg_65_tlast,
    output m_axis_oarg_65_tvalid,
    output [M_AXIS_OARG_65_DMWIDTH/8-1:0] m_axis_oarg_65_tkeep,
    output [M_AXIS_OARG_65_DMWIDTH/8-1:0] m_axis_oarg_65_tstrb,
    output [M_AXIS_OARG_65_DMWIDTH-1:0] m_axis_oarg_65_tdata,
    input m_axis_oarg_65_tready,
    input ap_axis_oarg_65_tlast,
    input ap_axis_oarg_65_tvalid,
    input [M_AXIS_OARG_65_WIDTH/8-1:0] ap_axis_oarg_65_tkeep,
    input [M_AXIS_OARG_65_WIDTH/8-1:0] ap_axis_oarg_65_tstrb,
    input [M_AXIS_OARG_65_WIDTH-1:0] ap_axis_oarg_65_tdata,
    output ap_axis_oarg_65_tready,
    //output AXIS to AXI-Stream interface 66
    input m_axis_oarg_66_aclk,
    input m_axis_oarg_66_aresetn,
    output m_axis_oarg_66_tlast,
    output m_axis_oarg_66_tvalid,
    output [M_AXIS_OARG_66_DMWIDTH/8-1:0] m_axis_oarg_66_tkeep,
    output [M_AXIS_OARG_66_DMWIDTH/8-1:0] m_axis_oarg_66_tstrb,
    output [M_AXIS_OARG_66_DMWIDTH-1:0] m_axis_oarg_66_tdata,
    input m_axis_oarg_66_tready,
    input ap_axis_oarg_66_tlast,
    input ap_axis_oarg_66_tvalid,
    input [M_AXIS_OARG_66_WIDTH/8-1:0] ap_axis_oarg_66_tkeep,
    input [M_AXIS_OARG_66_WIDTH/8-1:0] ap_axis_oarg_66_tstrb,
    input [M_AXIS_OARG_66_WIDTH-1:0] ap_axis_oarg_66_tdata,
    output ap_axis_oarg_66_tready,
    //output AXIS to AXI-Stream interface 67
    input m_axis_oarg_67_aclk,
    input m_axis_oarg_67_aresetn,
    output m_axis_oarg_67_tlast,
    output m_axis_oarg_67_tvalid,
    output [M_AXIS_OARG_67_DMWIDTH/8-1:0] m_axis_oarg_67_tkeep,
    output [M_AXIS_OARG_67_DMWIDTH/8-1:0] m_axis_oarg_67_tstrb,
    output [M_AXIS_OARG_67_DMWIDTH-1:0] m_axis_oarg_67_tdata,
    input m_axis_oarg_67_tready,
    input ap_axis_oarg_67_tlast,
    input ap_axis_oarg_67_tvalid,
    input [M_AXIS_OARG_67_WIDTH/8-1:0] ap_axis_oarg_67_tkeep,
    input [M_AXIS_OARG_67_WIDTH/8-1:0] ap_axis_oarg_67_tstrb,
    input [M_AXIS_OARG_67_WIDTH-1:0] ap_axis_oarg_67_tdata,
    output ap_axis_oarg_67_tready,
    //output AXIS to AXI-Stream interface 68
    input m_axis_oarg_68_aclk,
    input m_axis_oarg_68_aresetn,
    output m_axis_oarg_68_tlast,
    output m_axis_oarg_68_tvalid,
    output [M_AXIS_OARG_68_DMWIDTH/8-1:0] m_axis_oarg_68_tkeep,
    output [M_AXIS_OARG_68_DMWIDTH/8-1:0] m_axis_oarg_68_tstrb,
    output [M_AXIS_OARG_68_DMWIDTH-1:0] m_axis_oarg_68_tdata,
    input m_axis_oarg_68_tready,
    input ap_axis_oarg_68_tlast,
    input ap_axis_oarg_68_tvalid,
    input [M_AXIS_OARG_68_WIDTH/8-1:0] ap_axis_oarg_68_tkeep,
    input [M_AXIS_OARG_68_WIDTH/8-1:0] ap_axis_oarg_68_tstrb,
    input [M_AXIS_OARG_68_WIDTH-1:0] ap_axis_oarg_68_tdata,
    output ap_axis_oarg_68_tready,
    //output AXIS to AXI-Stream interface 69
    input m_axis_oarg_69_aclk,
    input m_axis_oarg_69_aresetn,
    output m_axis_oarg_69_tlast,
    output m_axis_oarg_69_tvalid,
    output [M_AXIS_OARG_69_DMWIDTH/8-1:0] m_axis_oarg_69_tkeep,
    output [M_AXIS_OARG_69_DMWIDTH/8-1:0] m_axis_oarg_69_tstrb,
    output [M_AXIS_OARG_69_DMWIDTH-1:0] m_axis_oarg_69_tdata,
    input m_axis_oarg_69_tready,
    input ap_axis_oarg_69_tlast,
    input ap_axis_oarg_69_tvalid,
    input [M_AXIS_OARG_69_WIDTH/8-1:0] ap_axis_oarg_69_tkeep,
    input [M_AXIS_OARG_69_WIDTH/8-1:0] ap_axis_oarg_69_tstrb,
    input [M_AXIS_OARG_69_WIDTH-1:0] ap_axis_oarg_69_tdata,
    output ap_axis_oarg_69_tready,
    //output AXIS to AXI-Stream interface 70
    input m_axis_oarg_70_aclk,
    input m_axis_oarg_70_aresetn,
    output m_axis_oarg_70_tlast,
    output m_axis_oarg_70_tvalid,
    output [M_AXIS_OARG_70_DMWIDTH/8-1:0] m_axis_oarg_70_tkeep,
    output [M_AXIS_OARG_70_DMWIDTH/8-1:0] m_axis_oarg_70_tstrb,
    output [M_AXIS_OARG_70_DMWIDTH-1:0] m_axis_oarg_70_tdata,
    input m_axis_oarg_70_tready,
    input ap_axis_oarg_70_tlast,
    input ap_axis_oarg_70_tvalid,
    input [M_AXIS_OARG_70_WIDTH/8-1:0] ap_axis_oarg_70_tkeep,
    input [M_AXIS_OARG_70_WIDTH/8-1:0] ap_axis_oarg_70_tstrb,
    input [M_AXIS_OARG_70_WIDTH-1:0] ap_axis_oarg_70_tdata,
    output ap_axis_oarg_70_tready,
    //output AXIS to AXI-Stream interface 71
    input m_axis_oarg_71_aclk,
    input m_axis_oarg_71_aresetn,
    output m_axis_oarg_71_tlast,
    output m_axis_oarg_71_tvalid,
    output [M_AXIS_OARG_71_DMWIDTH/8-1:0] m_axis_oarg_71_tkeep,
    output [M_AXIS_OARG_71_DMWIDTH/8-1:0] m_axis_oarg_71_tstrb,
    output [M_AXIS_OARG_71_DMWIDTH-1:0] m_axis_oarg_71_tdata,
    input m_axis_oarg_71_tready,
    input ap_axis_oarg_71_tlast,
    input ap_axis_oarg_71_tvalid,
    input [M_AXIS_OARG_71_WIDTH/8-1:0] ap_axis_oarg_71_tkeep,
    input [M_AXIS_OARG_71_WIDTH/8-1:0] ap_axis_oarg_71_tstrb,
    input [M_AXIS_OARG_71_WIDTH-1:0] ap_axis_oarg_71_tdata,
    output ap_axis_oarg_71_tready,
    //output AXIS to AXI-Stream interface 72
    input m_axis_oarg_72_aclk,
    input m_axis_oarg_72_aresetn,
    output m_axis_oarg_72_tlast,
    output m_axis_oarg_72_tvalid,
    output [M_AXIS_OARG_72_DMWIDTH/8-1:0] m_axis_oarg_72_tkeep,
    output [M_AXIS_OARG_72_DMWIDTH/8-1:0] m_axis_oarg_72_tstrb,
    output [M_AXIS_OARG_72_DMWIDTH-1:0] m_axis_oarg_72_tdata,
    input m_axis_oarg_72_tready,
    input ap_axis_oarg_72_tlast,
    input ap_axis_oarg_72_tvalid,
    input [M_AXIS_OARG_72_WIDTH/8-1:0] ap_axis_oarg_72_tkeep,
    input [M_AXIS_OARG_72_WIDTH/8-1:0] ap_axis_oarg_72_tstrb,
    input [M_AXIS_OARG_72_WIDTH-1:0] ap_axis_oarg_72_tdata,
    output ap_axis_oarg_72_tready,
    //output AXIS to AXI-Stream interface 73
    input m_axis_oarg_73_aclk,
    input m_axis_oarg_73_aresetn,
    output m_axis_oarg_73_tlast,
    output m_axis_oarg_73_tvalid,
    output [M_AXIS_OARG_73_DMWIDTH/8-1:0] m_axis_oarg_73_tkeep,
    output [M_AXIS_OARG_73_DMWIDTH/8-1:0] m_axis_oarg_73_tstrb,
    output [M_AXIS_OARG_73_DMWIDTH-1:0] m_axis_oarg_73_tdata,
    input m_axis_oarg_73_tready,
    input ap_axis_oarg_73_tlast,
    input ap_axis_oarg_73_tvalid,
    input [M_AXIS_OARG_73_WIDTH/8-1:0] ap_axis_oarg_73_tkeep,
    input [M_AXIS_OARG_73_WIDTH/8-1:0] ap_axis_oarg_73_tstrb,
    input [M_AXIS_OARG_73_WIDTH-1:0] ap_axis_oarg_73_tdata,
    output ap_axis_oarg_73_tready,
    //output AXIS to AXI-Stream interface 74
    input m_axis_oarg_74_aclk,
    input m_axis_oarg_74_aresetn,
    output m_axis_oarg_74_tlast,
    output m_axis_oarg_74_tvalid,
    output [M_AXIS_OARG_74_DMWIDTH/8-1:0] m_axis_oarg_74_tkeep,
    output [M_AXIS_OARG_74_DMWIDTH/8-1:0] m_axis_oarg_74_tstrb,
    output [M_AXIS_OARG_74_DMWIDTH-1:0] m_axis_oarg_74_tdata,
    input m_axis_oarg_74_tready,
    input ap_axis_oarg_74_tlast,
    input ap_axis_oarg_74_tvalid,
    input [M_AXIS_OARG_74_WIDTH/8-1:0] ap_axis_oarg_74_tkeep,
    input [M_AXIS_OARG_74_WIDTH/8-1:0] ap_axis_oarg_74_tstrb,
    input [M_AXIS_OARG_74_WIDTH-1:0] ap_axis_oarg_74_tdata,
    output ap_axis_oarg_74_tready,
    //output AXIS to AXI-Stream interface 75
    input m_axis_oarg_75_aclk,
    input m_axis_oarg_75_aresetn,
    output m_axis_oarg_75_tlast,
    output m_axis_oarg_75_tvalid,
    output [M_AXIS_OARG_75_DMWIDTH/8-1:0] m_axis_oarg_75_tkeep,
    output [M_AXIS_OARG_75_DMWIDTH/8-1:0] m_axis_oarg_75_tstrb,
    output [M_AXIS_OARG_75_DMWIDTH-1:0] m_axis_oarg_75_tdata,
    input m_axis_oarg_75_tready,
    input ap_axis_oarg_75_tlast,
    input ap_axis_oarg_75_tvalid,
    input [M_AXIS_OARG_75_WIDTH/8-1:0] ap_axis_oarg_75_tkeep,
    input [M_AXIS_OARG_75_WIDTH/8-1:0] ap_axis_oarg_75_tstrb,
    input [M_AXIS_OARG_75_WIDTH-1:0] ap_axis_oarg_75_tdata,
    output ap_axis_oarg_75_tready,
    //output AXIS to AXI-Stream interface 76
    input m_axis_oarg_76_aclk,
    input m_axis_oarg_76_aresetn,
    output m_axis_oarg_76_tlast,
    output m_axis_oarg_76_tvalid,
    output [M_AXIS_OARG_76_DMWIDTH/8-1:0] m_axis_oarg_76_tkeep,
    output [M_AXIS_OARG_76_DMWIDTH/8-1:0] m_axis_oarg_76_tstrb,
    output [M_AXIS_OARG_76_DMWIDTH-1:0] m_axis_oarg_76_tdata,
    input m_axis_oarg_76_tready,
    input ap_axis_oarg_76_tlast,
    input ap_axis_oarg_76_tvalid,
    input [M_AXIS_OARG_76_WIDTH/8-1:0] ap_axis_oarg_76_tkeep,
    input [M_AXIS_OARG_76_WIDTH/8-1:0] ap_axis_oarg_76_tstrb,
    input [M_AXIS_OARG_76_WIDTH-1:0] ap_axis_oarg_76_tdata,
    output ap_axis_oarg_76_tready,
    //output AXIS to AXI-Stream interface 77
    input m_axis_oarg_77_aclk,
    input m_axis_oarg_77_aresetn,
    output m_axis_oarg_77_tlast,
    output m_axis_oarg_77_tvalid,
    output [M_AXIS_OARG_77_DMWIDTH/8-1:0] m_axis_oarg_77_tkeep,
    output [M_AXIS_OARG_77_DMWIDTH/8-1:0] m_axis_oarg_77_tstrb,
    output [M_AXIS_OARG_77_DMWIDTH-1:0] m_axis_oarg_77_tdata,
    input m_axis_oarg_77_tready,
    input ap_axis_oarg_77_tlast,
    input ap_axis_oarg_77_tvalid,
    input [M_AXIS_OARG_77_WIDTH/8-1:0] ap_axis_oarg_77_tkeep,
    input [M_AXIS_OARG_77_WIDTH/8-1:0] ap_axis_oarg_77_tstrb,
    input [M_AXIS_OARG_77_WIDTH-1:0] ap_axis_oarg_77_tdata,
    output ap_axis_oarg_77_tready,
    //output AXIS to AXI-Stream interface 78
    input m_axis_oarg_78_aclk,
    input m_axis_oarg_78_aresetn,
    output m_axis_oarg_78_tlast,
    output m_axis_oarg_78_tvalid,
    output [M_AXIS_OARG_78_DMWIDTH/8-1:0] m_axis_oarg_78_tkeep,
    output [M_AXIS_OARG_78_DMWIDTH/8-1:0] m_axis_oarg_78_tstrb,
    output [M_AXIS_OARG_78_DMWIDTH-1:0] m_axis_oarg_78_tdata,
    input m_axis_oarg_78_tready,
    input ap_axis_oarg_78_tlast,
    input ap_axis_oarg_78_tvalid,
    input [M_AXIS_OARG_78_WIDTH/8-1:0] ap_axis_oarg_78_tkeep,
    input [M_AXIS_OARG_78_WIDTH/8-1:0] ap_axis_oarg_78_tstrb,
    input [M_AXIS_OARG_78_WIDTH-1:0] ap_axis_oarg_78_tdata,
    output ap_axis_oarg_78_tready,
    //output AXIS to AXI-Stream interface 79
    input m_axis_oarg_79_aclk,
    input m_axis_oarg_79_aresetn,
    output m_axis_oarg_79_tlast,
    output m_axis_oarg_79_tvalid,
    output [M_AXIS_OARG_79_DMWIDTH/8-1:0] m_axis_oarg_79_tkeep,
    output [M_AXIS_OARG_79_DMWIDTH/8-1:0] m_axis_oarg_79_tstrb,
    output [M_AXIS_OARG_79_DMWIDTH-1:0] m_axis_oarg_79_tdata,
    input m_axis_oarg_79_tready,
    input ap_axis_oarg_79_tlast,
    input ap_axis_oarg_79_tvalid,
    input [M_AXIS_OARG_79_WIDTH/8-1:0] ap_axis_oarg_79_tkeep,
    input [M_AXIS_OARG_79_WIDTH/8-1:0] ap_axis_oarg_79_tstrb,
    input [M_AXIS_OARG_79_WIDTH-1:0] ap_axis_oarg_79_tdata,
    output ap_axis_oarg_79_tready,
    //output AXIS to AXI-Stream interface 80
    input m_axis_oarg_80_aclk,
    input m_axis_oarg_80_aresetn,
    output m_axis_oarg_80_tlast,
    output m_axis_oarg_80_tvalid,
    output [M_AXIS_OARG_80_DMWIDTH/8-1:0] m_axis_oarg_80_tkeep,
    output [M_AXIS_OARG_80_DMWIDTH/8-1:0] m_axis_oarg_80_tstrb,
    output [M_AXIS_OARG_80_DMWIDTH-1:0] m_axis_oarg_80_tdata,
    input m_axis_oarg_80_tready,
    input ap_axis_oarg_80_tlast,
    input ap_axis_oarg_80_tvalid,
    input [M_AXIS_OARG_80_WIDTH/8-1:0] ap_axis_oarg_80_tkeep,
    input [M_AXIS_OARG_80_WIDTH/8-1:0] ap_axis_oarg_80_tstrb,
    input [M_AXIS_OARG_80_WIDTH-1:0] ap_axis_oarg_80_tdata,
    output ap_axis_oarg_80_tready,
    //output AXIS to AXI-Stream interface 81
    input m_axis_oarg_81_aclk,
    input m_axis_oarg_81_aresetn,
    output m_axis_oarg_81_tlast,
    output m_axis_oarg_81_tvalid,
    output [M_AXIS_OARG_81_DMWIDTH/8-1:0] m_axis_oarg_81_tkeep,
    output [M_AXIS_OARG_81_DMWIDTH/8-1:0] m_axis_oarg_81_tstrb,
    output [M_AXIS_OARG_81_DMWIDTH-1:0] m_axis_oarg_81_tdata,
    input m_axis_oarg_81_tready,
    input ap_axis_oarg_81_tlast,
    input ap_axis_oarg_81_tvalid,
    input [M_AXIS_OARG_81_WIDTH/8-1:0] ap_axis_oarg_81_tkeep,
    input [M_AXIS_OARG_81_WIDTH/8-1:0] ap_axis_oarg_81_tstrb,
    input [M_AXIS_OARG_81_WIDTH-1:0] ap_axis_oarg_81_tdata,
    output ap_axis_oarg_81_tready,
    //output AXIS to AXI-Stream interface 82
    input m_axis_oarg_82_aclk,
    input m_axis_oarg_82_aresetn,
    output m_axis_oarg_82_tlast,
    output m_axis_oarg_82_tvalid,
    output [M_AXIS_OARG_82_DMWIDTH/8-1:0] m_axis_oarg_82_tkeep,
    output [M_AXIS_OARG_82_DMWIDTH/8-1:0] m_axis_oarg_82_tstrb,
    output [M_AXIS_OARG_82_DMWIDTH-1:0] m_axis_oarg_82_tdata,
    input m_axis_oarg_82_tready,
    input ap_axis_oarg_82_tlast,
    input ap_axis_oarg_82_tvalid,
    input [M_AXIS_OARG_82_WIDTH/8-1:0] ap_axis_oarg_82_tkeep,
    input [M_AXIS_OARG_82_WIDTH/8-1:0] ap_axis_oarg_82_tstrb,
    input [M_AXIS_OARG_82_WIDTH-1:0] ap_axis_oarg_82_tdata,
    output ap_axis_oarg_82_tready,
    //output AXIS to AXI-Stream interface 83
    input m_axis_oarg_83_aclk,
    input m_axis_oarg_83_aresetn,
    output m_axis_oarg_83_tlast,
    output m_axis_oarg_83_tvalid,
    output [M_AXIS_OARG_83_DMWIDTH/8-1:0] m_axis_oarg_83_tkeep,
    output [M_AXIS_OARG_83_DMWIDTH/8-1:0] m_axis_oarg_83_tstrb,
    output [M_AXIS_OARG_83_DMWIDTH-1:0] m_axis_oarg_83_tdata,
    input m_axis_oarg_83_tready,
    input ap_axis_oarg_83_tlast,
    input ap_axis_oarg_83_tvalid,
    input [M_AXIS_OARG_83_WIDTH/8-1:0] ap_axis_oarg_83_tkeep,
    input [M_AXIS_OARG_83_WIDTH/8-1:0] ap_axis_oarg_83_tstrb,
    input [M_AXIS_OARG_83_WIDTH-1:0] ap_axis_oarg_83_tdata,
    output ap_axis_oarg_83_tready,
    //output AXIS to AXI-Stream interface 84
    input m_axis_oarg_84_aclk,
    input m_axis_oarg_84_aresetn,
    output m_axis_oarg_84_tlast,
    output m_axis_oarg_84_tvalid,
    output [M_AXIS_OARG_84_DMWIDTH/8-1:0] m_axis_oarg_84_tkeep,
    output [M_AXIS_OARG_84_DMWIDTH/8-1:0] m_axis_oarg_84_tstrb,
    output [M_AXIS_OARG_84_DMWIDTH-1:0] m_axis_oarg_84_tdata,
    input m_axis_oarg_84_tready,
    input ap_axis_oarg_84_tlast,
    input ap_axis_oarg_84_tvalid,
    input [M_AXIS_OARG_84_WIDTH/8-1:0] ap_axis_oarg_84_tkeep,
    input [M_AXIS_OARG_84_WIDTH/8-1:0] ap_axis_oarg_84_tstrb,
    input [M_AXIS_OARG_84_WIDTH-1:0] ap_axis_oarg_84_tdata,
    output ap_axis_oarg_84_tready,
    //output AXIS to AXI-Stream interface 85
    input m_axis_oarg_85_aclk,
    input m_axis_oarg_85_aresetn,
    output m_axis_oarg_85_tlast,
    output m_axis_oarg_85_tvalid,
    output [M_AXIS_OARG_85_DMWIDTH/8-1:0] m_axis_oarg_85_tkeep,
    output [M_AXIS_OARG_85_DMWIDTH/8-1:0] m_axis_oarg_85_tstrb,
    output [M_AXIS_OARG_85_DMWIDTH-1:0] m_axis_oarg_85_tdata,
    input m_axis_oarg_85_tready,
    input ap_axis_oarg_85_tlast,
    input ap_axis_oarg_85_tvalid,
    input [M_AXIS_OARG_85_WIDTH/8-1:0] ap_axis_oarg_85_tkeep,
    input [M_AXIS_OARG_85_WIDTH/8-1:0] ap_axis_oarg_85_tstrb,
    input [M_AXIS_OARG_85_WIDTH-1:0] ap_axis_oarg_85_tdata,
    output ap_axis_oarg_85_tready,
    //output AXIS to AXI-Stream interface 86
    input m_axis_oarg_86_aclk,
    input m_axis_oarg_86_aresetn,
    output m_axis_oarg_86_tlast,
    output m_axis_oarg_86_tvalid,
    output [M_AXIS_OARG_86_DMWIDTH/8-1:0] m_axis_oarg_86_tkeep,
    output [M_AXIS_OARG_86_DMWIDTH/8-1:0] m_axis_oarg_86_tstrb,
    output [M_AXIS_OARG_86_DMWIDTH-1:0] m_axis_oarg_86_tdata,
    input m_axis_oarg_86_tready,
    input ap_axis_oarg_86_tlast,
    input ap_axis_oarg_86_tvalid,
    input [M_AXIS_OARG_86_WIDTH/8-1:0] ap_axis_oarg_86_tkeep,
    input [M_AXIS_OARG_86_WIDTH/8-1:0] ap_axis_oarg_86_tstrb,
    input [M_AXIS_OARG_86_WIDTH-1:0] ap_axis_oarg_86_tdata,
    output ap_axis_oarg_86_tready,
    //output AXIS to AXI-Stream interface 87
    input m_axis_oarg_87_aclk,
    input m_axis_oarg_87_aresetn,
    output m_axis_oarg_87_tlast,
    output m_axis_oarg_87_tvalid,
    output [M_AXIS_OARG_87_DMWIDTH/8-1:0] m_axis_oarg_87_tkeep,
    output [M_AXIS_OARG_87_DMWIDTH/8-1:0] m_axis_oarg_87_tstrb,
    output [M_AXIS_OARG_87_DMWIDTH-1:0] m_axis_oarg_87_tdata,
    input m_axis_oarg_87_tready,
    input ap_axis_oarg_87_tlast,
    input ap_axis_oarg_87_tvalid,
    input [M_AXIS_OARG_87_WIDTH/8-1:0] ap_axis_oarg_87_tkeep,
    input [M_AXIS_OARG_87_WIDTH/8-1:0] ap_axis_oarg_87_tstrb,
    input [M_AXIS_OARG_87_WIDTH-1:0] ap_axis_oarg_87_tdata,
    output ap_axis_oarg_87_tready,
    //output AXIS to AXI-Stream interface 88
    input m_axis_oarg_88_aclk,
    input m_axis_oarg_88_aresetn,
    output m_axis_oarg_88_tlast,
    output m_axis_oarg_88_tvalid,
    output [M_AXIS_OARG_88_DMWIDTH/8-1:0] m_axis_oarg_88_tkeep,
    output [M_AXIS_OARG_88_DMWIDTH/8-1:0] m_axis_oarg_88_tstrb,
    output [M_AXIS_OARG_88_DMWIDTH-1:0] m_axis_oarg_88_tdata,
    input m_axis_oarg_88_tready,
    input ap_axis_oarg_88_tlast,
    input ap_axis_oarg_88_tvalid,
    input [M_AXIS_OARG_88_WIDTH/8-1:0] ap_axis_oarg_88_tkeep,
    input [M_AXIS_OARG_88_WIDTH/8-1:0] ap_axis_oarg_88_tstrb,
    input [M_AXIS_OARG_88_WIDTH-1:0] ap_axis_oarg_88_tdata,
    output ap_axis_oarg_88_tready,
    //output AXIS to AXI-Stream interface 89
    input m_axis_oarg_89_aclk,
    input m_axis_oarg_89_aresetn,
    output m_axis_oarg_89_tlast,
    output m_axis_oarg_89_tvalid,
    output [M_AXIS_OARG_89_DMWIDTH/8-1:0] m_axis_oarg_89_tkeep,
    output [M_AXIS_OARG_89_DMWIDTH/8-1:0] m_axis_oarg_89_tstrb,
    output [M_AXIS_OARG_89_DMWIDTH-1:0] m_axis_oarg_89_tdata,
    input m_axis_oarg_89_tready,
    input ap_axis_oarg_89_tlast,
    input ap_axis_oarg_89_tvalid,
    input [M_AXIS_OARG_89_WIDTH/8-1:0] ap_axis_oarg_89_tkeep,
    input [M_AXIS_OARG_89_WIDTH/8-1:0] ap_axis_oarg_89_tstrb,
    input [M_AXIS_OARG_89_WIDTH-1:0] ap_axis_oarg_89_tdata,
    output ap_axis_oarg_89_tready,
    //output AXIS to AXI-Stream interface 90
    input m_axis_oarg_90_aclk,
    input m_axis_oarg_90_aresetn,
    output m_axis_oarg_90_tlast,
    output m_axis_oarg_90_tvalid,
    output [M_AXIS_OARG_90_DMWIDTH/8-1:0] m_axis_oarg_90_tkeep,
    output [M_AXIS_OARG_90_DMWIDTH/8-1:0] m_axis_oarg_90_tstrb,
    output [M_AXIS_OARG_90_DMWIDTH-1:0] m_axis_oarg_90_tdata,
    input m_axis_oarg_90_tready,
    input ap_axis_oarg_90_tlast,
    input ap_axis_oarg_90_tvalid,
    input [M_AXIS_OARG_90_WIDTH/8-1:0] ap_axis_oarg_90_tkeep,
    input [M_AXIS_OARG_90_WIDTH/8-1:0] ap_axis_oarg_90_tstrb,
    input [M_AXIS_OARG_90_WIDTH-1:0] ap_axis_oarg_90_tdata,
    output ap_axis_oarg_90_tready,
    //output AXIS to AXI-Stream interface 91
    input m_axis_oarg_91_aclk,
    input m_axis_oarg_91_aresetn,
    output m_axis_oarg_91_tlast,
    output m_axis_oarg_91_tvalid,
    output [M_AXIS_OARG_91_DMWIDTH/8-1:0] m_axis_oarg_91_tkeep,
    output [M_AXIS_OARG_91_DMWIDTH/8-1:0] m_axis_oarg_91_tstrb,
    output [M_AXIS_OARG_91_DMWIDTH-1:0] m_axis_oarg_91_tdata,
    input m_axis_oarg_91_tready,
    input ap_axis_oarg_91_tlast,
    input ap_axis_oarg_91_tvalid,
    input [M_AXIS_OARG_91_WIDTH/8-1:0] ap_axis_oarg_91_tkeep,
    input [M_AXIS_OARG_91_WIDTH/8-1:0] ap_axis_oarg_91_tstrb,
    input [M_AXIS_OARG_91_WIDTH-1:0] ap_axis_oarg_91_tdata,
    output ap_axis_oarg_91_tready,
    //output AXIS to AXI-Stream interface 92
    input m_axis_oarg_92_aclk,
    input m_axis_oarg_92_aresetn,
    output m_axis_oarg_92_tlast,
    output m_axis_oarg_92_tvalid,
    output [M_AXIS_OARG_92_DMWIDTH/8-1:0] m_axis_oarg_92_tkeep,
    output [M_AXIS_OARG_92_DMWIDTH/8-1:0] m_axis_oarg_92_tstrb,
    output [M_AXIS_OARG_92_DMWIDTH-1:0] m_axis_oarg_92_tdata,
    input m_axis_oarg_92_tready,
    input ap_axis_oarg_92_tlast,
    input ap_axis_oarg_92_tvalid,
    input [M_AXIS_OARG_92_WIDTH/8-1:0] ap_axis_oarg_92_tkeep,
    input [M_AXIS_OARG_92_WIDTH/8-1:0] ap_axis_oarg_92_tstrb,
    input [M_AXIS_OARG_92_WIDTH-1:0] ap_axis_oarg_92_tdata,
    output ap_axis_oarg_92_tready,
    //output AXIS to AXI-Stream interface 93
    input m_axis_oarg_93_aclk,
    input m_axis_oarg_93_aresetn,
    output m_axis_oarg_93_tlast,
    output m_axis_oarg_93_tvalid,
    output [M_AXIS_OARG_93_DMWIDTH/8-1:0] m_axis_oarg_93_tkeep,
    output [M_AXIS_OARG_93_DMWIDTH/8-1:0] m_axis_oarg_93_tstrb,
    output [M_AXIS_OARG_93_DMWIDTH-1:0] m_axis_oarg_93_tdata,
    input m_axis_oarg_93_tready,
    input ap_axis_oarg_93_tlast,
    input ap_axis_oarg_93_tvalid,
    input [M_AXIS_OARG_93_WIDTH/8-1:0] ap_axis_oarg_93_tkeep,
    input [M_AXIS_OARG_93_WIDTH/8-1:0] ap_axis_oarg_93_tstrb,
    input [M_AXIS_OARG_93_WIDTH-1:0] ap_axis_oarg_93_tdata,
    output ap_axis_oarg_93_tready,
    //output AXIS to AXI-Stream interface 94
    input m_axis_oarg_94_aclk,
    input m_axis_oarg_94_aresetn,
    output m_axis_oarg_94_tlast,
    output m_axis_oarg_94_tvalid,
    output [M_AXIS_OARG_94_DMWIDTH/8-1:0] m_axis_oarg_94_tkeep,
    output [M_AXIS_OARG_94_DMWIDTH/8-1:0] m_axis_oarg_94_tstrb,
    output [M_AXIS_OARG_94_DMWIDTH-1:0] m_axis_oarg_94_tdata,
    input m_axis_oarg_94_tready,
    input ap_axis_oarg_94_tlast,
    input ap_axis_oarg_94_tvalid,
    input [M_AXIS_OARG_94_WIDTH/8-1:0] ap_axis_oarg_94_tkeep,
    input [M_AXIS_OARG_94_WIDTH/8-1:0] ap_axis_oarg_94_tstrb,
    input [M_AXIS_OARG_94_WIDTH-1:0] ap_axis_oarg_94_tdata,
    output ap_axis_oarg_94_tready,
    //output AXIS to AXI-Stream interface 95
    input m_axis_oarg_95_aclk,
    input m_axis_oarg_95_aresetn,
    output m_axis_oarg_95_tlast,
    output m_axis_oarg_95_tvalid,
    output [M_AXIS_OARG_95_DMWIDTH/8-1:0] m_axis_oarg_95_tkeep,
    output [M_AXIS_OARG_95_DMWIDTH/8-1:0] m_axis_oarg_95_tstrb,
    output [M_AXIS_OARG_95_DMWIDTH-1:0] m_axis_oarg_95_tdata,
    input m_axis_oarg_95_tready,
    input ap_axis_oarg_95_tlast,
    input ap_axis_oarg_95_tvalid,
    input [M_AXIS_OARG_95_WIDTH/8-1:0] ap_axis_oarg_95_tkeep,
    input [M_AXIS_OARG_95_WIDTH/8-1:0] ap_axis_oarg_95_tstrb,
    input [M_AXIS_OARG_95_WIDTH-1:0] ap_axis_oarg_95_tdata,
    output ap_axis_oarg_95_tready,
    //output AXIS to AXI-Stream interface 96
    input m_axis_oarg_96_aclk,
    input m_axis_oarg_96_aresetn,
    output m_axis_oarg_96_tlast,
    output m_axis_oarg_96_tvalid,
    output [M_AXIS_OARG_96_DMWIDTH/8-1:0] m_axis_oarg_96_tkeep,
    output [M_AXIS_OARG_96_DMWIDTH/8-1:0] m_axis_oarg_96_tstrb,
    output [M_AXIS_OARG_96_DMWIDTH-1:0] m_axis_oarg_96_tdata,
    input m_axis_oarg_96_tready,
    input ap_axis_oarg_96_tlast,
    input ap_axis_oarg_96_tvalid,
    input [M_AXIS_OARG_96_WIDTH/8-1:0] ap_axis_oarg_96_tkeep,
    input [M_AXIS_OARG_96_WIDTH/8-1:0] ap_axis_oarg_96_tstrb,
    input [M_AXIS_OARG_96_WIDTH-1:0] ap_axis_oarg_96_tdata,
    output ap_axis_oarg_96_tready,
    //output AXIS to AXI-Stream interface 97
    input m_axis_oarg_97_aclk,
    input m_axis_oarg_97_aresetn,
    output m_axis_oarg_97_tlast,
    output m_axis_oarg_97_tvalid,
    output [M_AXIS_OARG_97_DMWIDTH/8-1:0] m_axis_oarg_97_tkeep,
    output [M_AXIS_OARG_97_DMWIDTH/8-1:0] m_axis_oarg_97_tstrb,
    output [M_AXIS_OARG_97_DMWIDTH-1:0] m_axis_oarg_97_tdata,
    input m_axis_oarg_97_tready,
    input ap_axis_oarg_97_tlast,
    input ap_axis_oarg_97_tvalid,
    input [M_AXIS_OARG_97_WIDTH/8-1:0] ap_axis_oarg_97_tkeep,
    input [M_AXIS_OARG_97_WIDTH/8-1:0] ap_axis_oarg_97_tstrb,
    input [M_AXIS_OARG_97_WIDTH-1:0] ap_axis_oarg_97_tdata,
    output ap_axis_oarg_97_tready,
    //output AXIS to AXI-Stream interface 98
    input m_axis_oarg_98_aclk,
    input m_axis_oarg_98_aresetn,
    output m_axis_oarg_98_tlast,
    output m_axis_oarg_98_tvalid,
    output [M_AXIS_OARG_98_DMWIDTH/8-1:0] m_axis_oarg_98_tkeep,
    output [M_AXIS_OARG_98_DMWIDTH/8-1:0] m_axis_oarg_98_tstrb,
    output [M_AXIS_OARG_98_DMWIDTH-1:0] m_axis_oarg_98_tdata,
    input m_axis_oarg_98_tready,
    input ap_axis_oarg_98_tlast,
    input ap_axis_oarg_98_tvalid,
    input [M_AXIS_OARG_98_WIDTH/8-1:0] ap_axis_oarg_98_tkeep,
    input [M_AXIS_OARG_98_WIDTH/8-1:0] ap_axis_oarg_98_tstrb,
    input [M_AXIS_OARG_98_WIDTH-1:0] ap_axis_oarg_98_tdata,
    output ap_axis_oarg_98_tready,
    //output AXIS to AXI-Stream interface 99
    input m_axis_oarg_99_aclk,
    input m_axis_oarg_99_aresetn,
    output m_axis_oarg_99_tlast,
    output m_axis_oarg_99_tvalid,
    output [M_AXIS_OARG_99_DMWIDTH/8-1:0] m_axis_oarg_99_tkeep,
    output [M_AXIS_OARG_99_DMWIDTH/8-1:0] m_axis_oarg_99_tstrb,
    output [M_AXIS_OARG_99_DMWIDTH-1:0] m_axis_oarg_99_tdata,
    input m_axis_oarg_99_tready,
    input ap_axis_oarg_99_tlast,
    input ap_axis_oarg_99_tvalid,
    input [M_AXIS_OARG_99_WIDTH/8-1:0] ap_axis_oarg_99_tkeep,
    input [M_AXIS_OARG_99_WIDTH/8-1:0] ap_axis_oarg_99_tstrb,
    input [M_AXIS_OARG_99_WIDTH-1:0] ap_axis_oarg_99_tdata,
    output ap_axis_oarg_99_tready,
    //output AXIS to AXI-Stream interface 100
    input m_axis_oarg_100_aclk,
    input m_axis_oarg_100_aresetn,
    output m_axis_oarg_100_tlast,
    output m_axis_oarg_100_tvalid,
    output [M_AXIS_OARG_100_DMWIDTH/8-1:0] m_axis_oarg_100_tkeep,
    output [M_AXIS_OARG_100_DMWIDTH/8-1:0] m_axis_oarg_100_tstrb,
    output [M_AXIS_OARG_100_DMWIDTH-1:0] m_axis_oarg_100_tdata,
    input m_axis_oarg_100_tready,
    input ap_axis_oarg_100_tlast,
    input ap_axis_oarg_100_tvalid,
    input [M_AXIS_OARG_100_WIDTH/8-1:0] ap_axis_oarg_100_tkeep,
    input [M_AXIS_OARG_100_WIDTH/8-1:0] ap_axis_oarg_100_tstrb,
    input [M_AXIS_OARG_100_WIDTH-1:0] ap_axis_oarg_100_tdata,
    output ap_axis_oarg_100_tready,
    //output AXIS to AXI-Stream interface 101
    input m_axis_oarg_101_aclk,
    input m_axis_oarg_101_aresetn,
    output m_axis_oarg_101_tlast,
    output m_axis_oarg_101_tvalid,
    output [M_AXIS_OARG_101_DMWIDTH/8-1:0] m_axis_oarg_101_tkeep,
    output [M_AXIS_OARG_101_DMWIDTH/8-1:0] m_axis_oarg_101_tstrb,
    output [M_AXIS_OARG_101_DMWIDTH-1:0] m_axis_oarg_101_tdata,
    input m_axis_oarg_101_tready,
    input ap_axis_oarg_101_tlast,
    input ap_axis_oarg_101_tvalid,
    input [M_AXIS_OARG_101_WIDTH/8-1:0] ap_axis_oarg_101_tkeep,
    input [M_AXIS_OARG_101_WIDTH/8-1:0] ap_axis_oarg_101_tstrb,
    input [M_AXIS_OARG_101_WIDTH-1:0] ap_axis_oarg_101_tdata,
    output ap_axis_oarg_101_tready,
    //output AXIS to AXI-Stream interface 102
    input m_axis_oarg_102_aclk,
    input m_axis_oarg_102_aresetn,
    output m_axis_oarg_102_tlast,
    output m_axis_oarg_102_tvalid,
    output [M_AXIS_OARG_102_DMWIDTH/8-1:0] m_axis_oarg_102_tkeep,
    output [M_AXIS_OARG_102_DMWIDTH/8-1:0] m_axis_oarg_102_tstrb,
    output [M_AXIS_OARG_102_DMWIDTH-1:0] m_axis_oarg_102_tdata,
    input m_axis_oarg_102_tready,
    input ap_axis_oarg_102_tlast,
    input ap_axis_oarg_102_tvalid,
    input [M_AXIS_OARG_102_WIDTH/8-1:0] ap_axis_oarg_102_tkeep,
    input [M_AXIS_OARG_102_WIDTH/8-1:0] ap_axis_oarg_102_tstrb,
    input [M_AXIS_OARG_102_WIDTH-1:0] ap_axis_oarg_102_tdata,
    output ap_axis_oarg_102_tready,
    //output AXIS to AXI-Stream interface 103
    input m_axis_oarg_103_aclk,
    input m_axis_oarg_103_aresetn,
    output m_axis_oarg_103_tlast,
    output m_axis_oarg_103_tvalid,
    output [M_AXIS_OARG_103_DMWIDTH/8-1:0] m_axis_oarg_103_tkeep,
    output [M_AXIS_OARG_103_DMWIDTH/8-1:0] m_axis_oarg_103_tstrb,
    output [M_AXIS_OARG_103_DMWIDTH-1:0] m_axis_oarg_103_tdata,
    input m_axis_oarg_103_tready,
    input ap_axis_oarg_103_tlast,
    input ap_axis_oarg_103_tvalid,
    input [M_AXIS_OARG_103_WIDTH/8-1:0] ap_axis_oarg_103_tkeep,
    input [M_AXIS_OARG_103_WIDTH/8-1:0] ap_axis_oarg_103_tstrb,
    input [M_AXIS_OARG_103_WIDTH-1:0] ap_axis_oarg_103_tdata,
    output ap_axis_oarg_103_tready,
    //output AXIS to AXI-Stream interface 104
    input m_axis_oarg_104_aclk,
    input m_axis_oarg_104_aresetn,
    output m_axis_oarg_104_tlast,
    output m_axis_oarg_104_tvalid,
    output [M_AXIS_OARG_104_DMWIDTH/8-1:0] m_axis_oarg_104_tkeep,
    output [M_AXIS_OARG_104_DMWIDTH/8-1:0] m_axis_oarg_104_tstrb,
    output [M_AXIS_OARG_104_DMWIDTH-1:0] m_axis_oarg_104_tdata,
    input m_axis_oarg_104_tready,
    input ap_axis_oarg_104_tlast,
    input ap_axis_oarg_104_tvalid,
    input [M_AXIS_OARG_104_WIDTH/8-1:0] ap_axis_oarg_104_tkeep,
    input [M_AXIS_OARG_104_WIDTH/8-1:0] ap_axis_oarg_104_tstrb,
    input [M_AXIS_OARG_104_WIDTH-1:0] ap_axis_oarg_104_tdata,
    output ap_axis_oarg_104_tready,
    //output AXIS to AXI-Stream interface 105
    input m_axis_oarg_105_aclk,
    input m_axis_oarg_105_aresetn,
    output m_axis_oarg_105_tlast,
    output m_axis_oarg_105_tvalid,
    output [M_AXIS_OARG_105_DMWIDTH/8-1:0] m_axis_oarg_105_tkeep,
    output [M_AXIS_OARG_105_DMWIDTH/8-1:0] m_axis_oarg_105_tstrb,
    output [M_AXIS_OARG_105_DMWIDTH-1:0] m_axis_oarg_105_tdata,
    input m_axis_oarg_105_tready,
    input ap_axis_oarg_105_tlast,
    input ap_axis_oarg_105_tvalid,
    input [M_AXIS_OARG_105_WIDTH/8-1:0] ap_axis_oarg_105_tkeep,
    input [M_AXIS_OARG_105_WIDTH/8-1:0] ap_axis_oarg_105_tstrb,
    input [M_AXIS_OARG_105_WIDTH-1:0] ap_axis_oarg_105_tdata,
    output ap_axis_oarg_105_tready,
    //output AXIS to AXI-Stream interface 106
    input m_axis_oarg_106_aclk,
    input m_axis_oarg_106_aresetn,
    output m_axis_oarg_106_tlast,
    output m_axis_oarg_106_tvalid,
    output [M_AXIS_OARG_106_DMWIDTH/8-1:0] m_axis_oarg_106_tkeep,
    output [M_AXIS_OARG_106_DMWIDTH/8-1:0] m_axis_oarg_106_tstrb,
    output [M_AXIS_OARG_106_DMWIDTH-1:0] m_axis_oarg_106_tdata,
    input m_axis_oarg_106_tready,
    input ap_axis_oarg_106_tlast,
    input ap_axis_oarg_106_tvalid,
    input [M_AXIS_OARG_106_WIDTH/8-1:0] ap_axis_oarg_106_tkeep,
    input [M_AXIS_OARG_106_WIDTH/8-1:0] ap_axis_oarg_106_tstrb,
    input [M_AXIS_OARG_106_WIDTH-1:0] ap_axis_oarg_106_tdata,
    output ap_axis_oarg_106_tready,
    //output AXIS to AXI-Stream interface 107
    input m_axis_oarg_107_aclk,
    input m_axis_oarg_107_aresetn,
    output m_axis_oarg_107_tlast,
    output m_axis_oarg_107_tvalid,
    output [M_AXIS_OARG_107_DMWIDTH/8-1:0] m_axis_oarg_107_tkeep,
    output [M_AXIS_OARG_107_DMWIDTH/8-1:0] m_axis_oarg_107_tstrb,
    output [M_AXIS_OARG_107_DMWIDTH-1:0] m_axis_oarg_107_tdata,
    input m_axis_oarg_107_tready,
    input ap_axis_oarg_107_tlast,
    input ap_axis_oarg_107_tvalid,
    input [M_AXIS_OARG_107_WIDTH/8-1:0] ap_axis_oarg_107_tkeep,
    input [M_AXIS_OARG_107_WIDTH/8-1:0] ap_axis_oarg_107_tstrb,
    input [M_AXIS_OARG_107_WIDTH-1:0] ap_axis_oarg_107_tdata,
    output ap_axis_oarg_107_tready,
    //output AXIS to AXI-Stream interface 108
    input m_axis_oarg_108_aclk,
    input m_axis_oarg_108_aresetn,
    output m_axis_oarg_108_tlast,
    output m_axis_oarg_108_tvalid,
    output [M_AXIS_OARG_108_DMWIDTH/8-1:0] m_axis_oarg_108_tkeep,
    output [M_AXIS_OARG_108_DMWIDTH/8-1:0] m_axis_oarg_108_tstrb,
    output [M_AXIS_OARG_108_DMWIDTH-1:0] m_axis_oarg_108_tdata,
    input m_axis_oarg_108_tready,
    input ap_axis_oarg_108_tlast,
    input ap_axis_oarg_108_tvalid,
    input [M_AXIS_OARG_108_WIDTH/8-1:0] ap_axis_oarg_108_tkeep,
    input [M_AXIS_OARG_108_WIDTH/8-1:0] ap_axis_oarg_108_tstrb,
    input [M_AXIS_OARG_108_WIDTH-1:0] ap_axis_oarg_108_tdata,
    output ap_axis_oarg_108_tready,
    //output AXIS to AXI-Stream interface 109
    input m_axis_oarg_109_aclk,
    input m_axis_oarg_109_aresetn,
    output m_axis_oarg_109_tlast,
    output m_axis_oarg_109_tvalid,
    output [M_AXIS_OARG_109_DMWIDTH/8-1:0] m_axis_oarg_109_tkeep,
    output [M_AXIS_OARG_109_DMWIDTH/8-1:0] m_axis_oarg_109_tstrb,
    output [M_AXIS_OARG_109_DMWIDTH-1:0] m_axis_oarg_109_tdata,
    input m_axis_oarg_109_tready,
    input ap_axis_oarg_109_tlast,
    input ap_axis_oarg_109_tvalid,
    input [M_AXIS_OARG_109_WIDTH/8-1:0] ap_axis_oarg_109_tkeep,
    input [M_AXIS_OARG_109_WIDTH/8-1:0] ap_axis_oarg_109_tstrb,
    input [M_AXIS_OARG_109_WIDTH-1:0] ap_axis_oarg_109_tdata,
    output ap_axis_oarg_109_tready,
    //output AXIS to AXI-Stream interface 110
    input m_axis_oarg_110_aclk,
    input m_axis_oarg_110_aresetn,
    output m_axis_oarg_110_tlast,
    output m_axis_oarg_110_tvalid,
    output [M_AXIS_OARG_110_DMWIDTH/8-1:0] m_axis_oarg_110_tkeep,
    output [M_AXIS_OARG_110_DMWIDTH/8-1:0] m_axis_oarg_110_tstrb,
    output [M_AXIS_OARG_110_DMWIDTH-1:0] m_axis_oarg_110_tdata,
    input m_axis_oarg_110_tready,
    input ap_axis_oarg_110_tlast,
    input ap_axis_oarg_110_tvalid,
    input [M_AXIS_OARG_110_WIDTH/8-1:0] ap_axis_oarg_110_tkeep,
    input [M_AXIS_OARG_110_WIDTH/8-1:0] ap_axis_oarg_110_tstrb,
    input [M_AXIS_OARG_110_WIDTH-1:0] ap_axis_oarg_110_tdata,
    output ap_axis_oarg_110_tready,
    //output AXIS to AXI-Stream interface 111
    input m_axis_oarg_111_aclk,
    input m_axis_oarg_111_aresetn,
    output m_axis_oarg_111_tlast,
    output m_axis_oarg_111_tvalid,
    output [M_AXIS_OARG_111_DMWIDTH/8-1:0] m_axis_oarg_111_tkeep,
    output [M_AXIS_OARG_111_DMWIDTH/8-1:0] m_axis_oarg_111_tstrb,
    output [M_AXIS_OARG_111_DMWIDTH-1:0] m_axis_oarg_111_tdata,
    input m_axis_oarg_111_tready,
    input ap_axis_oarg_111_tlast,
    input ap_axis_oarg_111_tvalid,
    input [M_AXIS_OARG_111_WIDTH/8-1:0] ap_axis_oarg_111_tkeep,
    input [M_AXIS_OARG_111_WIDTH/8-1:0] ap_axis_oarg_111_tstrb,
    input [M_AXIS_OARG_111_WIDTH-1:0] ap_axis_oarg_111_tdata,
    output ap_axis_oarg_111_tready,
    //output AXIS to AXI-Stream interface 112
    input m_axis_oarg_112_aclk,
    input m_axis_oarg_112_aresetn,
    output m_axis_oarg_112_tlast,
    output m_axis_oarg_112_tvalid,
    output [M_AXIS_OARG_112_DMWIDTH/8-1:0] m_axis_oarg_112_tkeep,
    output [M_AXIS_OARG_112_DMWIDTH/8-1:0] m_axis_oarg_112_tstrb,
    output [M_AXIS_OARG_112_DMWIDTH-1:0] m_axis_oarg_112_tdata,
    input m_axis_oarg_112_tready,
    input ap_axis_oarg_112_tlast,
    input ap_axis_oarg_112_tvalid,
    input [M_AXIS_OARG_112_WIDTH/8-1:0] ap_axis_oarg_112_tkeep,
    input [M_AXIS_OARG_112_WIDTH/8-1:0] ap_axis_oarg_112_tstrb,
    input [M_AXIS_OARG_112_WIDTH-1:0] ap_axis_oarg_112_tdata,
    output ap_axis_oarg_112_tready,
    //output AXIS to AXI-Stream interface 113
    input m_axis_oarg_113_aclk,
    input m_axis_oarg_113_aresetn,
    output m_axis_oarg_113_tlast,
    output m_axis_oarg_113_tvalid,
    output [M_AXIS_OARG_113_DMWIDTH/8-1:0] m_axis_oarg_113_tkeep,
    output [M_AXIS_OARG_113_DMWIDTH/8-1:0] m_axis_oarg_113_tstrb,
    output [M_AXIS_OARG_113_DMWIDTH-1:0] m_axis_oarg_113_tdata,
    input m_axis_oarg_113_tready,
    input ap_axis_oarg_113_tlast,
    input ap_axis_oarg_113_tvalid,
    input [M_AXIS_OARG_113_WIDTH/8-1:0] ap_axis_oarg_113_tkeep,
    input [M_AXIS_OARG_113_WIDTH/8-1:0] ap_axis_oarg_113_tstrb,
    input [M_AXIS_OARG_113_WIDTH-1:0] ap_axis_oarg_113_tdata,
    output ap_axis_oarg_113_tready,
    //output AXIS to AXI-Stream interface 114
    input m_axis_oarg_114_aclk,
    input m_axis_oarg_114_aresetn,
    output m_axis_oarg_114_tlast,
    output m_axis_oarg_114_tvalid,
    output [M_AXIS_OARG_114_DMWIDTH/8-1:0] m_axis_oarg_114_tkeep,
    output [M_AXIS_OARG_114_DMWIDTH/8-1:0] m_axis_oarg_114_tstrb,
    output [M_AXIS_OARG_114_DMWIDTH-1:0] m_axis_oarg_114_tdata,
    input m_axis_oarg_114_tready,
    input ap_axis_oarg_114_tlast,
    input ap_axis_oarg_114_tvalid,
    input [M_AXIS_OARG_114_WIDTH/8-1:0] ap_axis_oarg_114_tkeep,
    input [M_AXIS_OARG_114_WIDTH/8-1:0] ap_axis_oarg_114_tstrb,
    input [M_AXIS_OARG_114_WIDTH-1:0] ap_axis_oarg_114_tdata,
    output ap_axis_oarg_114_tready,
    //output AXIS to AXI-Stream interface 115
    input m_axis_oarg_115_aclk,
    input m_axis_oarg_115_aresetn,
    output m_axis_oarg_115_tlast,
    output m_axis_oarg_115_tvalid,
    output [M_AXIS_OARG_115_DMWIDTH/8-1:0] m_axis_oarg_115_tkeep,
    output [M_AXIS_OARG_115_DMWIDTH/8-1:0] m_axis_oarg_115_tstrb,
    output [M_AXIS_OARG_115_DMWIDTH-1:0] m_axis_oarg_115_tdata,
    input m_axis_oarg_115_tready,
    input ap_axis_oarg_115_tlast,
    input ap_axis_oarg_115_tvalid,
    input [M_AXIS_OARG_115_WIDTH/8-1:0] ap_axis_oarg_115_tkeep,
    input [M_AXIS_OARG_115_WIDTH/8-1:0] ap_axis_oarg_115_tstrb,
    input [M_AXIS_OARG_115_WIDTH-1:0] ap_axis_oarg_115_tdata,
    output ap_axis_oarg_115_tready,
    //output AXIS to AXI-Stream interface 116
    input m_axis_oarg_116_aclk,
    input m_axis_oarg_116_aresetn,
    output m_axis_oarg_116_tlast,
    output m_axis_oarg_116_tvalid,
    output [M_AXIS_OARG_116_DMWIDTH/8-1:0] m_axis_oarg_116_tkeep,
    output [M_AXIS_OARG_116_DMWIDTH/8-1:0] m_axis_oarg_116_tstrb,
    output [M_AXIS_OARG_116_DMWIDTH-1:0] m_axis_oarg_116_tdata,
    input m_axis_oarg_116_tready,
    input ap_axis_oarg_116_tlast,
    input ap_axis_oarg_116_tvalid,
    input [M_AXIS_OARG_116_WIDTH/8-1:0] ap_axis_oarg_116_tkeep,
    input [M_AXIS_OARG_116_WIDTH/8-1:0] ap_axis_oarg_116_tstrb,
    input [M_AXIS_OARG_116_WIDTH-1:0] ap_axis_oarg_116_tdata,
    output ap_axis_oarg_116_tready,
    //output AXIS to AXI-Stream interface 117
    input m_axis_oarg_117_aclk,
    input m_axis_oarg_117_aresetn,
    output m_axis_oarg_117_tlast,
    output m_axis_oarg_117_tvalid,
    output [M_AXIS_OARG_117_DMWIDTH/8-1:0] m_axis_oarg_117_tkeep,
    output [M_AXIS_OARG_117_DMWIDTH/8-1:0] m_axis_oarg_117_tstrb,
    output [M_AXIS_OARG_117_DMWIDTH-1:0] m_axis_oarg_117_tdata,
    input m_axis_oarg_117_tready,
    input ap_axis_oarg_117_tlast,
    input ap_axis_oarg_117_tvalid,
    input [M_AXIS_OARG_117_WIDTH/8-1:0] ap_axis_oarg_117_tkeep,
    input [M_AXIS_OARG_117_WIDTH/8-1:0] ap_axis_oarg_117_tstrb,
    input [M_AXIS_OARG_117_WIDTH-1:0] ap_axis_oarg_117_tdata,
    output ap_axis_oarg_117_tready,
    //output AXIS to AXI-Stream interface 118
    input m_axis_oarg_118_aclk,
    input m_axis_oarg_118_aresetn,
    output m_axis_oarg_118_tlast,
    output m_axis_oarg_118_tvalid,
    output [M_AXIS_OARG_118_DMWIDTH/8-1:0] m_axis_oarg_118_tkeep,
    output [M_AXIS_OARG_118_DMWIDTH/8-1:0] m_axis_oarg_118_tstrb,
    output [M_AXIS_OARG_118_DMWIDTH-1:0] m_axis_oarg_118_tdata,
    input m_axis_oarg_118_tready,
    input ap_axis_oarg_118_tlast,
    input ap_axis_oarg_118_tvalid,
    input [M_AXIS_OARG_118_WIDTH/8-1:0] ap_axis_oarg_118_tkeep,
    input [M_AXIS_OARG_118_WIDTH/8-1:0] ap_axis_oarg_118_tstrb,
    input [M_AXIS_OARG_118_WIDTH-1:0] ap_axis_oarg_118_tdata,
    output ap_axis_oarg_118_tready,
    //output AXIS to AXI-Stream interface 119
    input m_axis_oarg_119_aclk,
    input m_axis_oarg_119_aresetn,
    output m_axis_oarg_119_tlast,
    output m_axis_oarg_119_tvalid,
    output [M_AXIS_OARG_119_DMWIDTH/8-1:0] m_axis_oarg_119_tkeep,
    output [M_AXIS_OARG_119_DMWIDTH/8-1:0] m_axis_oarg_119_tstrb,
    output [M_AXIS_OARG_119_DMWIDTH-1:0] m_axis_oarg_119_tdata,
    input m_axis_oarg_119_tready,
    input ap_axis_oarg_119_tlast,
    input ap_axis_oarg_119_tvalid,
    input [M_AXIS_OARG_119_WIDTH/8-1:0] ap_axis_oarg_119_tkeep,
    input [M_AXIS_OARG_119_WIDTH/8-1:0] ap_axis_oarg_119_tstrb,
    input [M_AXIS_OARG_119_WIDTH-1:0] ap_axis_oarg_119_tdata,
    output ap_axis_oarg_119_tready,
    //output AXIS to AXI-Stream interface 120
    input m_axis_oarg_120_aclk,
    input m_axis_oarg_120_aresetn,
    output m_axis_oarg_120_tlast,
    output m_axis_oarg_120_tvalid,
    output [M_AXIS_OARG_120_DMWIDTH/8-1:0] m_axis_oarg_120_tkeep,
    output [M_AXIS_OARG_120_DMWIDTH/8-1:0] m_axis_oarg_120_tstrb,
    output [M_AXIS_OARG_120_DMWIDTH-1:0] m_axis_oarg_120_tdata,
    input m_axis_oarg_120_tready,
    input ap_axis_oarg_120_tlast,
    input ap_axis_oarg_120_tvalid,
    input [M_AXIS_OARG_120_WIDTH/8-1:0] ap_axis_oarg_120_tkeep,
    input [M_AXIS_OARG_120_WIDTH/8-1:0] ap_axis_oarg_120_tstrb,
    input [M_AXIS_OARG_120_WIDTH-1:0] ap_axis_oarg_120_tdata,
    output ap_axis_oarg_120_tready,
    //output AXIS to AXI-Stream interface 121
    input m_axis_oarg_121_aclk,
    input m_axis_oarg_121_aresetn,
    output m_axis_oarg_121_tlast,
    output m_axis_oarg_121_tvalid,
    output [M_AXIS_OARG_121_DMWIDTH/8-1:0] m_axis_oarg_121_tkeep,
    output [M_AXIS_OARG_121_DMWIDTH/8-1:0] m_axis_oarg_121_tstrb,
    output [M_AXIS_OARG_121_DMWIDTH-1:0] m_axis_oarg_121_tdata,
    input m_axis_oarg_121_tready,
    input ap_axis_oarg_121_tlast,
    input ap_axis_oarg_121_tvalid,
    input [M_AXIS_OARG_121_WIDTH/8-1:0] ap_axis_oarg_121_tkeep,
    input [M_AXIS_OARG_121_WIDTH/8-1:0] ap_axis_oarg_121_tstrb,
    input [M_AXIS_OARG_121_WIDTH-1:0] ap_axis_oarg_121_tdata,
    output ap_axis_oarg_121_tready,
    //output AXIS to AXI-Stream interface 122
    input m_axis_oarg_122_aclk,
    input m_axis_oarg_122_aresetn,
    output m_axis_oarg_122_tlast,
    output m_axis_oarg_122_tvalid,
    output [M_AXIS_OARG_122_DMWIDTH/8-1:0] m_axis_oarg_122_tkeep,
    output [M_AXIS_OARG_122_DMWIDTH/8-1:0] m_axis_oarg_122_tstrb,
    output [M_AXIS_OARG_122_DMWIDTH-1:0] m_axis_oarg_122_tdata,
    input m_axis_oarg_122_tready,
    input ap_axis_oarg_122_tlast,
    input ap_axis_oarg_122_tvalid,
    input [M_AXIS_OARG_122_WIDTH/8-1:0] ap_axis_oarg_122_tkeep,
    input [M_AXIS_OARG_122_WIDTH/8-1:0] ap_axis_oarg_122_tstrb,
    input [M_AXIS_OARG_122_WIDTH-1:0] ap_axis_oarg_122_tdata,
    output ap_axis_oarg_122_tready,
    //output AXIS to AXI-Stream interface 123
    input m_axis_oarg_123_aclk,
    input m_axis_oarg_123_aresetn,
    output m_axis_oarg_123_tlast,
    output m_axis_oarg_123_tvalid,
    output [M_AXIS_OARG_123_DMWIDTH/8-1:0] m_axis_oarg_123_tkeep,
    output [M_AXIS_OARG_123_DMWIDTH/8-1:0] m_axis_oarg_123_tstrb,
    output [M_AXIS_OARG_123_DMWIDTH-1:0] m_axis_oarg_123_tdata,
    input m_axis_oarg_123_tready,
    input ap_axis_oarg_123_tlast,
    input ap_axis_oarg_123_tvalid,
    input [M_AXIS_OARG_123_WIDTH/8-1:0] ap_axis_oarg_123_tkeep,
    input [M_AXIS_OARG_123_WIDTH/8-1:0] ap_axis_oarg_123_tstrb,
    input [M_AXIS_OARG_123_WIDTH-1:0] ap_axis_oarg_123_tdata,
    output ap_axis_oarg_123_tready,
    //output AXIS to AXI-Stream interface 124
    input m_axis_oarg_124_aclk,
    input m_axis_oarg_124_aresetn,
    output m_axis_oarg_124_tlast,
    output m_axis_oarg_124_tvalid,
    output [M_AXIS_OARG_124_DMWIDTH/8-1:0] m_axis_oarg_124_tkeep,
    output [M_AXIS_OARG_124_DMWIDTH/8-1:0] m_axis_oarg_124_tstrb,
    output [M_AXIS_OARG_124_DMWIDTH-1:0] m_axis_oarg_124_tdata,
    input m_axis_oarg_124_tready,
    input ap_axis_oarg_124_tlast,
    input ap_axis_oarg_124_tvalid,
    input [M_AXIS_OARG_124_WIDTH/8-1:0] ap_axis_oarg_124_tkeep,
    input [M_AXIS_OARG_124_WIDTH/8-1:0] ap_axis_oarg_124_tstrb,
    input [M_AXIS_OARG_124_WIDTH-1:0] ap_axis_oarg_124_tdata,
    output ap_axis_oarg_124_tready,
    //output AXIS to AXI-Stream interface 125
    input m_axis_oarg_125_aclk,
    input m_axis_oarg_125_aresetn,
    output m_axis_oarg_125_tlast,
    output m_axis_oarg_125_tvalid,
    output [M_AXIS_OARG_125_DMWIDTH/8-1:0] m_axis_oarg_125_tkeep,
    output [M_AXIS_OARG_125_DMWIDTH/8-1:0] m_axis_oarg_125_tstrb,
    output [M_AXIS_OARG_125_DMWIDTH-1:0] m_axis_oarg_125_tdata,
    input m_axis_oarg_125_tready,
    input ap_axis_oarg_125_tlast,
    input ap_axis_oarg_125_tvalid,
    input [M_AXIS_OARG_125_WIDTH/8-1:0] ap_axis_oarg_125_tkeep,
    input [M_AXIS_OARG_125_WIDTH/8-1:0] ap_axis_oarg_125_tstrb,
    input [M_AXIS_OARG_125_WIDTH-1:0] ap_axis_oarg_125_tdata,
    output ap_axis_oarg_125_tready,
    //output AXIS to AXI-Stream interface 126
    input m_axis_oarg_126_aclk,
    input m_axis_oarg_126_aresetn,
    output m_axis_oarg_126_tlast,
    output m_axis_oarg_126_tvalid,
    output [M_AXIS_OARG_126_DMWIDTH/8-1:0] m_axis_oarg_126_tkeep,
    output [M_AXIS_OARG_126_DMWIDTH/8-1:0] m_axis_oarg_126_tstrb,
    output [M_AXIS_OARG_126_DMWIDTH-1:0] m_axis_oarg_126_tdata,
    input m_axis_oarg_126_tready,
    input ap_axis_oarg_126_tlast,
    input ap_axis_oarg_126_tvalid,
    input [M_AXIS_OARG_126_WIDTH/8-1:0] ap_axis_oarg_126_tkeep,
    input [M_AXIS_OARG_126_WIDTH/8-1:0] ap_axis_oarg_126_tstrb,
    input [M_AXIS_OARG_126_WIDTH-1:0] ap_axis_oarg_126_tdata,
    output ap_axis_oarg_126_tready,
    //output AXIS to AXI-Stream interface 127
    input m_axis_oarg_127_aclk,
    input m_axis_oarg_127_aresetn,
    output m_axis_oarg_127_tlast,
    output m_axis_oarg_127_tvalid,
    output [M_AXIS_OARG_127_DMWIDTH/8-1:0] m_axis_oarg_127_tkeep,
    output [M_AXIS_OARG_127_DMWIDTH/8-1:0] m_axis_oarg_127_tstrb,
    output [M_AXIS_OARG_127_DMWIDTH-1:0] m_axis_oarg_127_tdata,
    input m_axis_oarg_127_tready,
    input ap_axis_oarg_127_tlast,
    input ap_axis_oarg_127_tvalid,
    input [M_AXIS_OARG_127_WIDTH/8-1:0] ap_axis_oarg_127_tkeep,
    input [M_AXIS_OARG_127_WIDTH/8-1:0] ap_axis_oarg_127_tstrb,
    input [M_AXIS_OARG_127_WIDTH-1:0] ap_axis_oarg_127_tdata,
    output ap_axis_oarg_127_tready
    );


    localparam C_MAX_OUTPUT_AXISs = 128;
    localparam C_MAX_BIT_WIDTH = 1024;
    localparam [(C_MAX_OUTPUT_AXISs*32)-1:0] C_OUTAXIS_BIT_ARRAY = {M_AXIS_OARG_127_WIDTH,M_AXIS_OARG_126_WIDTH,M_AXIS_OARG_125_WIDTH,M_AXIS_OARG_124_WIDTH,M_AXIS_OARG_123_WIDTH,M_AXIS_OARG_122_WIDTH,M_AXIS_OARG_121_WIDTH,M_AXIS_OARG_120_WIDTH,M_AXIS_OARG_119_WIDTH,M_AXIS_OARG_118_WIDTH,M_AXIS_OARG_117_WIDTH,M_AXIS_OARG_116_WIDTH,M_AXIS_OARG_115_WIDTH,M_AXIS_OARG_114_WIDTH,M_AXIS_OARG_113_WIDTH,M_AXIS_OARG_112_WIDTH,M_AXIS_OARG_111_WIDTH,M_AXIS_OARG_110_WIDTH,M_AXIS_OARG_109_WIDTH,M_AXIS_OARG_108_WIDTH,M_AXIS_OARG_107_WIDTH,M_AXIS_OARG_106_WIDTH,M_AXIS_OARG_105_WIDTH,M_AXIS_OARG_104_WIDTH,M_AXIS_OARG_103_WIDTH,M_AXIS_OARG_102_WIDTH,M_AXIS_OARG_101_WIDTH,M_AXIS_OARG_100_WIDTH,M_AXIS_OARG_99_WIDTH,M_AXIS_OARG_98_WIDTH,M_AXIS_OARG_97_WIDTH,M_AXIS_OARG_96_WIDTH,M_AXIS_OARG_95_WIDTH,M_AXIS_OARG_94_WIDTH,M_AXIS_OARG_93_WIDTH,M_AXIS_OARG_92_WIDTH,M_AXIS_OARG_91_WIDTH,M_AXIS_OARG_90_WIDTH,M_AXIS_OARG_89_WIDTH,M_AXIS_OARG_88_WIDTH,M_AXIS_OARG_87_WIDTH,M_AXIS_OARG_86_WIDTH,M_AXIS_OARG_85_WIDTH,M_AXIS_OARG_84_WIDTH,M_AXIS_OARG_83_WIDTH,M_AXIS_OARG_82_WIDTH,M_AXIS_OARG_81_WIDTH,M_AXIS_OARG_80_WIDTH,M_AXIS_OARG_79_WIDTH,M_AXIS_OARG_78_WIDTH,M_AXIS_OARG_77_WIDTH,M_AXIS_OARG_76_WIDTH,M_AXIS_OARG_75_WIDTH,M_AXIS_OARG_74_WIDTH,M_AXIS_OARG_73_WIDTH,M_AXIS_OARG_72_WIDTH,M_AXIS_OARG_71_WIDTH,M_AXIS_OARG_70_WIDTH,M_AXIS_OARG_69_WIDTH,M_AXIS_OARG_68_WIDTH,M_AXIS_OARG_67_WIDTH,M_AXIS_OARG_66_WIDTH,M_AXIS_OARG_65_WIDTH,M_AXIS_OARG_64_WIDTH,M_AXIS_OARG_63_WIDTH,M_AXIS_OARG_62_WIDTH,M_AXIS_OARG_61_WIDTH,M_AXIS_OARG_60_WIDTH,M_AXIS_OARG_59_WIDTH,M_AXIS_OARG_58_WIDTH,M_AXIS_OARG_57_WIDTH,M_AXIS_OARG_56_WIDTH,M_AXIS_OARG_55_WIDTH,M_AXIS_OARG_54_WIDTH,M_AXIS_OARG_53_WIDTH,M_AXIS_OARG_52_WIDTH,M_AXIS_OARG_51_WIDTH,M_AXIS_OARG_50_WIDTH,M_AXIS_OARG_49_WIDTH,M_AXIS_OARG_48_WIDTH,M_AXIS_OARG_47_WIDTH,M_AXIS_OARG_46_WIDTH,M_AXIS_OARG_45_WIDTH,M_AXIS_OARG_44_WIDTH,M_AXIS_OARG_43_WIDTH,M_AXIS_OARG_42_WIDTH,M_AXIS_OARG_41_WIDTH,M_AXIS_OARG_40_WIDTH,M_AXIS_OARG_39_WIDTH,M_AXIS_OARG_38_WIDTH,M_AXIS_OARG_37_WIDTH,M_AXIS_OARG_36_WIDTH,M_AXIS_OARG_35_WIDTH,M_AXIS_OARG_34_WIDTH,M_AXIS_OARG_33_WIDTH,M_AXIS_OARG_32_WIDTH,M_AXIS_OARG_31_WIDTH,M_AXIS_OARG_30_WIDTH,M_AXIS_OARG_29_WIDTH,M_AXIS_OARG_28_WIDTH,M_AXIS_OARG_27_WIDTH,M_AXIS_OARG_26_WIDTH,M_AXIS_OARG_25_WIDTH,M_AXIS_OARG_24_WIDTH,M_AXIS_OARG_23_WIDTH,M_AXIS_OARG_22_WIDTH,M_AXIS_OARG_21_WIDTH,M_AXIS_OARG_20_WIDTH,M_AXIS_OARG_19_WIDTH,M_AXIS_OARG_18_WIDTH,M_AXIS_OARG_17_WIDTH,M_AXIS_OARG_16_WIDTH,M_AXIS_OARG_15_WIDTH,M_AXIS_OARG_14_WIDTH,M_AXIS_OARG_13_WIDTH,M_AXIS_OARG_12_WIDTH,M_AXIS_OARG_11_WIDTH,M_AXIS_OARG_10_WIDTH,M_AXIS_OARG_9_WIDTH,M_AXIS_OARG_8_WIDTH,M_AXIS_OARG_7_WIDTH,M_AXIS_OARG_6_WIDTH,M_AXIS_OARG_5_WIDTH,M_AXIS_OARG_4_WIDTH,M_AXIS_OARG_3_WIDTH,M_AXIS_OARG_2_WIDTH,M_AXIS_OARG_1_WIDTH,M_AXIS_OARG_0_WIDTH};
    localparam [(C_MAX_OUTPUT_AXISs*32)-1:0] C_DEPTH_BIT_ARRAY = {M_AXIS_OARG_127_DEPTH,M_AXIS_OARG_126_DEPTH,M_AXIS_OARG_125_DEPTH,M_AXIS_OARG_124_DEPTH,M_AXIS_OARG_123_DEPTH,M_AXIS_OARG_122_DEPTH,M_AXIS_OARG_121_DEPTH,M_AXIS_OARG_120_DEPTH,M_AXIS_OARG_119_DEPTH,M_AXIS_OARG_118_DEPTH,M_AXIS_OARG_117_DEPTH,M_AXIS_OARG_116_DEPTH,M_AXIS_OARG_115_DEPTH,M_AXIS_OARG_114_DEPTH,M_AXIS_OARG_113_DEPTH,M_AXIS_OARG_112_DEPTH,M_AXIS_OARG_111_DEPTH,M_AXIS_OARG_110_DEPTH,M_AXIS_OARG_109_DEPTH,M_AXIS_OARG_108_DEPTH,M_AXIS_OARG_107_DEPTH,M_AXIS_OARG_106_DEPTH,M_AXIS_OARG_105_DEPTH,M_AXIS_OARG_104_DEPTH,M_AXIS_OARG_103_DEPTH,M_AXIS_OARG_102_DEPTH,M_AXIS_OARG_101_DEPTH,M_AXIS_OARG_100_DEPTH,M_AXIS_OARG_99_DEPTH,M_AXIS_OARG_98_DEPTH,M_AXIS_OARG_97_DEPTH,M_AXIS_OARG_96_DEPTH,M_AXIS_OARG_95_DEPTH,M_AXIS_OARG_94_DEPTH,M_AXIS_OARG_93_DEPTH,M_AXIS_OARG_92_DEPTH,M_AXIS_OARG_91_DEPTH,M_AXIS_OARG_90_DEPTH,M_AXIS_OARG_89_DEPTH,M_AXIS_OARG_88_DEPTH,M_AXIS_OARG_87_DEPTH,M_AXIS_OARG_86_DEPTH,M_AXIS_OARG_85_DEPTH,M_AXIS_OARG_84_DEPTH,M_AXIS_OARG_83_DEPTH,M_AXIS_OARG_82_DEPTH,M_AXIS_OARG_81_DEPTH,M_AXIS_OARG_80_DEPTH,M_AXIS_OARG_79_DEPTH,M_AXIS_OARG_78_DEPTH,M_AXIS_OARG_77_DEPTH,M_AXIS_OARG_76_DEPTH,M_AXIS_OARG_75_DEPTH,M_AXIS_OARG_74_DEPTH,M_AXIS_OARG_73_DEPTH,M_AXIS_OARG_72_DEPTH,M_AXIS_OARG_71_DEPTH,M_AXIS_OARG_70_DEPTH,M_AXIS_OARG_69_DEPTH,M_AXIS_OARG_68_DEPTH,M_AXIS_OARG_67_DEPTH,M_AXIS_OARG_66_DEPTH,M_AXIS_OARG_65_DEPTH,M_AXIS_OARG_64_DEPTH,M_AXIS_OARG_63_DEPTH,M_AXIS_OARG_62_DEPTH,M_AXIS_OARG_61_DEPTH,M_AXIS_OARG_60_DEPTH,M_AXIS_OARG_59_DEPTH,M_AXIS_OARG_58_DEPTH,M_AXIS_OARG_57_DEPTH,M_AXIS_OARG_56_DEPTH,M_AXIS_OARG_55_DEPTH,M_AXIS_OARG_54_DEPTH,M_AXIS_OARG_53_DEPTH,M_AXIS_OARG_52_DEPTH,M_AXIS_OARG_51_DEPTH,M_AXIS_OARG_50_DEPTH,M_AXIS_OARG_49_DEPTH,M_AXIS_OARG_48_DEPTH,M_AXIS_OARG_47_DEPTH,M_AXIS_OARG_46_DEPTH,M_AXIS_OARG_45_DEPTH,M_AXIS_OARG_44_DEPTH,M_AXIS_OARG_43_DEPTH,M_AXIS_OARG_42_DEPTH,M_AXIS_OARG_41_DEPTH,M_AXIS_OARG_40_DEPTH,M_AXIS_OARG_39_DEPTH,M_AXIS_OARG_38_DEPTH,M_AXIS_OARG_37_DEPTH,M_AXIS_OARG_36_DEPTH,M_AXIS_OARG_35_DEPTH,M_AXIS_OARG_34_DEPTH,M_AXIS_OARG_33_DEPTH,M_AXIS_OARG_32_DEPTH,M_AXIS_OARG_31_DEPTH,M_AXIS_OARG_30_DEPTH,M_AXIS_OARG_29_DEPTH,M_AXIS_OARG_28_DEPTH,M_AXIS_OARG_27_DEPTH,M_AXIS_OARG_26_DEPTH,M_AXIS_OARG_25_DEPTH,M_AXIS_OARG_24_DEPTH,M_AXIS_OARG_23_DEPTH,M_AXIS_OARG_22_DEPTH,M_AXIS_OARG_21_DEPTH,M_AXIS_OARG_20_DEPTH,M_AXIS_OARG_19_DEPTH,M_AXIS_OARG_18_DEPTH,M_AXIS_OARG_17_DEPTH,M_AXIS_OARG_16_DEPTH,M_AXIS_OARG_15_DEPTH,M_AXIS_OARG_14_DEPTH,M_AXIS_OARG_13_DEPTH,M_AXIS_OARG_12_DEPTH,M_AXIS_OARG_11_DEPTH,M_AXIS_OARG_10_DEPTH,M_AXIS_OARG_9_DEPTH,M_AXIS_OARG_8_DEPTH,M_AXIS_OARG_7_DEPTH,M_AXIS_OARG_6_DEPTH,M_AXIS_OARG_5_DEPTH,M_AXIS_OARG_4_DEPTH,M_AXIS_OARG_3_DEPTH,M_AXIS_OARG_2_DEPTH,M_AXIS_OARG_1_DEPTH,M_AXIS_OARG_0_DEPTH};
    localparam [(C_MAX_OUTPUT_AXISs*32)-1:0] C_DMWIDTH_BIT_ARRAY = {M_AXIS_OARG_127_DMWIDTH,M_AXIS_OARG_126_DMWIDTH,M_AXIS_OARG_125_DMWIDTH,M_AXIS_OARG_124_DMWIDTH,M_AXIS_OARG_123_DMWIDTH,M_AXIS_OARG_122_DMWIDTH,M_AXIS_OARG_121_DMWIDTH,M_AXIS_OARG_120_DMWIDTH,M_AXIS_OARG_119_DMWIDTH,M_AXIS_OARG_118_DMWIDTH,M_AXIS_OARG_117_DMWIDTH,M_AXIS_OARG_116_DMWIDTH,M_AXIS_OARG_115_DMWIDTH,M_AXIS_OARG_114_DMWIDTH,M_AXIS_OARG_113_DMWIDTH,M_AXIS_OARG_112_DMWIDTH,M_AXIS_OARG_111_DMWIDTH,M_AXIS_OARG_110_DMWIDTH,M_AXIS_OARG_109_DMWIDTH,M_AXIS_OARG_108_DMWIDTH,M_AXIS_OARG_107_DMWIDTH,M_AXIS_OARG_106_DMWIDTH,M_AXIS_OARG_105_DMWIDTH,M_AXIS_OARG_104_DMWIDTH,M_AXIS_OARG_103_DMWIDTH,M_AXIS_OARG_102_DMWIDTH,M_AXIS_OARG_101_DMWIDTH,M_AXIS_OARG_100_DMWIDTH,M_AXIS_OARG_99_DMWIDTH,M_AXIS_OARG_98_DMWIDTH,M_AXIS_OARG_97_DMWIDTH,M_AXIS_OARG_96_DMWIDTH,M_AXIS_OARG_95_DMWIDTH,M_AXIS_OARG_94_DMWIDTH,M_AXIS_OARG_93_DMWIDTH,M_AXIS_OARG_92_DMWIDTH,M_AXIS_OARG_91_DMWIDTH,M_AXIS_OARG_90_DMWIDTH,M_AXIS_OARG_89_DMWIDTH,M_AXIS_OARG_88_DMWIDTH,M_AXIS_OARG_87_DMWIDTH,M_AXIS_OARG_86_DMWIDTH,M_AXIS_OARG_85_DMWIDTH,M_AXIS_OARG_84_DMWIDTH,M_AXIS_OARG_83_DMWIDTH,M_AXIS_OARG_82_DMWIDTH,M_AXIS_OARG_81_DMWIDTH,M_AXIS_OARG_80_DMWIDTH,M_AXIS_OARG_79_DMWIDTH,M_AXIS_OARG_78_DMWIDTH,M_AXIS_OARG_77_DMWIDTH,M_AXIS_OARG_76_DMWIDTH,M_AXIS_OARG_75_DMWIDTH,M_AXIS_OARG_74_DMWIDTH,M_AXIS_OARG_73_DMWIDTH,M_AXIS_OARG_72_DMWIDTH,M_AXIS_OARG_71_DMWIDTH,M_AXIS_OARG_70_DMWIDTH,M_AXIS_OARG_69_DMWIDTH,M_AXIS_OARG_68_DMWIDTH,M_AXIS_OARG_67_DMWIDTH,M_AXIS_OARG_66_DMWIDTH,M_AXIS_OARG_65_DMWIDTH,M_AXIS_OARG_64_DMWIDTH,M_AXIS_OARG_63_DMWIDTH,M_AXIS_OARG_62_DMWIDTH,M_AXIS_OARG_61_DMWIDTH,M_AXIS_OARG_60_DMWIDTH,M_AXIS_OARG_59_DMWIDTH,M_AXIS_OARG_58_DMWIDTH,M_AXIS_OARG_57_DMWIDTH,M_AXIS_OARG_56_DMWIDTH,M_AXIS_OARG_55_DMWIDTH,M_AXIS_OARG_54_DMWIDTH,M_AXIS_OARG_53_DMWIDTH,M_AXIS_OARG_52_DMWIDTH,M_AXIS_OARG_51_DMWIDTH,M_AXIS_OARG_50_DMWIDTH,M_AXIS_OARG_49_DMWIDTH,M_AXIS_OARG_48_DMWIDTH,M_AXIS_OARG_47_DMWIDTH,M_AXIS_OARG_46_DMWIDTH,M_AXIS_OARG_45_DMWIDTH,M_AXIS_OARG_44_DMWIDTH,M_AXIS_OARG_43_DMWIDTH,M_AXIS_OARG_42_DMWIDTH,M_AXIS_OARG_41_DMWIDTH,M_AXIS_OARG_40_DMWIDTH,M_AXIS_OARG_39_DMWIDTH,M_AXIS_OARG_38_DMWIDTH,M_AXIS_OARG_37_DMWIDTH,M_AXIS_OARG_36_DMWIDTH,M_AXIS_OARG_35_DMWIDTH,M_AXIS_OARG_34_DMWIDTH,M_AXIS_OARG_33_DMWIDTH,M_AXIS_OARG_32_DMWIDTH,M_AXIS_OARG_31_DMWIDTH,M_AXIS_OARG_30_DMWIDTH,M_AXIS_OARG_29_DMWIDTH,M_AXIS_OARG_28_DMWIDTH,M_AXIS_OARG_27_DMWIDTH,M_AXIS_OARG_26_DMWIDTH,M_AXIS_OARG_25_DMWIDTH,M_AXIS_OARG_24_DMWIDTH,M_AXIS_OARG_23_DMWIDTH,M_AXIS_OARG_22_DMWIDTH,M_AXIS_OARG_21_DMWIDTH,M_AXIS_OARG_20_DMWIDTH,M_AXIS_OARG_19_DMWIDTH,M_AXIS_OARG_18_DMWIDTH,M_AXIS_OARG_17_DMWIDTH,M_AXIS_OARG_16_DMWIDTH,M_AXIS_OARG_15_DMWIDTH,M_AXIS_OARG_14_DMWIDTH,M_AXIS_OARG_13_DMWIDTH,M_AXIS_OARG_12_DMWIDTH,M_AXIS_OARG_11_DMWIDTH,M_AXIS_OARG_10_DMWIDTH,M_AXIS_OARG_9_DMWIDTH,M_AXIS_OARG_8_DMWIDTH,M_AXIS_OARG_7_DMWIDTH,M_AXIS_OARG_6_DMWIDTH,M_AXIS_OARG_5_DMWIDTH,M_AXIS_OARG_4_DMWIDTH,M_AXIS_OARG_3_DMWIDTH,M_AXIS_OARG_2_DMWIDTH,M_AXIS_OARG_1_DMWIDTH,M_AXIS_OARG_0_DMWIDTH};
    localparam [(C_MAX_OUTPUT_AXISs*32)-1:0] C_IS_ASYNC_BIT_ARRAY = {M_AXIS_OARG_127_IS_ASYNC,M_AXIS_OARG_126_IS_ASYNC,M_AXIS_OARG_125_IS_ASYNC,M_AXIS_OARG_124_IS_ASYNC,M_AXIS_OARG_123_IS_ASYNC,M_AXIS_OARG_122_IS_ASYNC,M_AXIS_OARG_121_IS_ASYNC,M_AXIS_OARG_120_IS_ASYNC,M_AXIS_OARG_119_IS_ASYNC,M_AXIS_OARG_118_IS_ASYNC,M_AXIS_OARG_117_IS_ASYNC,M_AXIS_OARG_116_IS_ASYNC,M_AXIS_OARG_115_IS_ASYNC,M_AXIS_OARG_114_IS_ASYNC,M_AXIS_OARG_113_IS_ASYNC,M_AXIS_OARG_112_IS_ASYNC,M_AXIS_OARG_111_IS_ASYNC,M_AXIS_OARG_110_IS_ASYNC,M_AXIS_OARG_109_IS_ASYNC,M_AXIS_OARG_108_IS_ASYNC,M_AXIS_OARG_107_IS_ASYNC,M_AXIS_OARG_106_IS_ASYNC,M_AXIS_OARG_105_IS_ASYNC,M_AXIS_OARG_104_IS_ASYNC,M_AXIS_OARG_103_IS_ASYNC,M_AXIS_OARG_102_IS_ASYNC,M_AXIS_OARG_101_IS_ASYNC,M_AXIS_OARG_100_IS_ASYNC,M_AXIS_OARG_99_IS_ASYNC,M_AXIS_OARG_98_IS_ASYNC,M_AXIS_OARG_97_IS_ASYNC,M_AXIS_OARG_96_IS_ASYNC,M_AXIS_OARG_95_IS_ASYNC,M_AXIS_OARG_94_IS_ASYNC,M_AXIS_OARG_93_IS_ASYNC,M_AXIS_OARG_92_IS_ASYNC,M_AXIS_OARG_91_IS_ASYNC,M_AXIS_OARG_90_IS_ASYNC,M_AXIS_OARG_89_IS_ASYNC,M_AXIS_OARG_88_IS_ASYNC,M_AXIS_OARG_87_IS_ASYNC,M_AXIS_OARG_86_IS_ASYNC,M_AXIS_OARG_85_IS_ASYNC,M_AXIS_OARG_84_IS_ASYNC,M_AXIS_OARG_83_IS_ASYNC,M_AXIS_OARG_82_IS_ASYNC,M_AXIS_OARG_81_IS_ASYNC,M_AXIS_OARG_80_IS_ASYNC,M_AXIS_OARG_79_IS_ASYNC,M_AXIS_OARG_78_IS_ASYNC,M_AXIS_OARG_77_IS_ASYNC,M_AXIS_OARG_76_IS_ASYNC,M_AXIS_OARG_75_IS_ASYNC,M_AXIS_OARG_74_IS_ASYNC,M_AXIS_OARG_73_IS_ASYNC,M_AXIS_OARG_72_IS_ASYNC,M_AXIS_OARG_71_IS_ASYNC,M_AXIS_OARG_70_IS_ASYNC,M_AXIS_OARG_69_IS_ASYNC,M_AXIS_OARG_68_IS_ASYNC,M_AXIS_OARG_67_IS_ASYNC,M_AXIS_OARG_66_IS_ASYNC,M_AXIS_OARG_65_IS_ASYNC,M_AXIS_OARG_64_IS_ASYNC,M_AXIS_OARG_63_IS_ASYNC,M_AXIS_OARG_62_IS_ASYNC,M_AXIS_OARG_61_IS_ASYNC,M_AXIS_OARG_60_IS_ASYNC,M_AXIS_OARG_59_IS_ASYNC,M_AXIS_OARG_58_IS_ASYNC,M_AXIS_OARG_57_IS_ASYNC,M_AXIS_OARG_56_IS_ASYNC,M_AXIS_OARG_55_IS_ASYNC,M_AXIS_OARG_54_IS_ASYNC,M_AXIS_OARG_53_IS_ASYNC,M_AXIS_OARG_52_IS_ASYNC,M_AXIS_OARG_51_IS_ASYNC,M_AXIS_OARG_50_IS_ASYNC,M_AXIS_OARG_49_IS_ASYNC,M_AXIS_OARG_48_IS_ASYNC,M_AXIS_OARG_47_IS_ASYNC,M_AXIS_OARG_46_IS_ASYNC,M_AXIS_OARG_45_IS_ASYNC,M_AXIS_OARG_44_IS_ASYNC,M_AXIS_OARG_43_IS_ASYNC,M_AXIS_OARG_42_IS_ASYNC,M_AXIS_OARG_41_IS_ASYNC,M_AXIS_OARG_40_IS_ASYNC,M_AXIS_OARG_39_IS_ASYNC,M_AXIS_OARG_38_IS_ASYNC,M_AXIS_OARG_37_IS_ASYNC,M_AXIS_OARG_36_IS_ASYNC,M_AXIS_OARG_35_IS_ASYNC,M_AXIS_OARG_34_IS_ASYNC,M_AXIS_OARG_33_IS_ASYNC,M_AXIS_OARG_32_IS_ASYNC,M_AXIS_OARG_31_IS_ASYNC,M_AXIS_OARG_30_IS_ASYNC,M_AXIS_OARG_29_IS_ASYNC,M_AXIS_OARG_28_IS_ASYNC,M_AXIS_OARG_27_IS_ASYNC,M_AXIS_OARG_26_IS_ASYNC,M_AXIS_OARG_25_IS_ASYNC,M_AXIS_OARG_24_IS_ASYNC,M_AXIS_OARG_23_IS_ASYNC,M_AXIS_OARG_22_IS_ASYNC,M_AXIS_OARG_21_IS_ASYNC,M_AXIS_OARG_20_IS_ASYNC,M_AXIS_OARG_19_IS_ASYNC,M_AXIS_OARG_18_IS_ASYNC,M_AXIS_OARG_17_IS_ASYNC,M_AXIS_OARG_16_IS_ASYNC,M_AXIS_OARG_15_IS_ASYNC,M_AXIS_OARG_14_IS_ASYNC,M_AXIS_OARG_13_IS_ASYNC,M_AXIS_OARG_12_IS_ASYNC,M_AXIS_OARG_11_IS_ASYNC,M_AXIS_OARG_10_IS_ASYNC,M_AXIS_OARG_9_IS_ASYNC,M_AXIS_OARG_8_IS_ASYNC,M_AXIS_OARG_7_IS_ASYNC,M_AXIS_OARG_6_IS_ASYNC,M_AXIS_OARG_5_IS_ASYNC,M_AXIS_OARG_4_IS_ASYNC,M_AXIS_OARG_3_IS_ASYNC,M_AXIS_OARG_2_IS_ASYNC,M_AXIS_OARG_1_IS_ASYNC,M_AXIS_OARG_0_IS_ASYNC};
    localparam [(C_MAX_OUTPUT_AXISs*32)-1:0] C_GEN_TLAST_BIT_ARRAY = {M_AXIS_OARG_127_GEN_TLAST,M_AXIS_OARG_126_GEN_TLAST,M_AXIS_OARG_125_GEN_TLAST,M_AXIS_OARG_124_GEN_TLAST,M_AXIS_OARG_123_GEN_TLAST,M_AXIS_OARG_122_GEN_TLAST,M_AXIS_OARG_121_GEN_TLAST,M_AXIS_OARG_120_GEN_TLAST,M_AXIS_OARG_119_GEN_TLAST,M_AXIS_OARG_118_GEN_TLAST,M_AXIS_OARG_117_GEN_TLAST,M_AXIS_OARG_116_GEN_TLAST,M_AXIS_OARG_115_GEN_TLAST,M_AXIS_OARG_114_GEN_TLAST,M_AXIS_OARG_113_GEN_TLAST,M_AXIS_OARG_112_GEN_TLAST,M_AXIS_OARG_111_GEN_TLAST,M_AXIS_OARG_110_GEN_TLAST,M_AXIS_OARG_109_GEN_TLAST,M_AXIS_OARG_108_GEN_TLAST,M_AXIS_OARG_107_GEN_TLAST,M_AXIS_OARG_106_GEN_TLAST,M_AXIS_OARG_105_GEN_TLAST,M_AXIS_OARG_104_GEN_TLAST,M_AXIS_OARG_103_GEN_TLAST,M_AXIS_OARG_102_GEN_TLAST,M_AXIS_OARG_101_GEN_TLAST,M_AXIS_OARG_100_GEN_TLAST,M_AXIS_OARG_99_GEN_TLAST,M_AXIS_OARG_98_GEN_TLAST,M_AXIS_OARG_97_GEN_TLAST,M_AXIS_OARG_96_GEN_TLAST,M_AXIS_OARG_95_GEN_TLAST,M_AXIS_OARG_94_GEN_TLAST,M_AXIS_OARG_93_GEN_TLAST,M_AXIS_OARG_92_GEN_TLAST,M_AXIS_OARG_91_GEN_TLAST,M_AXIS_OARG_90_GEN_TLAST,M_AXIS_OARG_89_GEN_TLAST,M_AXIS_OARG_88_GEN_TLAST,M_AXIS_OARG_87_GEN_TLAST,M_AXIS_OARG_86_GEN_TLAST,M_AXIS_OARG_85_GEN_TLAST,M_AXIS_OARG_84_GEN_TLAST,M_AXIS_OARG_83_GEN_TLAST,M_AXIS_OARG_82_GEN_TLAST,M_AXIS_OARG_81_GEN_TLAST,M_AXIS_OARG_80_GEN_TLAST,M_AXIS_OARG_79_GEN_TLAST,M_AXIS_OARG_78_GEN_TLAST,M_AXIS_OARG_77_GEN_TLAST,M_AXIS_OARG_76_GEN_TLAST,M_AXIS_OARG_75_GEN_TLAST,M_AXIS_OARG_74_GEN_TLAST,M_AXIS_OARG_73_GEN_TLAST,M_AXIS_OARG_72_GEN_TLAST,M_AXIS_OARG_71_GEN_TLAST,M_AXIS_OARG_70_GEN_TLAST,M_AXIS_OARG_69_GEN_TLAST,M_AXIS_OARG_68_GEN_TLAST,M_AXIS_OARG_67_GEN_TLAST,M_AXIS_OARG_66_GEN_TLAST,M_AXIS_OARG_65_GEN_TLAST,M_AXIS_OARG_64_GEN_TLAST,M_AXIS_OARG_63_GEN_TLAST,M_AXIS_OARG_62_GEN_TLAST,M_AXIS_OARG_61_GEN_TLAST,M_AXIS_OARG_60_GEN_TLAST,M_AXIS_OARG_59_GEN_TLAST,M_AXIS_OARG_58_GEN_TLAST,M_AXIS_OARG_57_GEN_TLAST,M_AXIS_OARG_56_GEN_TLAST,M_AXIS_OARG_55_GEN_TLAST,M_AXIS_OARG_54_GEN_TLAST,M_AXIS_OARG_53_GEN_TLAST,M_AXIS_OARG_52_GEN_TLAST,M_AXIS_OARG_51_GEN_TLAST,M_AXIS_OARG_50_GEN_TLAST,M_AXIS_OARG_49_GEN_TLAST,M_AXIS_OARG_48_GEN_TLAST,M_AXIS_OARG_47_GEN_TLAST,M_AXIS_OARG_46_GEN_TLAST,M_AXIS_OARG_45_GEN_TLAST,M_AXIS_OARG_44_GEN_TLAST,M_AXIS_OARG_43_GEN_TLAST,M_AXIS_OARG_42_GEN_TLAST,M_AXIS_OARG_41_GEN_TLAST,M_AXIS_OARG_40_GEN_TLAST,M_AXIS_OARG_39_GEN_TLAST,M_AXIS_OARG_38_GEN_TLAST,M_AXIS_OARG_37_GEN_TLAST,M_AXIS_OARG_36_GEN_TLAST,M_AXIS_OARG_35_GEN_TLAST,M_AXIS_OARG_34_GEN_TLAST,M_AXIS_OARG_33_GEN_TLAST,M_AXIS_OARG_32_GEN_TLAST,M_AXIS_OARG_31_GEN_TLAST,M_AXIS_OARG_30_GEN_TLAST,M_AXIS_OARG_29_GEN_TLAST,M_AXIS_OARG_28_GEN_TLAST,M_AXIS_OARG_27_GEN_TLAST,M_AXIS_OARG_26_GEN_TLAST,M_AXIS_OARG_25_GEN_TLAST,M_AXIS_OARG_24_GEN_TLAST,M_AXIS_OARG_23_GEN_TLAST,M_AXIS_OARG_22_GEN_TLAST,M_AXIS_OARG_21_GEN_TLAST,M_AXIS_OARG_20_GEN_TLAST,M_AXIS_OARG_19_GEN_TLAST,M_AXIS_OARG_18_GEN_TLAST,M_AXIS_OARG_17_GEN_TLAST,M_AXIS_OARG_16_GEN_TLAST,M_AXIS_OARG_15_GEN_TLAST,M_AXIS_OARG_14_GEN_TLAST,M_AXIS_OARG_13_GEN_TLAST,M_AXIS_OARG_12_GEN_TLAST,M_AXIS_OARG_11_GEN_TLAST,M_AXIS_OARG_10_GEN_TLAST,M_AXIS_OARG_9_GEN_TLAST,M_AXIS_OARG_8_GEN_TLAST,M_AXIS_OARG_7_GEN_TLAST,M_AXIS_OARG_6_GEN_TLAST,M_AXIS_OARG_5_GEN_TLAST,M_AXIS_OARG_4_GEN_TLAST,M_AXIS_OARG_3_GEN_TLAST,M_AXIS_OARG_2_GEN_TLAST,M_AXIS_OARG_1_GEN_TLAST,M_AXIS_OARG_0_GEN_TLAST};
    
    wire [C_MAX_OUTPUT_AXISs-1:0] axis_clk;
    wire [C_MAX_OUTPUT_AXISs-1:0] axis_rst;
    
    wire [C_MAX_OUTPUT_AXISs-1:0] dm_tlast;
    wire [C_MAX_OUTPUT_AXISs-1:0] dm_tvalid;
    wire [C_MAX_OUTPUT_AXISs-1:0] dm_tready;
    wire [C_MAX_BIT_WIDTH/8-1:0] dm_tkeep [C_NUM_OUTPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] dm_tstrb [C_NUM_OUTPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0] dm_tdata [C_MAX_OUTPUT_AXISs-1:0];
    
    wire [C_MAX_OUTPUT_AXISs-1:0] buf_tlast;
    wire [C_MAX_OUTPUT_AXISs-1:0] buf_tvalid;
    wire [C_MAX_OUTPUT_AXISs-1:0] buf_tready;
    wire [C_MAX_BIT_WIDTH-1:0] buf_tdata [C_MAX_OUTPUT_AXISs-1:0];
    
    wire [C_MAX_OUTPUT_AXISs-1:0] dwconv_tlast;
    wire [C_MAX_OUTPUT_AXISs-1:0] dwconv_tvalid;
    wire [C_MAX_OUTPUT_AXISs-1:0] dwconv_tready;
    wire [C_MAX_BIT_WIDTH/8-1:0] dwconv_tkeep [C_NUM_OUTPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] dwconv_tstrb [C_NUM_OUTPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0] dwconv_tdata [C_MAX_OUTPUT_AXISs-1:0];
    
    wire [C_MAX_OUTPUT_AXISs-1:0] ap_tlast;
    wire [C_MAX_OUTPUT_AXISs-1:0] ap_tvalid;
    wire [C_MAX_OUTPUT_AXISs-1:0] ap_tready;
    wire [C_MAX_BIT_WIDTH/8-1:0] ap_tkeep [C_NUM_OUTPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] ap_tstrb [C_NUM_OUTPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0] ap_tdata [C_MAX_OUTPUT_AXISs-1:0];
        
    //assign inputs to buses, and buses to outputs
    generate
        if(C_NUM_OUTPUT_AXISs > 0) begin
            assign axis_clk[0] = m_axis_oarg_0_aclk;
            assign axis_rst[0] = m_axis_oarg_0_aresetn;
            assign dm_tready[0] = m_axis_oarg_0_tready;
            assign m_axis_oarg_0_tlast = dm_tlast[0];
            assign m_axis_oarg_0_tvalid = dm_tvalid[0];
            assign m_axis_oarg_0_tkeep = dm_tkeep[0][M_AXIS_OARG_0_DMWIDTH/8-1:0];
            assign m_axis_oarg_0_tstrb = dm_tstrb[0][M_AXIS_OARG_0_DMWIDTH/8-1:0];
            assign m_axis_oarg_0_tdata = dm_tdata[0][M_AXIS_OARG_0_DMWIDTH-1:0];
            assign ap_axis_oarg_0_tready = ap_tready[0];
            assign ap_tlast[0] = ap_axis_oarg_0_tlast;
            assign ap_tvalid[0] = ap_axis_oarg_0_tvalid;
            assign ap_tdata[0][M_AXIS_OARG_0_WIDTH-1:0] = ap_axis_oarg_0_tdata;
            assign ap_tkeep[0] = {M_AXIS_OARG_0_WIDTH/8{1'b1}};
            assign ap_tstrb[0] = {M_AXIS_OARG_0_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 1) begin
            assign axis_clk[1] = m_axis_oarg_1_aclk;
            assign axis_rst[1] = m_axis_oarg_1_aresetn;
            assign dm_tready[1] = m_axis_oarg_1_tready;
            assign m_axis_oarg_1_tlast = dm_tlast[1];
            assign m_axis_oarg_1_tvalid = dm_tvalid[1];
            assign m_axis_oarg_1_tkeep = dm_tkeep[1][M_AXIS_OARG_1_DMWIDTH/8-1:0];
            assign m_axis_oarg_1_tstrb = dm_tstrb[1][M_AXIS_OARG_1_DMWIDTH/8-1:0];
            assign m_axis_oarg_1_tdata = dm_tdata[1][M_AXIS_OARG_1_DMWIDTH-1:0];
            assign ap_axis_oarg_1_tready = ap_tready[1];
            assign ap_tlast[1] = ap_axis_oarg_1_tlast;
            assign ap_tvalid[1] = ap_axis_oarg_1_tvalid;
            assign ap_tdata[1][M_AXIS_OARG_1_WIDTH-1:0] = ap_axis_oarg_1_tdata;
            assign ap_tkeep[1] = {M_AXIS_OARG_1_WIDTH/8{1'b1}};
            assign ap_tstrb[1] = {M_AXIS_OARG_1_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 2) begin
            assign axis_clk[2] = m_axis_oarg_2_aclk;
            assign axis_rst[2] = m_axis_oarg_2_aresetn;
            assign dm_tready[2] = m_axis_oarg_2_tready;
            assign m_axis_oarg_2_tlast = dm_tlast[2];
            assign m_axis_oarg_2_tvalid = dm_tvalid[2];
            assign m_axis_oarg_2_tkeep = dm_tkeep[2][M_AXIS_OARG_2_DMWIDTH/8-1:0];
            assign m_axis_oarg_2_tstrb = dm_tstrb[2][M_AXIS_OARG_2_DMWIDTH/8-1:0];
            assign m_axis_oarg_2_tdata = dm_tdata[2][M_AXIS_OARG_2_DMWIDTH-1:0];
            assign ap_axis_oarg_2_tready = ap_tready[2];
            assign ap_tlast[2] = ap_axis_oarg_2_tlast;
            assign ap_tvalid[2] = ap_axis_oarg_2_tvalid;
            assign ap_tdata[2][M_AXIS_OARG_2_WIDTH-1:0] = ap_axis_oarg_2_tdata;
            assign ap_tkeep[2] = {M_AXIS_OARG_2_WIDTH/8{1'b1}};
            assign ap_tstrb[2] = {M_AXIS_OARG_2_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 3) begin
            assign axis_clk[3] = m_axis_oarg_3_aclk;
            assign axis_rst[3] = m_axis_oarg_3_aresetn;
            assign dm_tready[3] = m_axis_oarg_3_tready;
            assign m_axis_oarg_3_tlast = dm_tlast[3];
            assign m_axis_oarg_3_tvalid = dm_tvalid[3];
            assign m_axis_oarg_3_tkeep = dm_tkeep[3][M_AXIS_OARG_3_DMWIDTH/8-1:0];
            assign m_axis_oarg_3_tstrb = dm_tstrb[3][M_AXIS_OARG_3_DMWIDTH/8-1:0];
            assign m_axis_oarg_3_tdata = dm_tdata[3][M_AXIS_OARG_3_DMWIDTH-1:0];
            assign ap_axis_oarg_3_tready = ap_tready[3];
            assign ap_tlast[3] = ap_axis_oarg_3_tlast;
            assign ap_tvalid[3] = ap_axis_oarg_3_tvalid;
            assign ap_tdata[3][M_AXIS_OARG_3_WIDTH-1:0] = ap_axis_oarg_3_tdata;
            assign ap_tkeep[3] = {M_AXIS_OARG_3_WIDTH/8{1'b1}};
            assign ap_tstrb[3] = {M_AXIS_OARG_3_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 4) begin
            assign axis_clk[4] = m_axis_oarg_4_aclk;
            assign axis_rst[4] = m_axis_oarg_4_aresetn;
            assign dm_tready[4] = m_axis_oarg_4_tready;
            assign m_axis_oarg_4_tlast = dm_tlast[4];
            assign m_axis_oarg_4_tvalid = dm_tvalid[4];
            assign m_axis_oarg_4_tkeep = dm_tkeep[4][M_AXIS_OARG_4_DMWIDTH/8-1:0];
            assign m_axis_oarg_4_tstrb = dm_tstrb[4][M_AXIS_OARG_4_DMWIDTH/8-1:0];
            assign m_axis_oarg_4_tdata = dm_tdata[4][M_AXIS_OARG_4_DMWIDTH-1:0];
            assign ap_axis_oarg_4_tready = ap_tready[4];
            assign ap_tlast[4] = ap_axis_oarg_4_tlast;
            assign ap_tvalid[4] = ap_axis_oarg_4_tvalid;
            assign ap_tdata[4][M_AXIS_OARG_4_WIDTH-1:0] = ap_axis_oarg_4_tdata;
            assign ap_tkeep[4] = {M_AXIS_OARG_4_WIDTH/8{1'b1}};
            assign ap_tstrb[4] = {M_AXIS_OARG_4_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 5) begin
            assign axis_clk[5] = m_axis_oarg_5_aclk;
            assign axis_rst[5] = m_axis_oarg_5_aresetn;
            assign dm_tready[5] = m_axis_oarg_5_tready;
            assign m_axis_oarg_5_tlast = dm_tlast[5];
            assign m_axis_oarg_5_tvalid = dm_tvalid[5];
            assign m_axis_oarg_5_tkeep = dm_tkeep[5][M_AXIS_OARG_5_DMWIDTH/8-1:0];
            assign m_axis_oarg_5_tstrb = dm_tstrb[5][M_AXIS_OARG_5_DMWIDTH/8-1:0];
            assign m_axis_oarg_5_tdata = dm_tdata[5][M_AXIS_OARG_5_DMWIDTH-1:0];
            assign ap_axis_oarg_5_tready = ap_tready[5];
            assign ap_tlast[5] = ap_axis_oarg_5_tlast;
            assign ap_tvalid[5] = ap_axis_oarg_5_tvalid;
            assign ap_tdata[5][M_AXIS_OARG_5_WIDTH-1:0] = ap_axis_oarg_5_tdata;
            assign ap_tkeep[5] = {M_AXIS_OARG_5_WIDTH/8{1'b1}};
            assign ap_tstrb[5] = {M_AXIS_OARG_5_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 6) begin
            assign axis_clk[6] = m_axis_oarg_6_aclk;
            assign axis_rst[6] = m_axis_oarg_6_aresetn;
            assign dm_tready[6] = m_axis_oarg_6_tready;
            assign m_axis_oarg_6_tlast = dm_tlast[6];
            assign m_axis_oarg_6_tvalid = dm_tvalid[6];
            assign m_axis_oarg_6_tkeep = dm_tkeep[6][M_AXIS_OARG_6_DMWIDTH/8-1:0];
            assign m_axis_oarg_6_tstrb = dm_tstrb[6][M_AXIS_OARG_6_DMWIDTH/8-1:0];
            assign m_axis_oarg_6_tdata = dm_tdata[6][M_AXIS_OARG_6_DMWIDTH-1:0];
            assign ap_axis_oarg_6_tready = ap_tready[6];
            assign ap_tlast[6] = ap_axis_oarg_6_tlast;
            assign ap_tvalid[6] = ap_axis_oarg_6_tvalid;
            assign ap_tdata[6][M_AXIS_OARG_6_WIDTH-1:0] = ap_axis_oarg_6_tdata;
            assign ap_tkeep[6] = {M_AXIS_OARG_6_WIDTH/8{1'b1}};
            assign ap_tstrb[6] = {M_AXIS_OARG_6_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 7) begin
            assign axis_clk[7] = m_axis_oarg_7_aclk;
            assign axis_rst[7] = m_axis_oarg_7_aresetn;
            assign dm_tready[7] = m_axis_oarg_7_tready;
            assign m_axis_oarg_7_tlast = dm_tlast[7];
            assign m_axis_oarg_7_tvalid = dm_tvalid[7];
            assign m_axis_oarg_7_tkeep = dm_tkeep[7][M_AXIS_OARG_7_DMWIDTH/8-1:0];
            assign m_axis_oarg_7_tstrb = dm_tstrb[7][M_AXIS_OARG_7_DMWIDTH/8-1:0];
            assign m_axis_oarg_7_tdata = dm_tdata[7][M_AXIS_OARG_7_DMWIDTH-1:0];
            assign ap_axis_oarg_7_tready = ap_tready[7];
            assign ap_tlast[7] = ap_axis_oarg_7_tlast;
            assign ap_tvalid[7] = ap_axis_oarg_7_tvalid;
            assign ap_tdata[7][M_AXIS_OARG_7_WIDTH-1:0] = ap_axis_oarg_7_tdata;
            assign ap_tkeep[7] = {M_AXIS_OARG_7_WIDTH/8{1'b1}};
            assign ap_tstrb[7] = {M_AXIS_OARG_7_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 8) begin
            assign axis_clk[8] = m_axis_oarg_8_aclk;
            assign axis_rst[8] = m_axis_oarg_8_aresetn;
            assign dm_tready[8] = m_axis_oarg_8_tready;
            assign m_axis_oarg_8_tlast = dm_tlast[8];
            assign m_axis_oarg_8_tvalid = dm_tvalid[8];
            assign m_axis_oarg_8_tkeep = dm_tkeep[8][M_AXIS_OARG_8_DMWIDTH/8-1:0];
            assign m_axis_oarg_8_tstrb = dm_tstrb[8][M_AXIS_OARG_8_DMWIDTH/8-1:0];
            assign m_axis_oarg_8_tdata = dm_tdata[8][M_AXIS_OARG_8_DMWIDTH-1:0];
            assign ap_axis_oarg_8_tready = ap_tready[8];
            assign ap_tlast[8] = ap_axis_oarg_8_tlast;
            assign ap_tvalid[8] = ap_axis_oarg_8_tvalid;
            assign ap_tdata[8][M_AXIS_OARG_8_WIDTH-1:0] = ap_axis_oarg_8_tdata;
            assign ap_tkeep[8] = {M_AXIS_OARG_8_WIDTH/8{1'b1}};
            assign ap_tstrb[8] = {M_AXIS_OARG_8_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 9) begin
            assign axis_clk[9] = m_axis_oarg_9_aclk;
            assign axis_rst[9] = m_axis_oarg_9_aresetn;
            assign dm_tready[9] = m_axis_oarg_9_tready;
            assign m_axis_oarg_9_tlast = dm_tlast[9];
            assign m_axis_oarg_9_tvalid = dm_tvalid[9];
            assign m_axis_oarg_9_tkeep = dm_tkeep[9][M_AXIS_OARG_9_DMWIDTH/8-1:0];
            assign m_axis_oarg_9_tstrb = dm_tstrb[9][M_AXIS_OARG_9_DMWIDTH/8-1:0];
            assign m_axis_oarg_9_tdata = dm_tdata[9][M_AXIS_OARG_9_DMWIDTH-1:0];
            assign ap_axis_oarg_9_tready = ap_tready[9];
            assign ap_tlast[9] = ap_axis_oarg_9_tlast;
            assign ap_tvalid[9] = ap_axis_oarg_9_tvalid;
            assign ap_tdata[9][M_AXIS_OARG_9_WIDTH-1:0] = ap_axis_oarg_9_tdata;
            assign ap_tkeep[9] = {M_AXIS_OARG_9_WIDTH/8{1'b1}};
            assign ap_tstrb[9] = {M_AXIS_OARG_9_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 10) begin
            assign axis_clk[10] = m_axis_oarg_10_aclk;
            assign axis_rst[10] = m_axis_oarg_10_aresetn;
            assign dm_tready[10] = m_axis_oarg_10_tready;
            assign m_axis_oarg_10_tlast = dm_tlast[10];
            assign m_axis_oarg_10_tvalid = dm_tvalid[10];
            assign m_axis_oarg_10_tkeep = dm_tkeep[10][M_AXIS_OARG_10_DMWIDTH/8-1:0];
            assign m_axis_oarg_10_tstrb = dm_tstrb[10][M_AXIS_OARG_10_DMWIDTH/8-1:0];
            assign m_axis_oarg_10_tdata = dm_tdata[10][M_AXIS_OARG_10_DMWIDTH-1:0];
            assign ap_axis_oarg_10_tready = ap_tready[10];
            assign ap_tlast[10] = ap_axis_oarg_10_tlast;
            assign ap_tvalid[10] = ap_axis_oarg_10_tvalid;
            assign ap_tdata[10][M_AXIS_OARG_10_WIDTH-1:0] = ap_axis_oarg_10_tdata;
            assign ap_tkeep[10] = {M_AXIS_OARG_10_WIDTH/8{1'b1}};
            assign ap_tstrb[10] = {M_AXIS_OARG_10_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 11) begin
            assign axis_clk[11] = m_axis_oarg_11_aclk;
            assign axis_rst[11] = m_axis_oarg_11_aresetn;
            assign dm_tready[11] = m_axis_oarg_11_tready;
            assign m_axis_oarg_11_tlast = dm_tlast[11];
            assign m_axis_oarg_11_tvalid = dm_tvalid[11];
            assign m_axis_oarg_11_tkeep = dm_tkeep[11][M_AXIS_OARG_11_DMWIDTH/8-1:0];
            assign m_axis_oarg_11_tstrb = dm_tstrb[11][M_AXIS_OARG_11_DMWIDTH/8-1:0];
            assign m_axis_oarg_11_tdata = dm_tdata[11][M_AXIS_OARG_11_DMWIDTH-1:0];
            assign ap_axis_oarg_11_tready = ap_tready[11];
            assign ap_tlast[11] = ap_axis_oarg_11_tlast;
            assign ap_tvalid[11] = ap_axis_oarg_11_tvalid;
            assign ap_tdata[11][M_AXIS_OARG_11_WIDTH-1:0] = ap_axis_oarg_11_tdata;
            assign ap_tkeep[11] = {M_AXIS_OARG_11_WIDTH/8{1'b1}};
            assign ap_tstrb[11] = {M_AXIS_OARG_11_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 12) begin
            assign axis_clk[12] = m_axis_oarg_12_aclk;
            assign axis_rst[12] = m_axis_oarg_12_aresetn;
            assign dm_tready[12] = m_axis_oarg_12_tready;
            assign m_axis_oarg_12_tlast = dm_tlast[12];
            assign m_axis_oarg_12_tvalid = dm_tvalid[12];
            assign m_axis_oarg_12_tkeep = dm_tkeep[12][M_AXIS_OARG_12_DMWIDTH/8-1:0];
            assign m_axis_oarg_12_tstrb = dm_tstrb[12][M_AXIS_OARG_12_DMWIDTH/8-1:0];
            assign m_axis_oarg_12_tdata = dm_tdata[12][M_AXIS_OARG_12_DMWIDTH-1:0];
            assign ap_axis_oarg_12_tready = ap_tready[12];
            assign ap_tlast[12] = ap_axis_oarg_12_tlast;
            assign ap_tvalid[12] = ap_axis_oarg_12_tvalid;
            assign ap_tdata[12][M_AXIS_OARG_12_WIDTH-1:0] = ap_axis_oarg_12_tdata;
            assign ap_tkeep[12] = {M_AXIS_OARG_12_WIDTH/8{1'b1}};
            assign ap_tstrb[12] = {M_AXIS_OARG_12_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 13) begin
            assign axis_clk[13] = m_axis_oarg_13_aclk;
            assign axis_rst[13] = m_axis_oarg_13_aresetn;
            assign dm_tready[13] = m_axis_oarg_13_tready;
            assign m_axis_oarg_13_tlast = dm_tlast[13];
            assign m_axis_oarg_13_tvalid = dm_tvalid[13];
            assign m_axis_oarg_13_tkeep = dm_tkeep[13][M_AXIS_OARG_13_DMWIDTH/8-1:0];
            assign m_axis_oarg_13_tstrb = dm_tstrb[13][M_AXIS_OARG_13_DMWIDTH/8-1:0];
            assign m_axis_oarg_13_tdata = dm_tdata[13][M_AXIS_OARG_13_DMWIDTH-1:0];
            assign ap_axis_oarg_13_tready = ap_tready[13];
            assign ap_tlast[13] = ap_axis_oarg_13_tlast;
            assign ap_tvalid[13] = ap_axis_oarg_13_tvalid;
            assign ap_tdata[13][M_AXIS_OARG_13_WIDTH-1:0] = ap_axis_oarg_13_tdata;
            assign ap_tkeep[13] = {M_AXIS_OARG_13_WIDTH/8{1'b1}};
            assign ap_tstrb[13] = {M_AXIS_OARG_13_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 14) begin
            assign axis_clk[14] = m_axis_oarg_14_aclk;
            assign axis_rst[14] = m_axis_oarg_14_aresetn;
            assign dm_tready[14] = m_axis_oarg_14_tready;
            assign m_axis_oarg_14_tlast = dm_tlast[14];
            assign m_axis_oarg_14_tvalid = dm_tvalid[14];
            assign m_axis_oarg_14_tkeep = dm_tkeep[14][M_AXIS_OARG_14_DMWIDTH/8-1:0];
            assign m_axis_oarg_14_tstrb = dm_tstrb[14][M_AXIS_OARG_14_DMWIDTH/8-1:0];
            assign m_axis_oarg_14_tdata = dm_tdata[14][M_AXIS_OARG_14_DMWIDTH-1:0];
            assign ap_axis_oarg_14_tready = ap_tready[14];
            assign ap_tlast[14] = ap_axis_oarg_14_tlast;
            assign ap_tvalid[14] = ap_axis_oarg_14_tvalid;
            assign ap_tdata[14][M_AXIS_OARG_14_WIDTH-1:0] = ap_axis_oarg_14_tdata;
            assign ap_tkeep[14] = {M_AXIS_OARG_14_WIDTH/8{1'b1}};
            assign ap_tstrb[14] = {M_AXIS_OARG_14_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 15) begin
            assign axis_clk[15] = m_axis_oarg_15_aclk;
            assign axis_rst[15] = m_axis_oarg_15_aresetn;
            assign dm_tready[15] = m_axis_oarg_15_tready;
            assign m_axis_oarg_15_tlast = dm_tlast[15];
            assign m_axis_oarg_15_tvalid = dm_tvalid[15];
            assign m_axis_oarg_15_tkeep = dm_tkeep[15][M_AXIS_OARG_15_DMWIDTH/8-1:0];
            assign m_axis_oarg_15_tstrb = dm_tstrb[15][M_AXIS_OARG_15_DMWIDTH/8-1:0];
            assign m_axis_oarg_15_tdata = dm_tdata[15][M_AXIS_OARG_15_DMWIDTH-1:0];
            assign ap_axis_oarg_15_tready = ap_tready[15];
            assign ap_tlast[15] = ap_axis_oarg_15_tlast;
            assign ap_tvalid[15] = ap_axis_oarg_15_tvalid;
            assign ap_tdata[15][M_AXIS_OARG_15_WIDTH-1:0] = ap_axis_oarg_15_tdata;
            assign ap_tkeep[15] = {M_AXIS_OARG_15_WIDTH/8{1'b1}};
            assign ap_tstrb[15] = {M_AXIS_OARG_15_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 16) begin
            assign axis_clk[16] = m_axis_oarg_16_aclk;
            assign axis_rst[16] = m_axis_oarg_16_aresetn;
            assign dm_tready[16] = m_axis_oarg_16_tready;
            assign m_axis_oarg_16_tlast = dm_tlast[16];
            assign m_axis_oarg_16_tvalid = dm_tvalid[16];
            assign m_axis_oarg_16_tkeep = dm_tkeep[16][M_AXIS_OARG_16_DMWIDTH/8-1:0];
            assign m_axis_oarg_16_tstrb = dm_tstrb[16][M_AXIS_OARG_16_DMWIDTH/8-1:0];
            assign m_axis_oarg_16_tdata = dm_tdata[16][M_AXIS_OARG_16_DMWIDTH-1:0];
            assign ap_axis_oarg_16_tready = ap_tready[16];
            assign ap_tlast[16] = ap_axis_oarg_16_tlast;
            assign ap_tvalid[16] = ap_axis_oarg_16_tvalid;
            assign ap_tdata[16][M_AXIS_OARG_16_WIDTH-1:0] = ap_axis_oarg_16_tdata;
            assign ap_tkeep[16] = {M_AXIS_OARG_16_WIDTH/8{1'b1}};
            assign ap_tstrb[16] = {M_AXIS_OARG_16_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 17) begin
            assign axis_clk[17] = m_axis_oarg_17_aclk;
            assign axis_rst[17] = m_axis_oarg_17_aresetn;
            assign dm_tready[17] = m_axis_oarg_17_tready;
            assign m_axis_oarg_17_tlast = dm_tlast[17];
            assign m_axis_oarg_17_tvalid = dm_tvalid[17];
            assign m_axis_oarg_17_tkeep = dm_tkeep[17][M_AXIS_OARG_17_DMWIDTH/8-1:0];
            assign m_axis_oarg_17_tstrb = dm_tstrb[17][M_AXIS_OARG_17_DMWIDTH/8-1:0];
            assign m_axis_oarg_17_tdata = dm_tdata[17][M_AXIS_OARG_17_DMWIDTH-1:0];
            assign ap_axis_oarg_17_tready = ap_tready[17];
            assign ap_tlast[17] = ap_axis_oarg_17_tlast;
            assign ap_tvalid[17] = ap_axis_oarg_17_tvalid;
            assign ap_tdata[17][M_AXIS_OARG_17_WIDTH-1:0] = ap_axis_oarg_17_tdata;
            assign ap_tkeep[17] = {M_AXIS_OARG_17_WIDTH/8{1'b1}};
            assign ap_tstrb[17] = {M_AXIS_OARG_17_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 18) begin
            assign axis_clk[18] = m_axis_oarg_18_aclk;
            assign axis_rst[18] = m_axis_oarg_18_aresetn;
            assign dm_tready[18] = m_axis_oarg_18_tready;
            assign m_axis_oarg_18_tlast = dm_tlast[18];
            assign m_axis_oarg_18_tvalid = dm_tvalid[18];
            assign m_axis_oarg_18_tkeep = dm_tkeep[18][M_AXIS_OARG_18_DMWIDTH/8-1:0];
            assign m_axis_oarg_18_tstrb = dm_tstrb[18][M_AXIS_OARG_18_DMWIDTH/8-1:0];
            assign m_axis_oarg_18_tdata = dm_tdata[18][M_AXIS_OARG_18_DMWIDTH-1:0];
            assign ap_axis_oarg_18_tready = ap_tready[18];
            assign ap_tlast[18] = ap_axis_oarg_18_tlast;
            assign ap_tvalid[18] = ap_axis_oarg_18_tvalid;
            assign ap_tdata[18][M_AXIS_OARG_18_WIDTH-1:0] = ap_axis_oarg_18_tdata;
            assign ap_tkeep[18] = {M_AXIS_OARG_18_WIDTH/8{1'b1}};
            assign ap_tstrb[18] = {M_AXIS_OARG_18_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 19) begin
            assign axis_clk[19] = m_axis_oarg_19_aclk;
            assign axis_rst[19] = m_axis_oarg_19_aresetn;
            assign dm_tready[19] = m_axis_oarg_19_tready;
            assign m_axis_oarg_19_tlast = dm_tlast[19];
            assign m_axis_oarg_19_tvalid = dm_tvalid[19];
            assign m_axis_oarg_19_tkeep = dm_tkeep[19][M_AXIS_OARG_19_DMWIDTH/8-1:0];
            assign m_axis_oarg_19_tstrb = dm_tstrb[19][M_AXIS_OARG_19_DMWIDTH/8-1:0];
            assign m_axis_oarg_19_tdata = dm_tdata[19][M_AXIS_OARG_19_DMWIDTH-1:0];
            assign ap_axis_oarg_19_tready = ap_tready[19];
            assign ap_tlast[19] = ap_axis_oarg_19_tlast;
            assign ap_tvalid[19] = ap_axis_oarg_19_tvalid;
            assign ap_tdata[19][M_AXIS_OARG_19_WIDTH-1:0] = ap_axis_oarg_19_tdata;
            assign ap_tkeep[19] = {M_AXIS_OARG_19_WIDTH/8{1'b1}};
            assign ap_tstrb[19] = {M_AXIS_OARG_19_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 20) begin
            assign axis_clk[20] = m_axis_oarg_20_aclk;
            assign axis_rst[20] = m_axis_oarg_20_aresetn;
            assign dm_tready[20] = m_axis_oarg_20_tready;
            assign m_axis_oarg_20_tlast = dm_tlast[20];
            assign m_axis_oarg_20_tvalid = dm_tvalid[20];
            assign m_axis_oarg_20_tkeep = dm_tkeep[20][M_AXIS_OARG_20_DMWIDTH/8-1:0];
            assign m_axis_oarg_20_tstrb = dm_tstrb[20][M_AXIS_OARG_20_DMWIDTH/8-1:0];
            assign m_axis_oarg_20_tdata = dm_tdata[20][M_AXIS_OARG_20_DMWIDTH-1:0];
            assign ap_axis_oarg_20_tready = ap_tready[20];
            assign ap_tlast[20] = ap_axis_oarg_20_tlast;
            assign ap_tvalid[20] = ap_axis_oarg_20_tvalid;
            assign ap_tdata[20][M_AXIS_OARG_20_WIDTH-1:0] = ap_axis_oarg_20_tdata;
            assign ap_tkeep[20] = {M_AXIS_OARG_20_WIDTH/8{1'b1}};
            assign ap_tstrb[20] = {M_AXIS_OARG_20_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 21) begin
            assign axis_clk[21] = m_axis_oarg_21_aclk;
            assign axis_rst[21] = m_axis_oarg_21_aresetn;
            assign dm_tready[21] = m_axis_oarg_21_tready;
            assign m_axis_oarg_21_tlast = dm_tlast[21];
            assign m_axis_oarg_21_tvalid = dm_tvalid[21];
            assign m_axis_oarg_21_tkeep = dm_tkeep[21][M_AXIS_OARG_21_DMWIDTH/8-1:0];
            assign m_axis_oarg_21_tstrb = dm_tstrb[21][M_AXIS_OARG_21_DMWIDTH/8-1:0];
            assign m_axis_oarg_21_tdata = dm_tdata[21][M_AXIS_OARG_21_DMWIDTH-1:0];
            assign ap_axis_oarg_21_tready = ap_tready[21];
            assign ap_tlast[21] = ap_axis_oarg_21_tlast;
            assign ap_tvalid[21] = ap_axis_oarg_21_tvalid;
            assign ap_tdata[21][M_AXIS_OARG_21_WIDTH-1:0] = ap_axis_oarg_21_tdata;
            assign ap_tkeep[21] = {M_AXIS_OARG_21_WIDTH/8{1'b1}};
            assign ap_tstrb[21] = {M_AXIS_OARG_21_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 22) begin
            assign axis_clk[22] = m_axis_oarg_22_aclk;
            assign axis_rst[22] = m_axis_oarg_22_aresetn;
            assign dm_tready[22] = m_axis_oarg_22_tready;
            assign m_axis_oarg_22_tlast = dm_tlast[22];
            assign m_axis_oarg_22_tvalid = dm_tvalid[22];
            assign m_axis_oarg_22_tkeep = dm_tkeep[22][M_AXIS_OARG_22_DMWIDTH/8-1:0];
            assign m_axis_oarg_22_tstrb = dm_tstrb[22][M_AXIS_OARG_22_DMWIDTH/8-1:0];
            assign m_axis_oarg_22_tdata = dm_tdata[22][M_AXIS_OARG_22_DMWIDTH-1:0];
            assign ap_axis_oarg_22_tready = ap_tready[22];
            assign ap_tlast[22] = ap_axis_oarg_22_tlast;
            assign ap_tvalid[22] = ap_axis_oarg_22_tvalid;
            assign ap_tdata[22][M_AXIS_OARG_22_WIDTH-1:0] = ap_axis_oarg_22_tdata;
            assign ap_tkeep[22] = {M_AXIS_OARG_22_WIDTH/8{1'b1}};
            assign ap_tstrb[22] = {M_AXIS_OARG_22_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 23) begin
            assign axis_clk[23] = m_axis_oarg_23_aclk;
            assign axis_rst[23] = m_axis_oarg_23_aresetn;
            assign dm_tready[23] = m_axis_oarg_23_tready;
            assign m_axis_oarg_23_tlast = dm_tlast[23];
            assign m_axis_oarg_23_tvalid = dm_tvalid[23];
            assign m_axis_oarg_23_tkeep = dm_tkeep[23][M_AXIS_OARG_23_DMWIDTH/8-1:0];
            assign m_axis_oarg_23_tstrb = dm_tstrb[23][M_AXIS_OARG_23_DMWIDTH/8-1:0];
            assign m_axis_oarg_23_tdata = dm_tdata[23][M_AXIS_OARG_23_DMWIDTH-1:0];
            assign ap_axis_oarg_23_tready = ap_tready[23];
            assign ap_tlast[23] = ap_axis_oarg_23_tlast;
            assign ap_tvalid[23] = ap_axis_oarg_23_tvalid;
            assign ap_tdata[23][M_AXIS_OARG_23_WIDTH-1:0] = ap_axis_oarg_23_tdata;
            assign ap_tkeep[23] = {M_AXIS_OARG_23_WIDTH/8{1'b1}};
            assign ap_tstrb[23] = {M_AXIS_OARG_23_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 24) begin
            assign axis_clk[24] = m_axis_oarg_24_aclk;
            assign axis_rst[24] = m_axis_oarg_24_aresetn;
            assign dm_tready[24] = m_axis_oarg_24_tready;
            assign m_axis_oarg_24_tlast = dm_tlast[24];
            assign m_axis_oarg_24_tvalid = dm_tvalid[24];
            assign m_axis_oarg_24_tkeep = dm_tkeep[24][M_AXIS_OARG_24_DMWIDTH/8-1:0];
            assign m_axis_oarg_24_tstrb = dm_tstrb[24][M_AXIS_OARG_24_DMWIDTH/8-1:0];
            assign m_axis_oarg_24_tdata = dm_tdata[24][M_AXIS_OARG_24_DMWIDTH-1:0];
            assign ap_axis_oarg_24_tready = ap_tready[24];
            assign ap_tlast[24] = ap_axis_oarg_24_tlast;
            assign ap_tvalid[24] = ap_axis_oarg_24_tvalid;
            assign ap_tdata[24][M_AXIS_OARG_24_WIDTH-1:0] = ap_axis_oarg_24_tdata;
            assign ap_tkeep[24] = {M_AXIS_OARG_24_WIDTH/8{1'b1}};
            assign ap_tstrb[24] = {M_AXIS_OARG_24_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 25) begin
            assign axis_clk[25] = m_axis_oarg_25_aclk;
            assign axis_rst[25] = m_axis_oarg_25_aresetn;
            assign dm_tready[25] = m_axis_oarg_25_tready;
            assign m_axis_oarg_25_tlast = dm_tlast[25];
            assign m_axis_oarg_25_tvalid = dm_tvalid[25];
            assign m_axis_oarg_25_tkeep = dm_tkeep[25][M_AXIS_OARG_25_DMWIDTH/8-1:0];
            assign m_axis_oarg_25_tstrb = dm_tstrb[25][M_AXIS_OARG_25_DMWIDTH/8-1:0];
            assign m_axis_oarg_25_tdata = dm_tdata[25][M_AXIS_OARG_25_DMWIDTH-1:0];
            assign ap_axis_oarg_25_tready = ap_tready[25];
            assign ap_tlast[25] = ap_axis_oarg_25_tlast;
            assign ap_tvalid[25] = ap_axis_oarg_25_tvalid;
            assign ap_tdata[25][M_AXIS_OARG_25_WIDTH-1:0] = ap_axis_oarg_25_tdata;
            assign ap_tkeep[25] = {M_AXIS_OARG_25_WIDTH/8{1'b1}};
            assign ap_tstrb[25] = {M_AXIS_OARG_25_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 26) begin
            assign axis_clk[26] = m_axis_oarg_26_aclk;
            assign axis_rst[26] = m_axis_oarg_26_aresetn;
            assign dm_tready[26] = m_axis_oarg_26_tready;
            assign m_axis_oarg_26_tlast = dm_tlast[26];
            assign m_axis_oarg_26_tvalid = dm_tvalid[26];
            assign m_axis_oarg_26_tkeep = dm_tkeep[26][M_AXIS_OARG_26_DMWIDTH/8-1:0];
            assign m_axis_oarg_26_tstrb = dm_tstrb[26][M_AXIS_OARG_26_DMWIDTH/8-1:0];
            assign m_axis_oarg_26_tdata = dm_tdata[26][M_AXIS_OARG_26_DMWIDTH-1:0];
            assign ap_axis_oarg_26_tready = ap_tready[26];
            assign ap_tlast[26] = ap_axis_oarg_26_tlast;
            assign ap_tvalid[26] = ap_axis_oarg_26_tvalid;
            assign ap_tdata[26][M_AXIS_OARG_26_WIDTH-1:0] = ap_axis_oarg_26_tdata;
            assign ap_tkeep[26] = {M_AXIS_OARG_26_WIDTH/8{1'b1}};
            assign ap_tstrb[26] = {M_AXIS_OARG_26_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 27) begin
            assign axis_clk[27] = m_axis_oarg_27_aclk;
            assign axis_rst[27] = m_axis_oarg_27_aresetn;
            assign dm_tready[27] = m_axis_oarg_27_tready;
            assign m_axis_oarg_27_tlast = dm_tlast[27];
            assign m_axis_oarg_27_tvalid = dm_tvalid[27];
            assign m_axis_oarg_27_tkeep = dm_tkeep[27][M_AXIS_OARG_27_DMWIDTH/8-1:0];
            assign m_axis_oarg_27_tstrb = dm_tstrb[27][M_AXIS_OARG_27_DMWIDTH/8-1:0];
            assign m_axis_oarg_27_tdata = dm_tdata[27][M_AXIS_OARG_27_DMWIDTH-1:0];
            assign ap_axis_oarg_27_tready = ap_tready[27];
            assign ap_tlast[27] = ap_axis_oarg_27_tlast;
            assign ap_tvalid[27] = ap_axis_oarg_27_tvalid;
            assign ap_tdata[27][M_AXIS_OARG_27_WIDTH-1:0] = ap_axis_oarg_27_tdata;
            assign ap_tkeep[27] = {M_AXIS_OARG_27_WIDTH/8{1'b1}};
            assign ap_tstrb[27] = {M_AXIS_OARG_27_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 28) begin
            assign axis_clk[28] = m_axis_oarg_28_aclk;
            assign axis_rst[28] = m_axis_oarg_28_aresetn;
            assign dm_tready[28] = m_axis_oarg_28_tready;
            assign m_axis_oarg_28_tlast = dm_tlast[28];
            assign m_axis_oarg_28_tvalid = dm_tvalid[28];
            assign m_axis_oarg_28_tkeep = dm_tkeep[28][M_AXIS_OARG_28_DMWIDTH/8-1:0];
            assign m_axis_oarg_28_tstrb = dm_tstrb[28][M_AXIS_OARG_28_DMWIDTH/8-1:0];
            assign m_axis_oarg_28_tdata = dm_tdata[28][M_AXIS_OARG_28_DMWIDTH-1:0];
            assign ap_axis_oarg_28_tready = ap_tready[28];
            assign ap_tlast[28] = ap_axis_oarg_28_tlast;
            assign ap_tvalid[28] = ap_axis_oarg_28_tvalid;
            assign ap_tdata[28][M_AXIS_OARG_28_WIDTH-1:0] = ap_axis_oarg_28_tdata;
            assign ap_tkeep[28] = {M_AXIS_OARG_28_WIDTH/8{1'b1}};
            assign ap_tstrb[28] = {M_AXIS_OARG_28_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 29) begin
            assign axis_clk[29] = m_axis_oarg_29_aclk;
            assign axis_rst[29] = m_axis_oarg_29_aresetn;
            assign dm_tready[29] = m_axis_oarg_29_tready;
            assign m_axis_oarg_29_tlast = dm_tlast[29];
            assign m_axis_oarg_29_tvalid = dm_tvalid[29];
            assign m_axis_oarg_29_tkeep = dm_tkeep[29][M_AXIS_OARG_29_DMWIDTH/8-1:0];
            assign m_axis_oarg_29_tstrb = dm_tstrb[29][M_AXIS_OARG_29_DMWIDTH/8-1:0];
            assign m_axis_oarg_29_tdata = dm_tdata[29][M_AXIS_OARG_29_DMWIDTH-1:0];
            assign ap_axis_oarg_29_tready = ap_tready[29];
            assign ap_tlast[29] = ap_axis_oarg_29_tlast;
            assign ap_tvalid[29] = ap_axis_oarg_29_tvalid;
            assign ap_tdata[29][M_AXIS_OARG_29_WIDTH-1:0] = ap_axis_oarg_29_tdata;
            assign ap_tkeep[29] = {M_AXIS_OARG_29_WIDTH/8{1'b1}};
            assign ap_tstrb[29] = {M_AXIS_OARG_29_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 30) begin
            assign axis_clk[30] = m_axis_oarg_30_aclk;
            assign axis_rst[30] = m_axis_oarg_30_aresetn;
            assign dm_tready[30] = m_axis_oarg_30_tready;
            assign m_axis_oarg_30_tlast = dm_tlast[30];
            assign m_axis_oarg_30_tvalid = dm_tvalid[30];
            assign m_axis_oarg_30_tkeep = dm_tkeep[30][M_AXIS_OARG_30_DMWIDTH/8-1:0];
            assign m_axis_oarg_30_tstrb = dm_tstrb[30][M_AXIS_OARG_30_DMWIDTH/8-1:0];
            assign m_axis_oarg_30_tdata = dm_tdata[30][M_AXIS_OARG_30_DMWIDTH-1:0];
            assign ap_axis_oarg_30_tready = ap_tready[30];
            assign ap_tlast[30] = ap_axis_oarg_30_tlast;
            assign ap_tvalid[30] = ap_axis_oarg_30_tvalid;
            assign ap_tdata[30][M_AXIS_OARG_30_WIDTH-1:0] = ap_axis_oarg_30_tdata;
            assign ap_tkeep[30] = {M_AXIS_OARG_30_WIDTH/8{1'b1}};
            assign ap_tstrb[30] = {M_AXIS_OARG_30_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 31) begin
            assign axis_clk[31] = m_axis_oarg_31_aclk;
            assign axis_rst[31] = m_axis_oarg_31_aresetn;
            assign dm_tready[31] = m_axis_oarg_31_tready;
            assign m_axis_oarg_31_tlast = dm_tlast[31];
            assign m_axis_oarg_31_tvalid = dm_tvalid[31];
            assign m_axis_oarg_31_tkeep = dm_tkeep[31][M_AXIS_OARG_31_DMWIDTH/8-1:0];
            assign m_axis_oarg_31_tstrb = dm_tstrb[31][M_AXIS_OARG_31_DMWIDTH/8-1:0];
            assign m_axis_oarg_31_tdata = dm_tdata[31][M_AXIS_OARG_31_DMWIDTH-1:0];
            assign ap_axis_oarg_31_tready = ap_tready[31];
            assign ap_tlast[31] = ap_axis_oarg_31_tlast;
            assign ap_tvalid[31] = ap_axis_oarg_31_tvalid;
            assign ap_tdata[31][M_AXIS_OARG_31_WIDTH-1:0] = ap_axis_oarg_31_tdata;
            assign ap_tkeep[31] = {M_AXIS_OARG_31_WIDTH/8{1'b1}};
            assign ap_tstrb[31] = {M_AXIS_OARG_31_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 32) begin
            assign axis_clk[32] = m_axis_oarg_32_aclk;
            assign axis_rst[32] = m_axis_oarg_32_aresetn;
            assign dm_tready[32] = m_axis_oarg_32_tready;
            assign m_axis_oarg_32_tlast = dm_tlast[32];
            assign m_axis_oarg_32_tvalid = dm_tvalid[32];
            assign m_axis_oarg_32_tkeep = dm_tkeep[32][M_AXIS_OARG_32_DMWIDTH/8-1:0];
            assign m_axis_oarg_32_tstrb = dm_tstrb[32][M_AXIS_OARG_32_DMWIDTH/8-1:0];
            assign m_axis_oarg_32_tdata = dm_tdata[32][M_AXIS_OARG_32_DMWIDTH-1:0];
            assign ap_axis_oarg_32_tready = ap_tready[32];
            assign ap_tlast[32] = ap_axis_oarg_32_tlast;
            assign ap_tvalid[32] = ap_axis_oarg_32_tvalid;
            assign ap_tdata[32][M_AXIS_OARG_32_WIDTH-1:0] = ap_axis_oarg_32_tdata;
            assign ap_tkeep[32] = {M_AXIS_OARG_32_WIDTH/8{1'b1}};
            assign ap_tstrb[32] = {M_AXIS_OARG_32_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 33) begin
            assign axis_clk[33] = m_axis_oarg_33_aclk;
            assign axis_rst[33] = m_axis_oarg_33_aresetn;
            assign dm_tready[33] = m_axis_oarg_33_tready;
            assign m_axis_oarg_33_tlast = dm_tlast[33];
            assign m_axis_oarg_33_tvalid = dm_tvalid[33];
            assign m_axis_oarg_33_tkeep = dm_tkeep[33][M_AXIS_OARG_33_DMWIDTH/8-1:0];
            assign m_axis_oarg_33_tstrb = dm_tstrb[33][M_AXIS_OARG_33_DMWIDTH/8-1:0];
            assign m_axis_oarg_33_tdata = dm_tdata[33][M_AXIS_OARG_33_DMWIDTH-1:0];
            assign ap_axis_oarg_33_tready = ap_tready[33];
            assign ap_tlast[33] = ap_axis_oarg_33_tlast;
            assign ap_tvalid[33] = ap_axis_oarg_33_tvalid;
            assign ap_tdata[33][M_AXIS_OARG_33_WIDTH-1:0] = ap_axis_oarg_33_tdata;
            assign ap_tkeep[33] = {M_AXIS_OARG_33_WIDTH/8{1'b1}};
            assign ap_tstrb[33] = {M_AXIS_OARG_33_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 34) begin
            assign axis_clk[34] = m_axis_oarg_34_aclk;
            assign axis_rst[34] = m_axis_oarg_34_aresetn;
            assign dm_tready[34] = m_axis_oarg_34_tready;
            assign m_axis_oarg_34_tlast = dm_tlast[34];
            assign m_axis_oarg_34_tvalid = dm_tvalid[34];
            assign m_axis_oarg_34_tkeep = dm_tkeep[34][M_AXIS_OARG_34_DMWIDTH/8-1:0];
            assign m_axis_oarg_34_tstrb = dm_tstrb[34][M_AXIS_OARG_34_DMWIDTH/8-1:0];
            assign m_axis_oarg_34_tdata = dm_tdata[34][M_AXIS_OARG_34_DMWIDTH-1:0];
            assign ap_axis_oarg_34_tready = ap_tready[34];
            assign ap_tlast[34] = ap_axis_oarg_34_tlast;
            assign ap_tvalid[34] = ap_axis_oarg_34_tvalid;
            assign ap_tdata[34][M_AXIS_OARG_34_WIDTH-1:0] = ap_axis_oarg_34_tdata;
            assign ap_tkeep[34] = {M_AXIS_OARG_34_WIDTH/8{1'b1}};
            assign ap_tstrb[34] = {M_AXIS_OARG_34_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 35) begin
            assign axis_clk[35] = m_axis_oarg_35_aclk;
            assign axis_rst[35] = m_axis_oarg_35_aresetn;
            assign dm_tready[35] = m_axis_oarg_35_tready;
            assign m_axis_oarg_35_tlast = dm_tlast[35];
            assign m_axis_oarg_35_tvalid = dm_tvalid[35];
            assign m_axis_oarg_35_tkeep = dm_tkeep[35][M_AXIS_OARG_35_DMWIDTH/8-1:0];
            assign m_axis_oarg_35_tstrb = dm_tstrb[35][M_AXIS_OARG_35_DMWIDTH/8-1:0];
            assign m_axis_oarg_35_tdata = dm_tdata[35][M_AXIS_OARG_35_DMWIDTH-1:0];
            assign ap_axis_oarg_35_tready = ap_tready[35];
            assign ap_tlast[35] = ap_axis_oarg_35_tlast;
            assign ap_tvalid[35] = ap_axis_oarg_35_tvalid;
            assign ap_tdata[35][M_AXIS_OARG_35_WIDTH-1:0] = ap_axis_oarg_35_tdata;
            assign ap_tkeep[35] = {M_AXIS_OARG_35_WIDTH/8{1'b1}};
            assign ap_tstrb[35] = {M_AXIS_OARG_35_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 36) begin
            assign axis_clk[36] = m_axis_oarg_36_aclk;
            assign axis_rst[36] = m_axis_oarg_36_aresetn;
            assign dm_tready[36] = m_axis_oarg_36_tready;
            assign m_axis_oarg_36_tlast = dm_tlast[36];
            assign m_axis_oarg_36_tvalid = dm_tvalid[36];
            assign m_axis_oarg_36_tkeep = dm_tkeep[36][M_AXIS_OARG_36_DMWIDTH/8-1:0];
            assign m_axis_oarg_36_tstrb = dm_tstrb[36][M_AXIS_OARG_36_DMWIDTH/8-1:0];
            assign m_axis_oarg_36_tdata = dm_tdata[36][M_AXIS_OARG_36_DMWIDTH-1:0];
            assign ap_axis_oarg_36_tready = ap_tready[36];
            assign ap_tlast[36] = ap_axis_oarg_36_tlast;
            assign ap_tvalid[36] = ap_axis_oarg_36_tvalid;
            assign ap_tdata[36][M_AXIS_OARG_36_WIDTH-1:0] = ap_axis_oarg_36_tdata;
            assign ap_tkeep[36] = {M_AXIS_OARG_36_WIDTH/8{1'b1}};
            assign ap_tstrb[36] = {M_AXIS_OARG_36_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 37) begin
            assign axis_clk[37] = m_axis_oarg_37_aclk;
            assign axis_rst[37] = m_axis_oarg_37_aresetn;
            assign dm_tready[37] = m_axis_oarg_37_tready;
            assign m_axis_oarg_37_tlast = dm_tlast[37];
            assign m_axis_oarg_37_tvalid = dm_tvalid[37];
            assign m_axis_oarg_37_tkeep = dm_tkeep[37][M_AXIS_OARG_37_DMWIDTH/8-1:0];
            assign m_axis_oarg_37_tstrb = dm_tstrb[37][M_AXIS_OARG_37_DMWIDTH/8-1:0];
            assign m_axis_oarg_37_tdata = dm_tdata[37][M_AXIS_OARG_37_DMWIDTH-1:0];
            assign ap_axis_oarg_37_tready = ap_tready[37];
            assign ap_tlast[37] = ap_axis_oarg_37_tlast;
            assign ap_tvalid[37] = ap_axis_oarg_37_tvalid;
            assign ap_tdata[37][M_AXIS_OARG_37_WIDTH-1:0] = ap_axis_oarg_37_tdata;
            assign ap_tkeep[37] = {M_AXIS_OARG_37_WIDTH/8{1'b1}};
            assign ap_tstrb[37] = {M_AXIS_OARG_37_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 38) begin
            assign axis_clk[38] = m_axis_oarg_38_aclk;
            assign axis_rst[38] = m_axis_oarg_38_aresetn;
            assign dm_tready[38] = m_axis_oarg_38_tready;
            assign m_axis_oarg_38_tlast = dm_tlast[38];
            assign m_axis_oarg_38_tvalid = dm_tvalid[38];
            assign m_axis_oarg_38_tkeep = dm_tkeep[38][M_AXIS_OARG_38_DMWIDTH/8-1:0];
            assign m_axis_oarg_38_tstrb = dm_tstrb[38][M_AXIS_OARG_38_DMWIDTH/8-1:0];
            assign m_axis_oarg_38_tdata = dm_tdata[38][M_AXIS_OARG_38_DMWIDTH-1:0];
            assign ap_axis_oarg_38_tready = ap_tready[38];
            assign ap_tlast[38] = ap_axis_oarg_38_tlast;
            assign ap_tvalid[38] = ap_axis_oarg_38_tvalid;
            assign ap_tdata[38][M_AXIS_OARG_38_WIDTH-1:0] = ap_axis_oarg_38_tdata;
            assign ap_tkeep[38] = {M_AXIS_OARG_38_WIDTH/8{1'b1}};
            assign ap_tstrb[38] = {M_AXIS_OARG_38_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 39) begin
            assign axis_clk[39] = m_axis_oarg_39_aclk;
            assign axis_rst[39] = m_axis_oarg_39_aresetn;
            assign dm_tready[39] = m_axis_oarg_39_tready;
            assign m_axis_oarg_39_tlast = dm_tlast[39];
            assign m_axis_oarg_39_tvalid = dm_tvalid[39];
            assign m_axis_oarg_39_tkeep = dm_tkeep[39][M_AXIS_OARG_39_DMWIDTH/8-1:0];
            assign m_axis_oarg_39_tstrb = dm_tstrb[39][M_AXIS_OARG_39_DMWIDTH/8-1:0];
            assign m_axis_oarg_39_tdata = dm_tdata[39][M_AXIS_OARG_39_DMWIDTH-1:0];
            assign ap_axis_oarg_39_tready = ap_tready[39];
            assign ap_tlast[39] = ap_axis_oarg_39_tlast;
            assign ap_tvalid[39] = ap_axis_oarg_39_tvalid;
            assign ap_tdata[39][M_AXIS_OARG_39_WIDTH-1:0] = ap_axis_oarg_39_tdata;
            assign ap_tkeep[39] = {M_AXIS_OARG_39_WIDTH/8{1'b1}};
            assign ap_tstrb[39] = {M_AXIS_OARG_39_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 40) begin
            assign axis_clk[40] = m_axis_oarg_40_aclk;
            assign axis_rst[40] = m_axis_oarg_40_aresetn;
            assign dm_tready[40] = m_axis_oarg_40_tready;
            assign m_axis_oarg_40_tlast = dm_tlast[40];
            assign m_axis_oarg_40_tvalid = dm_tvalid[40];
            assign m_axis_oarg_40_tkeep = dm_tkeep[40][M_AXIS_OARG_40_DMWIDTH/8-1:0];
            assign m_axis_oarg_40_tstrb = dm_tstrb[40][M_AXIS_OARG_40_DMWIDTH/8-1:0];
            assign m_axis_oarg_40_tdata = dm_tdata[40][M_AXIS_OARG_40_DMWIDTH-1:0];
            assign ap_axis_oarg_40_tready = ap_tready[40];
            assign ap_tlast[40] = ap_axis_oarg_40_tlast;
            assign ap_tvalid[40] = ap_axis_oarg_40_tvalid;
            assign ap_tdata[40][M_AXIS_OARG_40_WIDTH-1:0] = ap_axis_oarg_40_tdata;
            assign ap_tkeep[40] = {M_AXIS_OARG_40_WIDTH/8{1'b1}};
            assign ap_tstrb[40] = {M_AXIS_OARG_40_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 41) begin
            assign axis_clk[41] = m_axis_oarg_41_aclk;
            assign axis_rst[41] = m_axis_oarg_41_aresetn;
            assign dm_tready[41] = m_axis_oarg_41_tready;
            assign m_axis_oarg_41_tlast = dm_tlast[41];
            assign m_axis_oarg_41_tvalid = dm_tvalid[41];
            assign m_axis_oarg_41_tkeep = dm_tkeep[41][M_AXIS_OARG_41_DMWIDTH/8-1:0];
            assign m_axis_oarg_41_tstrb = dm_tstrb[41][M_AXIS_OARG_41_DMWIDTH/8-1:0];
            assign m_axis_oarg_41_tdata = dm_tdata[41][M_AXIS_OARG_41_DMWIDTH-1:0];
            assign ap_axis_oarg_41_tready = ap_tready[41];
            assign ap_tlast[41] = ap_axis_oarg_41_tlast;
            assign ap_tvalid[41] = ap_axis_oarg_41_tvalid;
            assign ap_tdata[41][M_AXIS_OARG_41_WIDTH-1:0] = ap_axis_oarg_41_tdata;
            assign ap_tkeep[41] = {M_AXIS_OARG_41_WIDTH/8{1'b1}};
            assign ap_tstrb[41] = {M_AXIS_OARG_41_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 42) begin
            assign axis_clk[42] = m_axis_oarg_42_aclk;
            assign axis_rst[42] = m_axis_oarg_42_aresetn;
            assign dm_tready[42] = m_axis_oarg_42_tready;
            assign m_axis_oarg_42_tlast = dm_tlast[42];
            assign m_axis_oarg_42_tvalid = dm_tvalid[42];
            assign m_axis_oarg_42_tkeep = dm_tkeep[42][M_AXIS_OARG_42_DMWIDTH/8-1:0];
            assign m_axis_oarg_42_tstrb = dm_tstrb[42][M_AXIS_OARG_42_DMWIDTH/8-1:0];
            assign m_axis_oarg_42_tdata = dm_tdata[42][M_AXIS_OARG_42_DMWIDTH-1:0];
            assign ap_axis_oarg_42_tready = ap_tready[42];
            assign ap_tlast[42] = ap_axis_oarg_42_tlast;
            assign ap_tvalid[42] = ap_axis_oarg_42_tvalid;
            assign ap_tdata[42][M_AXIS_OARG_42_WIDTH-1:0] = ap_axis_oarg_42_tdata;
            assign ap_tkeep[42] = {M_AXIS_OARG_42_WIDTH/8{1'b1}};
            assign ap_tstrb[42] = {M_AXIS_OARG_42_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 43) begin
            assign axis_clk[43] = m_axis_oarg_43_aclk;
            assign axis_rst[43] = m_axis_oarg_43_aresetn;
            assign dm_tready[43] = m_axis_oarg_43_tready;
            assign m_axis_oarg_43_tlast = dm_tlast[43];
            assign m_axis_oarg_43_tvalid = dm_tvalid[43];
            assign m_axis_oarg_43_tkeep = dm_tkeep[43][M_AXIS_OARG_43_DMWIDTH/8-1:0];
            assign m_axis_oarg_43_tstrb = dm_tstrb[43][M_AXIS_OARG_43_DMWIDTH/8-1:0];
            assign m_axis_oarg_43_tdata = dm_tdata[43][M_AXIS_OARG_43_DMWIDTH-1:0];
            assign ap_axis_oarg_43_tready = ap_tready[43];
            assign ap_tlast[43] = ap_axis_oarg_43_tlast;
            assign ap_tvalid[43] = ap_axis_oarg_43_tvalid;
            assign ap_tdata[43][M_AXIS_OARG_43_WIDTH-1:0] = ap_axis_oarg_43_tdata;
            assign ap_tkeep[43] = {M_AXIS_OARG_43_WIDTH/8{1'b1}};
            assign ap_tstrb[43] = {M_AXIS_OARG_43_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 44) begin
            assign axis_clk[44] = m_axis_oarg_44_aclk;
            assign axis_rst[44] = m_axis_oarg_44_aresetn;
            assign dm_tready[44] = m_axis_oarg_44_tready;
            assign m_axis_oarg_44_tlast = dm_tlast[44];
            assign m_axis_oarg_44_tvalid = dm_tvalid[44];
            assign m_axis_oarg_44_tkeep = dm_tkeep[44][M_AXIS_OARG_44_DMWIDTH/8-1:0];
            assign m_axis_oarg_44_tstrb = dm_tstrb[44][M_AXIS_OARG_44_DMWIDTH/8-1:0];
            assign m_axis_oarg_44_tdata = dm_tdata[44][M_AXIS_OARG_44_DMWIDTH-1:0];
            assign ap_axis_oarg_44_tready = ap_tready[44];
            assign ap_tlast[44] = ap_axis_oarg_44_tlast;
            assign ap_tvalid[44] = ap_axis_oarg_44_tvalid;
            assign ap_tdata[44][M_AXIS_OARG_44_WIDTH-1:0] = ap_axis_oarg_44_tdata;
            assign ap_tkeep[44] = {M_AXIS_OARG_44_WIDTH/8{1'b1}};
            assign ap_tstrb[44] = {M_AXIS_OARG_44_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 45) begin
            assign axis_clk[45] = m_axis_oarg_45_aclk;
            assign axis_rst[45] = m_axis_oarg_45_aresetn;
            assign dm_tready[45] = m_axis_oarg_45_tready;
            assign m_axis_oarg_45_tlast = dm_tlast[45];
            assign m_axis_oarg_45_tvalid = dm_tvalid[45];
            assign m_axis_oarg_45_tkeep = dm_tkeep[45][M_AXIS_OARG_45_DMWIDTH/8-1:0];
            assign m_axis_oarg_45_tstrb = dm_tstrb[45][M_AXIS_OARG_45_DMWIDTH/8-1:0];
            assign m_axis_oarg_45_tdata = dm_tdata[45][M_AXIS_OARG_45_DMWIDTH-1:0];
            assign ap_axis_oarg_45_tready = ap_tready[45];
            assign ap_tlast[45] = ap_axis_oarg_45_tlast;
            assign ap_tvalid[45] = ap_axis_oarg_45_tvalid;
            assign ap_tdata[45][M_AXIS_OARG_45_WIDTH-1:0] = ap_axis_oarg_45_tdata;
            assign ap_tkeep[45] = {M_AXIS_OARG_45_WIDTH/8{1'b1}};
            assign ap_tstrb[45] = {M_AXIS_OARG_45_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 46) begin
            assign axis_clk[46] = m_axis_oarg_46_aclk;
            assign axis_rst[46] = m_axis_oarg_46_aresetn;
            assign dm_tready[46] = m_axis_oarg_46_tready;
            assign m_axis_oarg_46_tlast = dm_tlast[46];
            assign m_axis_oarg_46_tvalid = dm_tvalid[46];
            assign m_axis_oarg_46_tkeep = dm_tkeep[46][M_AXIS_OARG_46_DMWIDTH/8-1:0];
            assign m_axis_oarg_46_tstrb = dm_tstrb[46][M_AXIS_OARG_46_DMWIDTH/8-1:0];
            assign m_axis_oarg_46_tdata = dm_tdata[46][M_AXIS_OARG_46_DMWIDTH-1:0];
            assign ap_axis_oarg_46_tready = ap_tready[46];
            assign ap_tlast[46] = ap_axis_oarg_46_tlast;
            assign ap_tvalid[46] = ap_axis_oarg_46_tvalid;
            assign ap_tdata[46][M_AXIS_OARG_46_WIDTH-1:0] = ap_axis_oarg_46_tdata;
            assign ap_tkeep[46] = {M_AXIS_OARG_46_WIDTH/8{1'b1}};
            assign ap_tstrb[46] = {M_AXIS_OARG_46_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 47) begin
            assign axis_clk[47] = m_axis_oarg_47_aclk;
            assign axis_rst[47] = m_axis_oarg_47_aresetn;
            assign dm_tready[47] = m_axis_oarg_47_tready;
            assign m_axis_oarg_47_tlast = dm_tlast[47];
            assign m_axis_oarg_47_tvalid = dm_tvalid[47];
            assign m_axis_oarg_47_tkeep = dm_tkeep[47][M_AXIS_OARG_47_DMWIDTH/8-1:0];
            assign m_axis_oarg_47_tstrb = dm_tstrb[47][M_AXIS_OARG_47_DMWIDTH/8-1:0];
            assign m_axis_oarg_47_tdata = dm_tdata[47][M_AXIS_OARG_47_DMWIDTH-1:0];
            assign ap_axis_oarg_47_tready = ap_tready[47];
            assign ap_tlast[47] = ap_axis_oarg_47_tlast;
            assign ap_tvalid[47] = ap_axis_oarg_47_tvalid;
            assign ap_tdata[47][M_AXIS_OARG_47_WIDTH-1:0] = ap_axis_oarg_47_tdata;
            assign ap_tkeep[47] = {M_AXIS_OARG_47_WIDTH/8{1'b1}};
            assign ap_tstrb[47] = {M_AXIS_OARG_47_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 48) begin
            assign axis_clk[48] = m_axis_oarg_48_aclk;
            assign axis_rst[48] = m_axis_oarg_48_aresetn;
            assign dm_tready[48] = m_axis_oarg_48_tready;
            assign m_axis_oarg_48_tlast = dm_tlast[48];
            assign m_axis_oarg_48_tvalid = dm_tvalid[48];
            assign m_axis_oarg_48_tkeep = dm_tkeep[48][M_AXIS_OARG_48_DMWIDTH/8-1:0];
            assign m_axis_oarg_48_tstrb = dm_tstrb[48][M_AXIS_OARG_48_DMWIDTH/8-1:0];
            assign m_axis_oarg_48_tdata = dm_tdata[48][M_AXIS_OARG_48_DMWIDTH-1:0];
            assign ap_axis_oarg_48_tready = ap_tready[48];
            assign ap_tlast[48] = ap_axis_oarg_48_tlast;
            assign ap_tvalid[48] = ap_axis_oarg_48_tvalid;
            assign ap_tdata[48][M_AXIS_OARG_48_WIDTH-1:0] = ap_axis_oarg_48_tdata;
            assign ap_tkeep[48] = {M_AXIS_OARG_48_WIDTH/8{1'b1}};
            assign ap_tstrb[48] = {M_AXIS_OARG_48_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 49) begin
            assign axis_clk[49] = m_axis_oarg_49_aclk;
            assign axis_rst[49] = m_axis_oarg_49_aresetn;
            assign dm_tready[49] = m_axis_oarg_49_tready;
            assign m_axis_oarg_49_tlast = dm_tlast[49];
            assign m_axis_oarg_49_tvalid = dm_tvalid[49];
            assign m_axis_oarg_49_tkeep = dm_tkeep[49][M_AXIS_OARG_49_DMWIDTH/8-1:0];
            assign m_axis_oarg_49_tstrb = dm_tstrb[49][M_AXIS_OARG_49_DMWIDTH/8-1:0];
            assign m_axis_oarg_49_tdata = dm_tdata[49][M_AXIS_OARG_49_DMWIDTH-1:0];
            assign ap_axis_oarg_49_tready = ap_tready[49];
            assign ap_tlast[49] = ap_axis_oarg_49_tlast;
            assign ap_tvalid[49] = ap_axis_oarg_49_tvalid;
            assign ap_tdata[49][M_AXIS_OARG_49_WIDTH-1:0] = ap_axis_oarg_49_tdata;
            assign ap_tkeep[49] = {M_AXIS_OARG_49_WIDTH/8{1'b1}};
            assign ap_tstrb[49] = {M_AXIS_OARG_49_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 50) begin
            assign axis_clk[50] = m_axis_oarg_50_aclk;
            assign axis_rst[50] = m_axis_oarg_50_aresetn;
            assign dm_tready[50] = m_axis_oarg_50_tready;
            assign m_axis_oarg_50_tlast = dm_tlast[50];
            assign m_axis_oarg_50_tvalid = dm_tvalid[50];
            assign m_axis_oarg_50_tkeep = dm_tkeep[50][M_AXIS_OARG_50_DMWIDTH/8-1:0];
            assign m_axis_oarg_50_tstrb = dm_tstrb[50][M_AXIS_OARG_50_DMWIDTH/8-1:0];
            assign m_axis_oarg_50_tdata = dm_tdata[50][M_AXIS_OARG_50_DMWIDTH-1:0];
            assign ap_axis_oarg_50_tready = ap_tready[50];
            assign ap_tlast[50] = ap_axis_oarg_50_tlast;
            assign ap_tvalid[50] = ap_axis_oarg_50_tvalid;
            assign ap_tdata[50][M_AXIS_OARG_50_WIDTH-1:0] = ap_axis_oarg_50_tdata;
            assign ap_tkeep[50] = {M_AXIS_OARG_50_WIDTH/8{1'b1}};
            assign ap_tstrb[50] = {M_AXIS_OARG_50_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 51) begin
            assign axis_clk[51] = m_axis_oarg_51_aclk;
            assign axis_rst[51] = m_axis_oarg_51_aresetn;
            assign dm_tready[51] = m_axis_oarg_51_tready;
            assign m_axis_oarg_51_tlast = dm_tlast[51];
            assign m_axis_oarg_51_tvalid = dm_tvalid[51];
            assign m_axis_oarg_51_tkeep = dm_tkeep[51][M_AXIS_OARG_51_DMWIDTH/8-1:0];
            assign m_axis_oarg_51_tstrb = dm_tstrb[51][M_AXIS_OARG_51_DMWIDTH/8-1:0];
            assign m_axis_oarg_51_tdata = dm_tdata[51][M_AXIS_OARG_51_DMWIDTH-1:0];
            assign ap_axis_oarg_51_tready = ap_tready[51];
            assign ap_tlast[51] = ap_axis_oarg_51_tlast;
            assign ap_tvalid[51] = ap_axis_oarg_51_tvalid;
            assign ap_tdata[51][M_AXIS_OARG_51_WIDTH-1:0] = ap_axis_oarg_51_tdata;
            assign ap_tkeep[51] = {M_AXIS_OARG_51_WIDTH/8{1'b1}};
            assign ap_tstrb[51] = {M_AXIS_OARG_51_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 52) begin
            assign axis_clk[52] = m_axis_oarg_52_aclk;
            assign axis_rst[52] = m_axis_oarg_52_aresetn;
            assign dm_tready[52] = m_axis_oarg_52_tready;
            assign m_axis_oarg_52_tlast = dm_tlast[52];
            assign m_axis_oarg_52_tvalid = dm_tvalid[52];
            assign m_axis_oarg_52_tkeep = dm_tkeep[52][M_AXIS_OARG_52_DMWIDTH/8-1:0];
            assign m_axis_oarg_52_tstrb = dm_tstrb[52][M_AXIS_OARG_52_DMWIDTH/8-1:0];
            assign m_axis_oarg_52_tdata = dm_tdata[52][M_AXIS_OARG_52_DMWIDTH-1:0];
            assign ap_axis_oarg_52_tready = ap_tready[52];
            assign ap_tlast[52] = ap_axis_oarg_52_tlast;
            assign ap_tvalid[52] = ap_axis_oarg_52_tvalid;
            assign ap_tdata[52][M_AXIS_OARG_52_WIDTH-1:0] = ap_axis_oarg_52_tdata;
            assign ap_tkeep[52] = {M_AXIS_OARG_52_WIDTH/8{1'b1}};
            assign ap_tstrb[52] = {M_AXIS_OARG_52_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 53) begin
            assign axis_clk[53] = m_axis_oarg_53_aclk;
            assign axis_rst[53] = m_axis_oarg_53_aresetn;
            assign dm_tready[53] = m_axis_oarg_53_tready;
            assign m_axis_oarg_53_tlast = dm_tlast[53];
            assign m_axis_oarg_53_tvalid = dm_tvalid[53];
            assign m_axis_oarg_53_tkeep = dm_tkeep[53][M_AXIS_OARG_53_DMWIDTH/8-1:0];
            assign m_axis_oarg_53_tstrb = dm_tstrb[53][M_AXIS_OARG_53_DMWIDTH/8-1:0];
            assign m_axis_oarg_53_tdata = dm_tdata[53][M_AXIS_OARG_53_DMWIDTH-1:0];
            assign ap_axis_oarg_53_tready = ap_tready[53];
            assign ap_tlast[53] = ap_axis_oarg_53_tlast;
            assign ap_tvalid[53] = ap_axis_oarg_53_tvalid;
            assign ap_tdata[53][M_AXIS_OARG_53_WIDTH-1:0] = ap_axis_oarg_53_tdata;
            assign ap_tkeep[53] = {M_AXIS_OARG_53_WIDTH/8{1'b1}};
            assign ap_tstrb[53] = {M_AXIS_OARG_53_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 54) begin
            assign axis_clk[54] = m_axis_oarg_54_aclk;
            assign axis_rst[54] = m_axis_oarg_54_aresetn;
            assign dm_tready[54] = m_axis_oarg_54_tready;
            assign m_axis_oarg_54_tlast = dm_tlast[54];
            assign m_axis_oarg_54_tvalid = dm_tvalid[54];
            assign m_axis_oarg_54_tkeep = dm_tkeep[54][M_AXIS_OARG_54_DMWIDTH/8-1:0];
            assign m_axis_oarg_54_tstrb = dm_tstrb[54][M_AXIS_OARG_54_DMWIDTH/8-1:0];
            assign m_axis_oarg_54_tdata = dm_tdata[54][M_AXIS_OARG_54_DMWIDTH-1:0];
            assign ap_axis_oarg_54_tready = ap_tready[54];
            assign ap_tlast[54] = ap_axis_oarg_54_tlast;
            assign ap_tvalid[54] = ap_axis_oarg_54_tvalid;
            assign ap_tdata[54][M_AXIS_OARG_54_WIDTH-1:0] = ap_axis_oarg_54_tdata;
            assign ap_tkeep[54] = {M_AXIS_OARG_54_WIDTH/8{1'b1}};
            assign ap_tstrb[54] = {M_AXIS_OARG_54_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 55) begin
            assign axis_clk[55] = m_axis_oarg_55_aclk;
            assign axis_rst[55] = m_axis_oarg_55_aresetn;
            assign dm_tready[55] = m_axis_oarg_55_tready;
            assign m_axis_oarg_55_tlast = dm_tlast[55];
            assign m_axis_oarg_55_tvalid = dm_tvalid[55];
            assign m_axis_oarg_55_tkeep = dm_tkeep[55][M_AXIS_OARG_55_DMWIDTH/8-1:0];
            assign m_axis_oarg_55_tstrb = dm_tstrb[55][M_AXIS_OARG_55_DMWIDTH/8-1:0];
            assign m_axis_oarg_55_tdata = dm_tdata[55][M_AXIS_OARG_55_DMWIDTH-1:0];
            assign ap_axis_oarg_55_tready = ap_tready[55];
            assign ap_tlast[55] = ap_axis_oarg_55_tlast;
            assign ap_tvalid[55] = ap_axis_oarg_55_tvalid;
            assign ap_tdata[55][M_AXIS_OARG_55_WIDTH-1:0] = ap_axis_oarg_55_tdata;
            assign ap_tkeep[55] = {M_AXIS_OARG_55_WIDTH/8{1'b1}};
            assign ap_tstrb[55] = {M_AXIS_OARG_55_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 56) begin
            assign axis_clk[56] = m_axis_oarg_56_aclk;
            assign axis_rst[56] = m_axis_oarg_56_aresetn;
            assign dm_tready[56] = m_axis_oarg_56_tready;
            assign m_axis_oarg_56_tlast = dm_tlast[56];
            assign m_axis_oarg_56_tvalid = dm_tvalid[56];
            assign m_axis_oarg_56_tkeep = dm_tkeep[56][M_AXIS_OARG_56_DMWIDTH/8-1:0];
            assign m_axis_oarg_56_tstrb = dm_tstrb[56][M_AXIS_OARG_56_DMWIDTH/8-1:0];
            assign m_axis_oarg_56_tdata = dm_tdata[56][M_AXIS_OARG_56_DMWIDTH-1:0];
            assign ap_axis_oarg_56_tready = ap_tready[56];
            assign ap_tlast[56] = ap_axis_oarg_56_tlast;
            assign ap_tvalid[56] = ap_axis_oarg_56_tvalid;
            assign ap_tdata[56][M_AXIS_OARG_56_WIDTH-1:0] = ap_axis_oarg_56_tdata;
            assign ap_tkeep[56] = {M_AXIS_OARG_56_WIDTH/8{1'b1}};
            assign ap_tstrb[56] = {M_AXIS_OARG_56_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 57) begin
            assign axis_clk[57] = m_axis_oarg_57_aclk;
            assign axis_rst[57] = m_axis_oarg_57_aresetn;
            assign dm_tready[57] = m_axis_oarg_57_tready;
            assign m_axis_oarg_57_tlast = dm_tlast[57];
            assign m_axis_oarg_57_tvalid = dm_tvalid[57];
            assign m_axis_oarg_57_tkeep = dm_tkeep[57][M_AXIS_OARG_57_DMWIDTH/8-1:0];
            assign m_axis_oarg_57_tstrb = dm_tstrb[57][M_AXIS_OARG_57_DMWIDTH/8-1:0];
            assign m_axis_oarg_57_tdata = dm_tdata[57][M_AXIS_OARG_57_DMWIDTH-1:0];
            assign ap_axis_oarg_57_tready = ap_tready[57];
            assign ap_tlast[57] = ap_axis_oarg_57_tlast;
            assign ap_tvalid[57] = ap_axis_oarg_57_tvalid;
            assign ap_tdata[57][M_AXIS_OARG_57_WIDTH-1:0] = ap_axis_oarg_57_tdata;
            assign ap_tkeep[57] = {M_AXIS_OARG_57_WIDTH/8{1'b1}};
            assign ap_tstrb[57] = {M_AXIS_OARG_57_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 58) begin
            assign axis_clk[58] = m_axis_oarg_58_aclk;
            assign axis_rst[58] = m_axis_oarg_58_aresetn;
            assign dm_tready[58] = m_axis_oarg_58_tready;
            assign m_axis_oarg_58_tlast = dm_tlast[58];
            assign m_axis_oarg_58_tvalid = dm_tvalid[58];
            assign m_axis_oarg_58_tkeep = dm_tkeep[58][M_AXIS_OARG_58_DMWIDTH/8-1:0];
            assign m_axis_oarg_58_tstrb = dm_tstrb[58][M_AXIS_OARG_58_DMWIDTH/8-1:0];
            assign m_axis_oarg_58_tdata = dm_tdata[58][M_AXIS_OARG_58_DMWIDTH-1:0];
            assign ap_axis_oarg_58_tready = ap_tready[58];
            assign ap_tlast[58] = ap_axis_oarg_58_tlast;
            assign ap_tvalid[58] = ap_axis_oarg_58_tvalid;
            assign ap_tdata[58][M_AXIS_OARG_58_WIDTH-1:0] = ap_axis_oarg_58_tdata;
            assign ap_tkeep[58] = {M_AXIS_OARG_58_WIDTH/8{1'b1}};
            assign ap_tstrb[58] = {M_AXIS_OARG_58_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 59) begin
            assign axis_clk[59] = m_axis_oarg_59_aclk;
            assign axis_rst[59] = m_axis_oarg_59_aresetn;
            assign dm_tready[59] = m_axis_oarg_59_tready;
            assign m_axis_oarg_59_tlast = dm_tlast[59];
            assign m_axis_oarg_59_tvalid = dm_tvalid[59];
            assign m_axis_oarg_59_tkeep = dm_tkeep[59][M_AXIS_OARG_59_DMWIDTH/8-1:0];
            assign m_axis_oarg_59_tstrb = dm_tstrb[59][M_AXIS_OARG_59_DMWIDTH/8-1:0];
            assign m_axis_oarg_59_tdata = dm_tdata[59][M_AXIS_OARG_59_DMWIDTH-1:0];
            assign ap_axis_oarg_59_tready = ap_tready[59];
            assign ap_tlast[59] = ap_axis_oarg_59_tlast;
            assign ap_tvalid[59] = ap_axis_oarg_59_tvalid;
            assign ap_tdata[59][M_AXIS_OARG_59_WIDTH-1:0] = ap_axis_oarg_59_tdata;
            assign ap_tkeep[59] = {M_AXIS_OARG_59_WIDTH/8{1'b1}};
            assign ap_tstrb[59] = {M_AXIS_OARG_59_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 60) begin
            assign axis_clk[60] = m_axis_oarg_60_aclk;
            assign axis_rst[60] = m_axis_oarg_60_aresetn;
            assign dm_tready[60] = m_axis_oarg_60_tready;
            assign m_axis_oarg_60_tlast = dm_tlast[60];
            assign m_axis_oarg_60_tvalid = dm_tvalid[60];
            assign m_axis_oarg_60_tkeep = dm_tkeep[60][M_AXIS_OARG_60_DMWIDTH/8-1:0];
            assign m_axis_oarg_60_tstrb = dm_tstrb[60][M_AXIS_OARG_60_DMWIDTH/8-1:0];
            assign m_axis_oarg_60_tdata = dm_tdata[60][M_AXIS_OARG_60_DMWIDTH-1:0];
            assign ap_axis_oarg_60_tready = ap_tready[60];
            assign ap_tlast[60] = ap_axis_oarg_60_tlast;
            assign ap_tvalid[60] = ap_axis_oarg_60_tvalid;
            assign ap_tdata[60][M_AXIS_OARG_60_WIDTH-1:0] = ap_axis_oarg_60_tdata;
            assign ap_tkeep[60] = {M_AXIS_OARG_60_WIDTH/8{1'b1}};
            assign ap_tstrb[60] = {M_AXIS_OARG_60_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 61) begin
            assign axis_clk[61] = m_axis_oarg_61_aclk;
            assign axis_rst[61] = m_axis_oarg_61_aresetn;
            assign dm_tready[61] = m_axis_oarg_61_tready;
            assign m_axis_oarg_61_tlast = dm_tlast[61];
            assign m_axis_oarg_61_tvalid = dm_tvalid[61];
            assign m_axis_oarg_61_tkeep = dm_tkeep[61][M_AXIS_OARG_61_DMWIDTH/8-1:0];
            assign m_axis_oarg_61_tstrb = dm_tstrb[61][M_AXIS_OARG_61_DMWIDTH/8-1:0];
            assign m_axis_oarg_61_tdata = dm_tdata[61][M_AXIS_OARG_61_DMWIDTH-1:0];
            assign ap_axis_oarg_61_tready = ap_tready[61];
            assign ap_tlast[61] = ap_axis_oarg_61_tlast;
            assign ap_tvalid[61] = ap_axis_oarg_61_tvalid;
            assign ap_tdata[61][M_AXIS_OARG_61_WIDTH-1:0] = ap_axis_oarg_61_tdata;
            assign ap_tkeep[61] = {M_AXIS_OARG_61_WIDTH/8{1'b1}};
            assign ap_tstrb[61] = {M_AXIS_OARG_61_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 62) begin
            assign axis_clk[62] = m_axis_oarg_62_aclk;
            assign axis_rst[62] = m_axis_oarg_62_aresetn;
            assign dm_tready[62] = m_axis_oarg_62_tready;
            assign m_axis_oarg_62_tlast = dm_tlast[62];
            assign m_axis_oarg_62_tvalid = dm_tvalid[62];
            assign m_axis_oarg_62_tkeep = dm_tkeep[62][M_AXIS_OARG_62_DMWIDTH/8-1:0];
            assign m_axis_oarg_62_tstrb = dm_tstrb[62][M_AXIS_OARG_62_DMWIDTH/8-1:0];
            assign m_axis_oarg_62_tdata = dm_tdata[62][M_AXIS_OARG_62_DMWIDTH-1:0];
            assign ap_axis_oarg_62_tready = ap_tready[62];
            assign ap_tlast[62] = ap_axis_oarg_62_tlast;
            assign ap_tvalid[62] = ap_axis_oarg_62_tvalid;
            assign ap_tdata[62][M_AXIS_OARG_62_WIDTH-1:0] = ap_axis_oarg_62_tdata;
            assign ap_tkeep[62] = {M_AXIS_OARG_62_WIDTH/8{1'b1}};
            assign ap_tstrb[62] = {M_AXIS_OARG_62_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 63) begin
            assign axis_clk[63] = m_axis_oarg_63_aclk;
            assign axis_rst[63] = m_axis_oarg_63_aresetn;
            assign dm_tready[63] = m_axis_oarg_63_tready;
            assign m_axis_oarg_63_tlast = dm_tlast[63];
            assign m_axis_oarg_63_tvalid = dm_tvalid[63];
            assign m_axis_oarg_63_tkeep = dm_tkeep[63][M_AXIS_OARG_63_DMWIDTH/8-1:0];
            assign m_axis_oarg_63_tstrb = dm_tstrb[63][M_AXIS_OARG_63_DMWIDTH/8-1:0];
            assign m_axis_oarg_63_tdata = dm_tdata[63][M_AXIS_OARG_63_DMWIDTH-1:0];
            assign ap_axis_oarg_63_tready = ap_tready[63];
            assign ap_tlast[63] = ap_axis_oarg_63_tlast;
            assign ap_tvalid[63] = ap_axis_oarg_63_tvalid;
            assign ap_tdata[63][M_AXIS_OARG_63_WIDTH-1:0] = ap_axis_oarg_63_tdata;
            assign ap_tkeep[63] = {M_AXIS_OARG_63_WIDTH/8{1'b1}};
            assign ap_tstrb[63] = {M_AXIS_OARG_63_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 64) begin
            assign axis_clk[64] = m_axis_oarg_64_aclk;
            assign axis_rst[64] = m_axis_oarg_64_aresetn;
            assign dm_tready[64] = m_axis_oarg_64_tready;
            assign m_axis_oarg_64_tlast = dm_tlast[64];
            assign m_axis_oarg_64_tvalid = dm_tvalid[64];
            assign m_axis_oarg_64_tkeep = dm_tkeep[64][M_AXIS_OARG_64_DMWIDTH/8-1:0];
            assign m_axis_oarg_64_tstrb = dm_tstrb[64][M_AXIS_OARG_64_DMWIDTH/8-1:0];
            assign m_axis_oarg_64_tdata = dm_tdata[64][M_AXIS_OARG_64_DMWIDTH-1:0];
            assign ap_axis_oarg_64_tready = ap_tready[64];
            assign ap_tlast[64] = ap_axis_oarg_64_tlast;
            assign ap_tvalid[64] = ap_axis_oarg_64_tvalid;
            assign ap_tdata[64][M_AXIS_OARG_64_WIDTH-1:0] = ap_axis_oarg_64_tdata;
            assign ap_tkeep[64] = {M_AXIS_OARG_64_WIDTH/8{1'b1}};
            assign ap_tstrb[64] = {M_AXIS_OARG_64_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 65) begin
            assign axis_clk[65] = m_axis_oarg_65_aclk;
            assign axis_rst[65] = m_axis_oarg_65_aresetn;
            assign dm_tready[65] = m_axis_oarg_65_tready;
            assign m_axis_oarg_65_tlast = dm_tlast[65];
            assign m_axis_oarg_65_tvalid = dm_tvalid[65];
            assign m_axis_oarg_65_tkeep = dm_tkeep[65][M_AXIS_OARG_65_DMWIDTH/8-1:0];
            assign m_axis_oarg_65_tstrb = dm_tstrb[65][M_AXIS_OARG_65_DMWIDTH/8-1:0];
            assign m_axis_oarg_65_tdata = dm_tdata[65][M_AXIS_OARG_65_DMWIDTH-1:0];
            assign ap_axis_oarg_65_tready = ap_tready[65];
            assign ap_tlast[65] = ap_axis_oarg_65_tlast;
            assign ap_tvalid[65] = ap_axis_oarg_65_tvalid;
            assign ap_tdata[65][M_AXIS_OARG_65_WIDTH-1:0] = ap_axis_oarg_65_tdata;
            assign ap_tkeep[65] = {M_AXIS_OARG_65_WIDTH/8{1'b1}};
            assign ap_tstrb[65] = {M_AXIS_OARG_65_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 66) begin
            assign axis_clk[66] = m_axis_oarg_66_aclk;
            assign axis_rst[66] = m_axis_oarg_66_aresetn;
            assign dm_tready[66] = m_axis_oarg_66_tready;
            assign m_axis_oarg_66_tlast = dm_tlast[66];
            assign m_axis_oarg_66_tvalid = dm_tvalid[66];
            assign m_axis_oarg_66_tkeep = dm_tkeep[66][M_AXIS_OARG_66_DMWIDTH/8-1:0];
            assign m_axis_oarg_66_tstrb = dm_tstrb[66][M_AXIS_OARG_66_DMWIDTH/8-1:0];
            assign m_axis_oarg_66_tdata = dm_tdata[66][M_AXIS_OARG_66_DMWIDTH-1:0];
            assign ap_axis_oarg_66_tready = ap_tready[66];
            assign ap_tlast[66] = ap_axis_oarg_66_tlast;
            assign ap_tvalid[66] = ap_axis_oarg_66_tvalid;
            assign ap_tdata[66][M_AXIS_OARG_66_WIDTH-1:0] = ap_axis_oarg_66_tdata;
            assign ap_tkeep[66] = {M_AXIS_OARG_66_WIDTH/8{1'b1}};
            assign ap_tstrb[66] = {M_AXIS_OARG_66_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 67) begin
            assign axis_clk[67] = m_axis_oarg_67_aclk;
            assign axis_rst[67] = m_axis_oarg_67_aresetn;
            assign dm_tready[67] = m_axis_oarg_67_tready;
            assign m_axis_oarg_67_tlast = dm_tlast[67];
            assign m_axis_oarg_67_tvalid = dm_tvalid[67];
            assign m_axis_oarg_67_tkeep = dm_tkeep[67][M_AXIS_OARG_67_DMWIDTH/8-1:0];
            assign m_axis_oarg_67_tstrb = dm_tstrb[67][M_AXIS_OARG_67_DMWIDTH/8-1:0];
            assign m_axis_oarg_67_tdata = dm_tdata[67][M_AXIS_OARG_67_DMWIDTH-1:0];
            assign ap_axis_oarg_67_tready = ap_tready[67];
            assign ap_tlast[67] = ap_axis_oarg_67_tlast;
            assign ap_tvalid[67] = ap_axis_oarg_67_tvalid;
            assign ap_tdata[67][M_AXIS_OARG_67_WIDTH-1:0] = ap_axis_oarg_67_tdata;
            assign ap_tkeep[67] = {M_AXIS_OARG_67_WIDTH/8{1'b1}};
            assign ap_tstrb[67] = {M_AXIS_OARG_67_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 68) begin
            assign axis_clk[68] = m_axis_oarg_68_aclk;
            assign axis_rst[68] = m_axis_oarg_68_aresetn;
            assign dm_tready[68] = m_axis_oarg_68_tready;
            assign m_axis_oarg_68_tlast = dm_tlast[68];
            assign m_axis_oarg_68_tvalid = dm_tvalid[68];
            assign m_axis_oarg_68_tkeep = dm_tkeep[68][M_AXIS_OARG_68_DMWIDTH/8-1:0];
            assign m_axis_oarg_68_tstrb = dm_tstrb[68][M_AXIS_OARG_68_DMWIDTH/8-1:0];
            assign m_axis_oarg_68_tdata = dm_tdata[68][M_AXIS_OARG_68_DMWIDTH-1:0];
            assign ap_axis_oarg_68_tready = ap_tready[68];
            assign ap_tlast[68] = ap_axis_oarg_68_tlast;
            assign ap_tvalid[68] = ap_axis_oarg_68_tvalid;
            assign ap_tdata[68][M_AXIS_OARG_68_WIDTH-1:0] = ap_axis_oarg_68_tdata;
            assign ap_tkeep[68] = {M_AXIS_OARG_68_WIDTH/8{1'b1}};
            assign ap_tstrb[68] = {M_AXIS_OARG_68_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 69) begin
            assign axis_clk[69] = m_axis_oarg_69_aclk;
            assign axis_rst[69] = m_axis_oarg_69_aresetn;
            assign dm_tready[69] = m_axis_oarg_69_tready;
            assign m_axis_oarg_69_tlast = dm_tlast[69];
            assign m_axis_oarg_69_tvalid = dm_tvalid[69];
            assign m_axis_oarg_69_tkeep = dm_tkeep[69][M_AXIS_OARG_69_DMWIDTH/8-1:0];
            assign m_axis_oarg_69_tstrb = dm_tstrb[69][M_AXIS_OARG_69_DMWIDTH/8-1:0];
            assign m_axis_oarg_69_tdata = dm_tdata[69][M_AXIS_OARG_69_DMWIDTH-1:0];
            assign ap_axis_oarg_69_tready = ap_tready[69];
            assign ap_tlast[69] = ap_axis_oarg_69_tlast;
            assign ap_tvalid[69] = ap_axis_oarg_69_tvalid;
            assign ap_tdata[69][M_AXIS_OARG_69_WIDTH-1:0] = ap_axis_oarg_69_tdata;
            assign ap_tkeep[69] = {M_AXIS_OARG_69_WIDTH/8{1'b1}};
            assign ap_tstrb[69] = {M_AXIS_OARG_69_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 70) begin
            assign axis_clk[70] = m_axis_oarg_70_aclk;
            assign axis_rst[70] = m_axis_oarg_70_aresetn;
            assign dm_tready[70] = m_axis_oarg_70_tready;
            assign m_axis_oarg_70_tlast = dm_tlast[70];
            assign m_axis_oarg_70_tvalid = dm_tvalid[70];
            assign m_axis_oarg_70_tkeep = dm_tkeep[70][M_AXIS_OARG_70_DMWIDTH/8-1:0];
            assign m_axis_oarg_70_tstrb = dm_tstrb[70][M_AXIS_OARG_70_DMWIDTH/8-1:0];
            assign m_axis_oarg_70_tdata = dm_tdata[70][M_AXIS_OARG_70_DMWIDTH-1:0];
            assign ap_axis_oarg_70_tready = ap_tready[70];
            assign ap_tlast[70] = ap_axis_oarg_70_tlast;
            assign ap_tvalid[70] = ap_axis_oarg_70_tvalid;
            assign ap_tdata[70][M_AXIS_OARG_70_WIDTH-1:0] = ap_axis_oarg_70_tdata;
            assign ap_tkeep[70] = {M_AXIS_OARG_70_WIDTH/8{1'b1}};
            assign ap_tstrb[70] = {M_AXIS_OARG_70_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 71) begin
            assign axis_clk[71] = m_axis_oarg_71_aclk;
            assign axis_rst[71] = m_axis_oarg_71_aresetn;
            assign dm_tready[71] = m_axis_oarg_71_tready;
            assign m_axis_oarg_71_tlast = dm_tlast[71];
            assign m_axis_oarg_71_tvalid = dm_tvalid[71];
            assign m_axis_oarg_71_tkeep = dm_tkeep[71][M_AXIS_OARG_71_DMWIDTH/8-1:0];
            assign m_axis_oarg_71_tstrb = dm_tstrb[71][M_AXIS_OARG_71_DMWIDTH/8-1:0];
            assign m_axis_oarg_71_tdata = dm_tdata[71][M_AXIS_OARG_71_DMWIDTH-1:0];
            assign ap_axis_oarg_71_tready = ap_tready[71];
            assign ap_tlast[71] = ap_axis_oarg_71_tlast;
            assign ap_tvalid[71] = ap_axis_oarg_71_tvalid;
            assign ap_tdata[71][M_AXIS_OARG_71_WIDTH-1:0] = ap_axis_oarg_71_tdata;
            assign ap_tkeep[71] = {M_AXIS_OARG_71_WIDTH/8{1'b1}};
            assign ap_tstrb[71] = {M_AXIS_OARG_71_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 72) begin
            assign axis_clk[72] = m_axis_oarg_72_aclk;
            assign axis_rst[72] = m_axis_oarg_72_aresetn;
            assign dm_tready[72] = m_axis_oarg_72_tready;
            assign m_axis_oarg_72_tlast = dm_tlast[72];
            assign m_axis_oarg_72_tvalid = dm_tvalid[72];
            assign m_axis_oarg_72_tkeep = dm_tkeep[72][M_AXIS_OARG_72_DMWIDTH/8-1:0];
            assign m_axis_oarg_72_tstrb = dm_tstrb[72][M_AXIS_OARG_72_DMWIDTH/8-1:0];
            assign m_axis_oarg_72_tdata = dm_tdata[72][M_AXIS_OARG_72_DMWIDTH-1:0];
            assign ap_axis_oarg_72_tready = ap_tready[72];
            assign ap_tlast[72] = ap_axis_oarg_72_tlast;
            assign ap_tvalid[72] = ap_axis_oarg_72_tvalid;
            assign ap_tdata[72][M_AXIS_OARG_72_WIDTH-1:0] = ap_axis_oarg_72_tdata;
            assign ap_tkeep[72] = {M_AXIS_OARG_72_WIDTH/8{1'b1}};
            assign ap_tstrb[72] = {M_AXIS_OARG_72_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 73) begin
            assign axis_clk[73] = m_axis_oarg_73_aclk;
            assign axis_rst[73] = m_axis_oarg_73_aresetn;
            assign dm_tready[73] = m_axis_oarg_73_tready;
            assign m_axis_oarg_73_tlast = dm_tlast[73];
            assign m_axis_oarg_73_tvalid = dm_tvalid[73];
            assign m_axis_oarg_73_tkeep = dm_tkeep[73][M_AXIS_OARG_73_DMWIDTH/8-1:0];
            assign m_axis_oarg_73_tstrb = dm_tstrb[73][M_AXIS_OARG_73_DMWIDTH/8-1:0];
            assign m_axis_oarg_73_tdata = dm_tdata[73][M_AXIS_OARG_73_DMWIDTH-1:0];
            assign ap_axis_oarg_73_tready = ap_tready[73];
            assign ap_tlast[73] = ap_axis_oarg_73_tlast;
            assign ap_tvalid[73] = ap_axis_oarg_73_tvalid;
            assign ap_tdata[73][M_AXIS_OARG_73_WIDTH-1:0] = ap_axis_oarg_73_tdata;
            assign ap_tkeep[73] = {M_AXIS_OARG_73_WIDTH/8{1'b1}};
            assign ap_tstrb[73] = {M_AXIS_OARG_73_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 74) begin
            assign axis_clk[74] = m_axis_oarg_74_aclk;
            assign axis_rst[74] = m_axis_oarg_74_aresetn;
            assign dm_tready[74] = m_axis_oarg_74_tready;
            assign m_axis_oarg_74_tlast = dm_tlast[74];
            assign m_axis_oarg_74_tvalid = dm_tvalid[74];
            assign m_axis_oarg_74_tkeep = dm_tkeep[74][M_AXIS_OARG_74_DMWIDTH/8-1:0];
            assign m_axis_oarg_74_tstrb = dm_tstrb[74][M_AXIS_OARG_74_DMWIDTH/8-1:0];
            assign m_axis_oarg_74_tdata = dm_tdata[74][M_AXIS_OARG_74_DMWIDTH-1:0];
            assign ap_axis_oarg_74_tready = ap_tready[74];
            assign ap_tlast[74] = ap_axis_oarg_74_tlast;
            assign ap_tvalid[74] = ap_axis_oarg_74_tvalid;
            assign ap_tdata[74][M_AXIS_OARG_74_WIDTH-1:0] = ap_axis_oarg_74_tdata;
            assign ap_tkeep[74] = {M_AXIS_OARG_74_WIDTH/8{1'b1}};
            assign ap_tstrb[74] = {M_AXIS_OARG_74_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 75) begin
            assign axis_clk[75] = m_axis_oarg_75_aclk;
            assign axis_rst[75] = m_axis_oarg_75_aresetn;
            assign dm_tready[75] = m_axis_oarg_75_tready;
            assign m_axis_oarg_75_tlast = dm_tlast[75];
            assign m_axis_oarg_75_tvalid = dm_tvalid[75];
            assign m_axis_oarg_75_tkeep = dm_tkeep[75][M_AXIS_OARG_75_DMWIDTH/8-1:0];
            assign m_axis_oarg_75_tstrb = dm_tstrb[75][M_AXIS_OARG_75_DMWIDTH/8-1:0];
            assign m_axis_oarg_75_tdata = dm_tdata[75][M_AXIS_OARG_75_DMWIDTH-1:0];
            assign ap_axis_oarg_75_tready = ap_tready[75];
            assign ap_tlast[75] = ap_axis_oarg_75_tlast;
            assign ap_tvalid[75] = ap_axis_oarg_75_tvalid;
            assign ap_tdata[75][M_AXIS_OARG_75_WIDTH-1:0] = ap_axis_oarg_75_tdata;
            assign ap_tkeep[75] = {M_AXIS_OARG_75_WIDTH/8{1'b1}};
            assign ap_tstrb[75] = {M_AXIS_OARG_75_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 76) begin
            assign axis_clk[76] = m_axis_oarg_76_aclk;
            assign axis_rst[76] = m_axis_oarg_76_aresetn;
            assign dm_tready[76] = m_axis_oarg_76_tready;
            assign m_axis_oarg_76_tlast = dm_tlast[76];
            assign m_axis_oarg_76_tvalid = dm_tvalid[76];
            assign m_axis_oarg_76_tkeep = dm_tkeep[76][M_AXIS_OARG_76_DMWIDTH/8-1:0];
            assign m_axis_oarg_76_tstrb = dm_tstrb[76][M_AXIS_OARG_76_DMWIDTH/8-1:0];
            assign m_axis_oarg_76_tdata = dm_tdata[76][M_AXIS_OARG_76_DMWIDTH-1:0];
            assign ap_axis_oarg_76_tready = ap_tready[76];
            assign ap_tlast[76] = ap_axis_oarg_76_tlast;
            assign ap_tvalid[76] = ap_axis_oarg_76_tvalid;
            assign ap_tdata[76][M_AXIS_OARG_76_WIDTH-1:0] = ap_axis_oarg_76_tdata;
            assign ap_tkeep[76] = {M_AXIS_OARG_76_WIDTH/8{1'b1}};
            assign ap_tstrb[76] = {M_AXIS_OARG_76_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 77) begin
            assign axis_clk[77] = m_axis_oarg_77_aclk;
            assign axis_rst[77] = m_axis_oarg_77_aresetn;
            assign dm_tready[77] = m_axis_oarg_77_tready;
            assign m_axis_oarg_77_tlast = dm_tlast[77];
            assign m_axis_oarg_77_tvalid = dm_tvalid[77];
            assign m_axis_oarg_77_tkeep = dm_tkeep[77][M_AXIS_OARG_77_DMWIDTH/8-1:0];
            assign m_axis_oarg_77_tstrb = dm_tstrb[77][M_AXIS_OARG_77_DMWIDTH/8-1:0];
            assign m_axis_oarg_77_tdata = dm_tdata[77][M_AXIS_OARG_77_DMWIDTH-1:0];
            assign ap_axis_oarg_77_tready = ap_tready[77];
            assign ap_tlast[77] = ap_axis_oarg_77_tlast;
            assign ap_tvalid[77] = ap_axis_oarg_77_tvalid;
            assign ap_tdata[77][M_AXIS_OARG_77_WIDTH-1:0] = ap_axis_oarg_77_tdata;
            assign ap_tkeep[77] = {M_AXIS_OARG_77_WIDTH/8{1'b1}};
            assign ap_tstrb[77] = {M_AXIS_OARG_77_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 78) begin
            assign axis_clk[78] = m_axis_oarg_78_aclk;
            assign axis_rst[78] = m_axis_oarg_78_aresetn;
            assign dm_tready[78] = m_axis_oarg_78_tready;
            assign m_axis_oarg_78_tlast = dm_tlast[78];
            assign m_axis_oarg_78_tvalid = dm_tvalid[78];
            assign m_axis_oarg_78_tkeep = dm_tkeep[78][M_AXIS_OARG_78_DMWIDTH/8-1:0];
            assign m_axis_oarg_78_tstrb = dm_tstrb[78][M_AXIS_OARG_78_DMWIDTH/8-1:0];
            assign m_axis_oarg_78_tdata = dm_tdata[78][M_AXIS_OARG_78_DMWIDTH-1:0];
            assign ap_axis_oarg_78_tready = ap_tready[78];
            assign ap_tlast[78] = ap_axis_oarg_78_tlast;
            assign ap_tvalid[78] = ap_axis_oarg_78_tvalid;
            assign ap_tdata[78][M_AXIS_OARG_78_WIDTH-1:0] = ap_axis_oarg_78_tdata;
            assign ap_tkeep[78] = {M_AXIS_OARG_78_WIDTH/8{1'b1}};
            assign ap_tstrb[78] = {M_AXIS_OARG_78_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 79) begin
            assign axis_clk[79] = m_axis_oarg_79_aclk;
            assign axis_rst[79] = m_axis_oarg_79_aresetn;
            assign dm_tready[79] = m_axis_oarg_79_tready;
            assign m_axis_oarg_79_tlast = dm_tlast[79];
            assign m_axis_oarg_79_tvalid = dm_tvalid[79];
            assign m_axis_oarg_79_tkeep = dm_tkeep[79][M_AXIS_OARG_79_DMWIDTH/8-1:0];
            assign m_axis_oarg_79_tstrb = dm_tstrb[79][M_AXIS_OARG_79_DMWIDTH/8-1:0];
            assign m_axis_oarg_79_tdata = dm_tdata[79][M_AXIS_OARG_79_DMWIDTH-1:0];
            assign ap_axis_oarg_79_tready = ap_tready[79];
            assign ap_tlast[79] = ap_axis_oarg_79_tlast;
            assign ap_tvalid[79] = ap_axis_oarg_79_tvalid;
            assign ap_tdata[79][M_AXIS_OARG_79_WIDTH-1:0] = ap_axis_oarg_79_tdata;
            assign ap_tkeep[79] = {M_AXIS_OARG_79_WIDTH/8{1'b1}};
            assign ap_tstrb[79] = {M_AXIS_OARG_79_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 80) begin
            assign axis_clk[80] = m_axis_oarg_80_aclk;
            assign axis_rst[80] = m_axis_oarg_80_aresetn;
            assign dm_tready[80] = m_axis_oarg_80_tready;
            assign m_axis_oarg_80_tlast = dm_tlast[80];
            assign m_axis_oarg_80_tvalid = dm_tvalid[80];
            assign m_axis_oarg_80_tkeep = dm_tkeep[80][M_AXIS_OARG_80_DMWIDTH/8-1:0];
            assign m_axis_oarg_80_tstrb = dm_tstrb[80][M_AXIS_OARG_80_DMWIDTH/8-1:0];
            assign m_axis_oarg_80_tdata = dm_tdata[80][M_AXIS_OARG_80_DMWIDTH-1:0];
            assign ap_axis_oarg_80_tready = ap_tready[80];
            assign ap_tlast[80] = ap_axis_oarg_80_tlast;
            assign ap_tvalid[80] = ap_axis_oarg_80_tvalid;
            assign ap_tdata[80][M_AXIS_OARG_80_WIDTH-1:0] = ap_axis_oarg_80_tdata;
            assign ap_tkeep[80] = {M_AXIS_OARG_80_WIDTH/8{1'b1}};
            assign ap_tstrb[80] = {M_AXIS_OARG_80_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 81) begin
            assign axis_clk[81] = m_axis_oarg_81_aclk;
            assign axis_rst[81] = m_axis_oarg_81_aresetn;
            assign dm_tready[81] = m_axis_oarg_81_tready;
            assign m_axis_oarg_81_tlast = dm_tlast[81];
            assign m_axis_oarg_81_tvalid = dm_tvalid[81];
            assign m_axis_oarg_81_tkeep = dm_tkeep[81][M_AXIS_OARG_81_DMWIDTH/8-1:0];
            assign m_axis_oarg_81_tstrb = dm_tstrb[81][M_AXIS_OARG_81_DMWIDTH/8-1:0];
            assign m_axis_oarg_81_tdata = dm_tdata[81][M_AXIS_OARG_81_DMWIDTH-1:0];
            assign ap_axis_oarg_81_tready = ap_tready[81];
            assign ap_tlast[81] = ap_axis_oarg_81_tlast;
            assign ap_tvalid[81] = ap_axis_oarg_81_tvalid;
            assign ap_tdata[81][M_AXIS_OARG_81_WIDTH-1:0] = ap_axis_oarg_81_tdata;
            assign ap_tkeep[81] = {M_AXIS_OARG_81_WIDTH/8{1'b1}};
            assign ap_tstrb[81] = {M_AXIS_OARG_81_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 82) begin
            assign axis_clk[82] = m_axis_oarg_82_aclk;
            assign axis_rst[82] = m_axis_oarg_82_aresetn;
            assign dm_tready[82] = m_axis_oarg_82_tready;
            assign m_axis_oarg_82_tlast = dm_tlast[82];
            assign m_axis_oarg_82_tvalid = dm_tvalid[82];
            assign m_axis_oarg_82_tkeep = dm_tkeep[82][M_AXIS_OARG_82_DMWIDTH/8-1:0];
            assign m_axis_oarg_82_tstrb = dm_tstrb[82][M_AXIS_OARG_82_DMWIDTH/8-1:0];
            assign m_axis_oarg_82_tdata = dm_tdata[82][M_AXIS_OARG_82_DMWIDTH-1:0];
            assign ap_axis_oarg_82_tready = ap_tready[82];
            assign ap_tlast[82] = ap_axis_oarg_82_tlast;
            assign ap_tvalid[82] = ap_axis_oarg_82_tvalid;
            assign ap_tdata[82][M_AXIS_OARG_82_WIDTH-1:0] = ap_axis_oarg_82_tdata;
            assign ap_tkeep[82] = {M_AXIS_OARG_82_WIDTH/8{1'b1}};
            assign ap_tstrb[82] = {M_AXIS_OARG_82_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 83) begin
            assign axis_clk[83] = m_axis_oarg_83_aclk;
            assign axis_rst[83] = m_axis_oarg_83_aresetn;
            assign dm_tready[83] = m_axis_oarg_83_tready;
            assign m_axis_oarg_83_tlast = dm_tlast[83];
            assign m_axis_oarg_83_tvalid = dm_tvalid[83];
            assign m_axis_oarg_83_tkeep = dm_tkeep[83][M_AXIS_OARG_83_DMWIDTH/8-1:0];
            assign m_axis_oarg_83_tstrb = dm_tstrb[83][M_AXIS_OARG_83_DMWIDTH/8-1:0];
            assign m_axis_oarg_83_tdata = dm_tdata[83][M_AXIS_OARG_83_DMWIDTH-1:0];
            assign ap_axis_oarg_83_tready = ap_tready[83];
            assign ap_tlast[83] = ap_axis_oarg_83_tlast;
            assign ap_tvalid[83] = ap_axis_oarg_83_tvalid;
            assign ap_tdata[83][M_AXIS_OARG_83_WIDTH-1:0] = ap_axis_oarg_83_tdata;
            assign ap_tkeep[83] = {M_AXIS_OARG_83_WIDTH/8{1'b1}};
            assign ap_tstrb[83] = {M_AXIS_OARG_83_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 84) begin
            assign axis_clk[84] = m_axis_oarg_84_aclk;
            assign axis_rst[84] = m_axis_oarg_84_aresetn;
            assign dm_tready[84] = m_axis_oarg_84_tready;
            assign m_axis_oarg_84_tlast = dm_tlast[84];
            assign m_axis_oarg_84_tvalid = dm_tvalid[84];
            assign m_axis_oarg_84_tkeep = dm_tkeep[84][M_AXIS_OARG_84_DMWIDTH/8-1:0];
            assign m_axis_oarg_84_tstrb = dm_tstrb[84][M_AXIS_OARG_84_DMWIDTH/8-1:0];
            assign m_axis_oarg_84_tdata = dm_tdata[84][M_AXIS_OARG_84_DMWIDTH-1:0];
            assign ap_axis_oarg_84_tready = ap_tready[84];
            assign ap_tlast[84] = ap_axis_oarg_84_tlast;
            assign ap_tvalid[84] = ap_axis_oarg_84_tvalid;
            assign ap_tdata[84][M_AXIS_OARG_84_WIDTH-1:0] = ap_axis_oarg_84_tdata;
            assign ap_tkeep[84] = {M_AXIS_OARG_84_WIDTH/8{1'b1}};
            assign ap_tstrb[84] = {M_AXIS_OARG_84_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 85) begin
            assign axis_clk[85] = m_axis_oarg_85_aclk;
            assign axis_rst[85] = m_axis_oarg_85_aresetn;
            assign dm_tready[85] = m_axis_oarg_85_tready;
            assign m_axis_oarg_85_tlast = dm_tlast[85];
            assign m_axis_oarg_85_tvalid = dm_tvalid[85];
            assign m_axis_oarg_85_tkeep = dm_tkeep[85][M_AXIS_OARG_85_DMWIDTH/8-1:0];
            assign m_axis_oarg_85_tstrb = dm_tstrb[85][M_AXIS_OARG_85_DMWIDTH/8-1:0];
            assign m_axis_oarg_85_tdata = dm_tdata[85][M_AXIS_OARG_85_DMWIDTH-1:0];
            assign ap_axis_oarg_85_tready = ap_tready[85];
            assign ap_tlast[85] = ap_axis_oarg_85_tlast;
            assign ap_tvalid[85] = ap_axis_oarg_85_tvalid;
            assign ap_tdata[85][M_AXIS_OARG_85_WIDTH-1:0] = ap_axis_oarg_85_tdata;
            assign ap_tkeep[85] = {M_AXIS_OARG_85_WIDTH/8{1'b1}};
            assign ap_tstrb[85] = {M_AXIS_OARG_85_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 86) begin
            assign axis_clk[86] = m_axis_oarg_86_aclk;
            assign axis_rst[86] = m_axis_oarg_86_aresetn;
            assign dm_tready[86] = m_axis_oarg_86_tready;
            assign m_axis_oarg_86_tlast = dm_tlast[86];
            assign m_axis_oarg_86_tvalid = dm_tvalid[86];
            assign m_axis_oarg_86_tkeep = dm_tkeep[86][M_AXIS_OARG_86_DMWIDTH/8-1:0];
            assign m_axis_oarg_86_tstrb = dm_tstrb[86][M_AXIS_OARG_86_DMWIDTH/8-1:0];
            assign m_axis_oarg_86_tdata = dm_tdata[86][M_AXIS_OARG_86_DMWIDTH-1:0];
            assign ap_axis_oarg_86_tready = ap_tready[86];
            assign ap_tlast[86] = ap_axis_oarg_86_tlast;
            assign ap_tvalid[86] = ap_axis_oarg_86_tvalid;
            assign ap_tdata[86][M_AXIS_OARG_86_WIDTH-1:0] = ap_axis_oarg_86_tdata;
            assign ap_tkeep[86] = {M_AXIS_OARG_86_WIDTH/8{1'b1}};
            assign ap_tstrb[86] = {M_AXIS_OARG_86_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 87) begin
            assign axis_clk[87] = m_axis_oarg_87_aclk;
            assign axis_rst[87] = m_axis_oarg_87_aresetn;
            assign dm_tready[87] = m_axis_oarg_87_tready;
            assign m_axis_oarg_87_tlast = dm_tlast[87];
            assign m_axis_oarg_87_tvalid = dm_tvalid[87];
            assign m_axis_oarg_87_tkeep = dm_tkeep[87][M_AXIS_OARG_87_DMWIDTH/8-1:0];
            assign m_axis_oarg_87_tstrb = dm_tstrb[87][M_AXIS_OARG_87_DMWIDTH/8-1:0];
            assign m_axis_oarg_87_tdata = dm_tdata[87][M_AXIS_OARG_87_DMWIDTH-1:0];
            assign ap_axis_oarg_87_tready = ap_tready[87];
            assign ap_tlast[87] = ap_axis_oarg_87_tlast;
            assign ap_tvalid[87] = ap_axis_oarg_87_tvalid;
            assign ap_tdata[87][M_AXIS_OARG_87_WIDTH-1:0] = ap_axis_oarg_87_tdata;
            assign ap_tkeep[87] = {M_AXIS_OARG_87_WIDTH/8{1'b1}};
            assign ap_tstrb[87] = {M_AXIS_OARG_87_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 88) begin
            assign axis_clk[88] = m_axis_oarg_88_aclk;
            assign axis_rst[88] = m_axis_oarg_88_aresetn;
            assign dm_tready[88] = m_axis_oarg_88_tready;
            assign m_axis_oarg_88_tlast = dm_tlast[88];
            assign m_axis_oarg_88_tvalid = dm_tvalid[88];
            assign m_axis_oarg_88_tkeep = dm_tkeep[88][M_AXIS_OARG_88_DMWIDTH/8-1:0];
            assign m_axis_oarg_88_tstrb = dm_tstrb[88][M_AXIS_OARG_88_DMWIDTH/8-1:0];
            assign m_axis_oarg_88_tdata = dm_tdata[88][M_AXIS_OARG_88_DMWIDTH-1:0];
            assign ap_axis_oarg_88_tready = ap_tready[88];
            assign ap_tlast[88] = ap_axis_oarg_88_tlast;
            assign ap_tvalid[88] = ap_axis_oarg_88_tvalid;
            assign ap_tdata[88][M_AXIS_OARG_88_WIDTH-1:0] = ap_axis_oarg_88_tdata;
            assign ap_tkeep[88] = {M_AXIS_OARG_88_WIDTH/8{1'b1}};
            assign ap_tstrb[88] = {M_AXIS_OARG_88_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 89) begin
            assign axis_clk[89] = m_axis_oarg_89_aclk;
            assign axis_rst[89] = m_axis_oarg_89_aresetn;
            assign dm_tready[89] = m_axis_oarg_89_tready;
            assign m_axis_oarg_89_tlast = dm_tlast[89];
            assign m_axis_oarg_89_tvalid = dm_tvalid[89];
            assign m_axis_oarg_89_tkeep = dm_tkeep[89][M_AXIS_OARG_89_DMWIDTH/8-1:0];
            assign m_axis_oarg_89_tstrb = dm_tstrb[89][M_AXIS_OARG_89_DMWIDTH/8-1:0];
            assign m_axis_oarg_89_tdata = dm_tdata[89][M_AXIS_OARG_89_DMWIDTH-1:0];
            assign ap_axis_oarg_89_tready = ap_tready[89];
            assign ap_tlast[89] = ap_axis_oarg_89_tlast;
            assign ap_tvalid[89] = ap_axis_oarg_89_tvalid;
            assign ap_tdata[89][M_AXIS_OARG_89_WIDTH-1:0] = ap_axis_oarg_89_tdata;
            assign ap_tkeep[89] = {M_AXIS_OARG_89_WIDTH/8{1'b1}};
            assign ap_tstrb[89] = {M_AXIS_OARG_89_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 90) begin
            assign axis_clk[90] = m_axis_oarg_90_aclk;
            assign axis_rst[90] = m_axis_oarg_90_aresetn;
            assign dm_tready[90] = m_axis_oarg_90_tready;
            assign m_axis_oarg_90_tlast = dm_tlast[90];
            assign m_axis_oarg_90_tvalid = dm_tvalid[90];
            assign m_axis_oarg_90_tkeep = dm_tkeep[90][M_AXIS_OARG_90_DMWIDTH/8-1:0];
            assign m_axis_oarg_90_tstrb = dm_tstrb[90][M_AXIS_OARG_90_DMWIDTH/8-1:0];
            assign m_axis_oarg_90_tdata = dm_tdata[90][M_AXIS_OARG_90_DMWIDTH-1:0];
            assign ap_axis_oarg_90_tready = ap_tready[90];
            assign ap_tlast[90] = ap_axis_oarg_90_tlast;
            assign ap_tvalid[90] = ap_axis_oarg_90_tvalid;
            assign ap_tdata[90][M_AXIS_OARG_90_WIDTH-1:0] = ap_axis_oarg_90_tdata;
            assign ap_tkeep[90] = {M_AXIS_OARG_90_WIDTH/8{1'b1}};
            assign ap_tstrb[90] = {M_AXIS_OARG_90_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 91) begin
            assign axis_clk[91] = m_axis_oarg_91_aclk;
            assign axis_rst[91] = m_axis_oarg_91_aresetn;
            assign dm_tready[91] = m_axis_oarg_91_tready;
            assign m_axis_oarg_91_tlast = dm_tlast[91];
            assign m_axis_oarg_91_tvalid = dm_tvalid[91];
            assign m_axis_oarg_91_tkeep = dm_tkeep[91][M_AXIS_OARG_91_DMWIDTH/8-1:0];
            assign m_axis_oarg_91_tstrb = dm_tstrb[91][M_AXIS_OARG_91_DMWIDTH/8-1:0];
            assign m_axis_oarg_91_tdata = dm_tdata[91][M_AXIS_OARG_91_DMWIDTH-1:0];
            assign ap_axis_oarg_91_tready = ap_tready[91];
            assign ap_tlast[91] = ap_axis_oarg_91_tlast;
            assign ap_tvalid[91] = ap_axis_oarg_91_tvalid;
            assign ap_tdata[91][M_AXIS_OARG_91_WIDTH-1:0] = ap_axis_oarg_91_tdata;
            assign ap_tkeep[91] = {M_AXIS_OARG_91_WIDTH/8{1'b1}};
            assign ap_tstrb[91] = {M_AXIS_OARG_91_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 92) begin
            assign axis_clk[92] = m_axis_oarg_92_aclk;
            assign axis_rst[92] = m_axis_oarg_92_aresetn;
            assign dm_tready[92] = m_axis_oarg_92_tready;
            assign m_axis_oarg_92_tlast = dm_tlast[92];
            assign m_axis_oarg_92_tvalid = dm_tvalid[92];
            assign m_axis_oarg_92_tkeep = dm_tkeep[92][M_AXIS_OARG_92_DMWIDTH/8-1:0];
            assign m_axis_oarg_92_tstrb = dm_tstrb[92][M_AXIS_OARG_92_DMWIDTH/8-1:0];
            assign m_axis_oarg_92_tdata = dm_tdata[92][M_AXIS_OARG_92_DMWIDTH-1:0];
            assign ap_axis_oarg_92_tready = ap_tready[92];
            assign ap_tlast[92] = ap_axis_oarg_92_tlast;
            assign ap_tvalid[92] = ap_axis_oarg_92_tvalid;
            assign ap_tdata[92][M_AXIS_OARG_92_WIDTH-1:0] = ap_axis_oarg_92_tdata;
            assign ap_tkeep[92] = {M_AXIS_OARG_92_WIDTH/8{1'b1}};
            assign ap_tstrb[92] = {M_AXIS_OARG_92_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 93) begin
            assign axis_clk[93] = m_axis_oarg_93_aclk;
            assign axis_rst[93] = m_axis_oarg_93_aresetn;
            assign dm_tready[93] = m_axis_oarg_93_tready;
            assign m_axis_oarg_93_tlast = dm_tlast[93];
            assign m_axis_oarg_93_tvalid = dm_tvalid[93];
            assign m_axis_oarg_93_tkeep = dm_tkeep[93][M_AXIS_OARG_93_DMWIDTH/8-1:0];
            assign m_axis_oarg_93_tstrb = dm_tstrb[93][M_AXIS_OARG_93_DMWIDTH/8-1:0];
            assign m_axis_oarg_93_tdata = dm_tdata[93][M_AXIS_OARG_93_DMWIDTH-1:0];
            assign ap_axis_oarg_93_tready = ap_tready[93];
            assign ap_tlast[93] = ap_axis_oarg_93_tlast;
            assign ap_tvalid[93] = ap_axis_oarg_93_tvalid;
            assign ap_tdata[93][M_AXIS_OARG_93_WIDTH-1:0] = ap_axis_oarg_93_tdata;
            assign ap_tkeep[93] = {M_AXIS_OARG_93_WIDTH/8{1'b1}};
            assign ap_tstrb[93] = {M_AXIS_OARG_93_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 94) begin
            assign axis_clk[94] = m_axis_oarg_94_aclk;
            assign axis_rst[94] = m_axis_oarg_94_aresetn;
            assign dm_tready[94] = m_axis_oarg_94_tready;
            assign m_axis_oarg_94_tlast = dm_tlast[94];
            assign m_axis_oarg_94_tvalid = dm_tvalid[94];
            assign m_axis_oarg_94_tkeep = dm_tkeep[94][M_AXIS_OARG_94_DMWIDTH/8-1:0];
            assign m_axis_oarg_94_tstrb = dm_tstrb[94][M_AXIS_OARG_94_DMWIDTH/8-1:0];
            assign m_axis_oarg_94_tdata = dm_tdata[94][M_AXIS_OARG_94_DMWIDTH-1:0];
            assign ap_axis_oarg_94_tready = ap_tready[94];
            assign ap_tlast[94] = ap_axis_oarg_94_tlast;
            assign ap_tvalid[94] = ap_axis_oarg_94_tvalid;
            assign ap_tdata[94][M_AXIS_OARG_94_WIDTH-1:0] = ap_axis_oarg_94_tdata;
            assign ap_tkeep[94] = {M_AXIS_OARG_94_WIDTH/8{1'b1}};
            assign ap_tstrb[94] = {M_AXIS_OARG_94_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 95) begin
            assign axis_clk[95] = m_axis_oarg_95_aclk;
            assign axis_rst[95] = m_axis_oarg_95_aresetn;
            assign dm_tready[95] = m_axis_oarg_95_tready;
            assign m_axis_oarg_95_tlast = dm_tlast[95];
            assign m_axis_oarg_95_tvalid = dm_tvalid[95];
            assign m_axis_oarg_95_tkeep = dm_tkeep[95][M_AXIS_OARG_95_DMWIDTH/8-1:0];
            assign m_axis_oarg_95_tstrb = dm_tstrb[95][M_AXIS_OARG_95_DMWIDTH/8-1:0];
            assign m_axis_oarg_95_tdata = dm_tdata[95][M_AXIS_OARG_95_DMWIDTH-1:0];
            assign ap_axis_oarg_95_tready = ap_tready[95];
            assign ap_tlast[95] = ap_axis_oarg_95_tlast;
            assign ap_tvalid[95] = ap_axis_oarg_95_tvalid;
            assign ap_tdata[95][M_AXIS_OARG_95_WIDTH-1:0] = ap_axis_oarg_95_tdata;
            assign ap_tkeep[95] = {M_AXIS_OARG_95_WIDTH/8{1'b1}};
            assign ap_tstrb[95] = {M_AXIS_OARG_95_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 96) begin
            assign axis_clk[96] = m_axis_oarg_96_aclk;
            assign axis_rst[96] = m_axis_oarg_96_aresetn;
            assign dm_tready[96] = m_axis_oarg_96_tready;
            assign m_axis_oarg_96_tlast = dm_tlast[96];
            assign m_axis_oarg_96_tvalid = dm_tvalid[96];
            assign m_axis_oarg_96_tkeep = dm_tkeep[96][M_AXIS_OARG_96_DMWIDTH/8-1:0];
            assign m_axis_oarg_96_tstrb = dm_tstrb[96][M_AXIS_OARG_96_DMWIDTH/8-1:0];
            assign m_axis_oarg_96_tdata = dm_tdata[96][M_AXIS_OARG_96_DMWIDTH-1:0];
            assign ap_axis_oarg_96_tready = ap_tready[96];
            assign ap_tlast[96] = ap_axis_oarg_96_tlast;
            assign ap_tvalid[96] = ap_axis_oarg_96_tvalid;
            assign ap_tdata[96][M_AXIS_OARG_96_WIDTH-1:0] = ap_axis_oarg_96_tdata;
            assign ap_tkeep[96] = {M_AXIS_OARG_96_WIDTH/8{1'b1}};
            assign ap_tstrb[96] = {M_AXIS_OARG_96_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 97) begin
            assign axis_clk[97] = m_axis_oarg_97_aclk;
            assign axis_rst[97] = m_axis_oarg_97_aresetn;
            assign dm_tready[97] = m_axis_oarg_97_tready;
            assign m_axis_oarg_97_tlast = dm_tlast[97];
            assign m_axis_oarg_97_tvalid = dm_tvalid[97];
            assign m_axis_oarg_97_tkeep = dm_tkeep[97][M_AXIS_OARG_97_DMWIDTH/8-1:0];
            assign m_axis_oarg_97_tstrb = dm_tstrb[97][M_AXIS_OARG_97_DMWIDTH/8-1:0];
            assign m_axis_oarg_97_tdata = dm_tdata[97][M_AXIS_OARG_97_DMWIDTH-1:0];
            assign ap_axis_oarg_97_tready = ap_tready[97];
            assign ap_tlast[97] = ap_axis_oarg_97_tlast;
            assign ap_tvalid[97] = ap_axis_oarg_97_tvalid;
            assign ap_tdata[97][M_AXIS_OARG_97_WIDTH-1:0] = ap_axis_oarg_97_tdata;
            assign ap_tkeep[97] = {M_AXIS_OARG_97_WIDTH/8{1'b1}};
            assign ap_tstrb[97] = {M_AXIS_OARG_97_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 98) begin
            assign axis_clk[98] = m_axis_oarg_98_aclk;
            assign axis_rst[98] = m_axis_oarg_98_aresetn;
            assign dm_tready[98] = m_axis_oarg_98_tready;
            assign m_axis_oarg_98_tlast = dm_tlast[98];
            assign m_axis_oarg_98_tvalid = dm_tvalid[98];
            assign m_axis_oarg_98_tkeep = dm_tkeep[98][M_AXIS_OARG_98_DMWIDTH/8-1:0];
            assign m_axis_oarg_98_tstrb = dm_tstrb[98][M_AXIS_OARG_98_DMWIDTH/8-1:0];
            assign m_axis_oarg_98_tdata = dm_tdata[98][M_AXIS_OARG_98_DMWIDTH-1:0];
            assign ap_axis_oarg_98_tready = ap_tready[98];
            assign ap_tlast[98] = ap_axis_oarg_98_tlast;
            assign ap_tvalid[98] = ap_axis_oarg_98_tvalid;
            assign ap_tdata[98][M_AXIS_OARG_98_WIDTH-1:0] = ap_axis_oarg_98_tdata;
            assign ap_tkeep[98] = {M_AXIS_OARG_98_WIDTH/8{1'b1}};
            assign ap_tstrb[98] = {M_AXIS_OARG_98_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 99) begin
            assign axis_clk[99] = m_axis_oarg_99_aclk;
            assign axis_rst[99] = m_axis_oarg_99_aresetn;
            assign dm_tready[99] = m_axis_oarg_99_tready;
            assign m_axis_oarg_99_tlast = dm_tlast[99];
            assign m_axis_oarg_99_tvalid = dm_tvalid[99];
            assign m_axis_oarg_99_tkeep = dm_tkeep[99][M_AXIS_OARG_99_DMWIDTH/8-1:0];
            assign m_axis_oarg_99_tstrb = dm_tstrb[99][M_AXIS_OARG_99_DMWIDTH/8-1:0];
            assign m_axis_oarg_99_tdata = dm_tdata[99][M_AXIS_OARG_99_DMWIDTH-1:0];
            assign ap_axis_oarg_99_tready = ap_tready[99];
            assign ap_tlast[99] = ap_axis_oarg_99_tlast;
            assign ap_tvalid[99] = ap_axis_oarg_99_tvalid;
            assign ap_tdata[99][M_AXIS_OARG_99_WIDTH-1:0] = ap_axis_oarg_99_tdata;
            assign ap_tkeep[99] = {M_AXIS_OARG_99_WIDTH/8{1'b1}};
            assign ap_tstrb[99] = {M_AXIS_OARG_99_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 100) begin
            assign axis_clk[100] = m_axis_oarg_100_aclk;
            assign axis_rst[100] = m_axis_oarg_100_aresetn;
            assign dm_tready[100] = m_axis_oarg_100_tready;
            assign m_axis_oarg_100_tlast = dm_tlast[100];
            assign m_axis_oarg_100_tvalid = dm_tvalid[100];
            assign m_axis_oarg_100_tkeep = dm_tkeep[100][M_AXIS_OARG_100_DMWIDTH/8-1:0];
            assign m_axis_oarg_100_tstrb = dm_tstrb[100][M_AXIS_OARG_100_DMWIDTH/8-1:0];
            assign m_axis_oarg_100_tdata = dm_tdata[100][M_AXIS_OARG_100_DMWIDTH-1:0];
            assign ap_axis_oarg_100_tready = ap_tready[100];
            assign ap_tlast[100] = ap_axis_oarg_100_tlast;
            assign ap_tvalid[100] = ap_axis_oarg_100_tvalid;
            assign ap_tdata[100][M_AXIS_OARG_100_WIDTH-1:0] = ap_axis_oarg_100_tdata;
            assign ap_tkeep[100] = {M_AXIS_OARG_100_WIDTH/8{1'b1}};
            assign ap_tstrb[100] = {M_AXIS_OARG_100_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 101) begin
            assign axis_clk[101] = m_axis_oarg_101_aclk;
            assign axis_rst[101] = m_axis_oarg_101_aresetn;
            assign dm_tready[101] = m_axis_oarg_101_tready;
            assign m_axis_oarg_101_tlast = dm_tlast[101];
            assign m_axis_oarg_101_tvalid = dm_tvalid[101];
            assign m_axis_oarg_101_tkeep = dm_tkeep[101][M_AXIS_OARG_101_DMWIDTH/8-1:0];
            assign m_axis_oarg_101_tstrb = dm_tstrb[101][M_AXIS_OARG_101_DMWIDTH/8-1:0];
            assign m_axis_oarg_101_tdata = dm_tdata[101][M_AXIS_OARG_101_DMWIDTH-1:0];
            assign ap_axis_oarg_101_tready = ap_tready[101];
            assign ap_tlast[101] = ap_axis_oarg_101_tlast;
            assign ap_tvalid[101] = ap_axis_oarg_101_tvalid;
            assign ap_tdata[101][M_AXIS_OARG_101_WIDTH-1:0] = ap_axis_oarg_101_tdata;
            assign ap_tkeep[101] = {M_AXIS_OARG_101_WIDTH/8{1'b1}};
            assign ap_tstrb[101] = {M_AXIS_OARG_101_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 102) begin
            assign axis_clk[102] = m_axis_oarg_102_aclk;
            assign axis_rst[102] = m_axis_oarg_102_aresetn;
            assign dm_tready[102] = m_axis_oarg_102_tready;
            assign m_axis_oarg_102_tlast = dm_tlast[102];
            assign m_axis_oarg_102_tvalid = dm_tvalid[102];
            assign m_axis_oarg_102_tkeep = dm_tkeep[102][M_AXIS_OARG_102_DMWIDTH/8-1:0];
            assign m_axis_oarg_102_tstrb = dm_tstrb[102][M_AXIS_OARG_102_DMWIDTH/8-1:0];
            assign m_axis_oarg_102_tdata = dm_tdata[102][M_AXIS_OARG_102_DMWIDTH-1:0];
            assign ap_axis_oarg_102_tready = ap_tready[102];
            assign ap_tlast[102] = ap_axis_oarg_102_tlast;
            assign ap_tvalid[102] = ap_axis_oarg_102_tvalid;
            assign ap_tdata[102][M_AXIS_OARG_102_WIDTH-1:0] = ap_axis_oarg_102_tdata;
            assign ap_tkeep[102] = {M_AXIS_OARG_102_WIDTH/8{1'b1}};
            assign ap_tstrb[102] = {M_AXIS_OARG_102_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 103) begin
            assign axis_clk[103] = m_axis_oarg_103_aclk;
            assign axis_rst[103] = m_axis_oarg_103_aresetn;
            assign dm_tready[103] = m_axis_oarg_103_tready;
            assign m_axis_oarg_103_tlast = dm_tlast[103];
            assign m_axis_oarg_103_tvalid = dm_tvalid[103];
            assign m_axis_oarg_103_tkeep = dm_tkeep[103][M_AXIS_OARG_103_DMWIDTH/8-1:0];
            assign m_axis_oarg_103_tstrb = dm_tstrb[103][M_AXIS_OARG_103_DMWIDTH/8-1:0];
            assign m_axis_oarg_103_tdata = dm_tdata[103][M_AXIS_OARG_103_DMWIDTH-1:0];
            assign ap_axis_oarg_103_tready = ap_tready[103];
            assign ap_tlast[103] = ap_axis_oarg_103_tlast;
            assign ap_tvalid[103] = ap_axis_oarg_103_tvalid;
            assign ap_tdata[103][M_AXIS_OARG_103_WIDTH-1:0] = ap_axis_oarg_103_tdata;
            assign ap_tkeep[103] = {M_AXIS_OARG_103_WIDTH/8{1'b1}};
            assign ap_tstrb[103] = {M_AXIS_OARG_103_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 104) begin
            assign axis_clk[104] = m_axis_oarg_104_aclk;
            assign axis_rst[104] = m_axis_oarg_104_aresetn;
            assign dm_tready[104] = m_axis_oarg_104_tready;
            assign m_axis_oarg_104_tlast = dm_tlast[104];
            assign m_axis_oarg_104_tvalid = dm_tvalid[104];
            assign m_axis_oarg_104_tkeep = dm_tkeep[104][M_AXIS_OARG_104_DMWIDTH/8-1:0];
            assign m_axis_oarg_104_tstrb = dm_tstrb[104][M_AXIS_OARG_104_DMWIDTH/8-1:0];
            assign m_axis_oarg_104_tdata = dm_tdata[104][M_AXIS_OARG_104_DMWIDTH-1:0];
            assign ap_axis_oarg_104_tready = ap_tready[104];
            assign ap_tlast[104] = ap_axis_oarg_104_tlast;
            assign ap_tvalid[104] = ap_axis_oarg_104_tvalid;
            assign ap_tdata[104][M_AXIS_OARG_104_WIDTH-1:0] = ap_axis_oarg_104_tdata;
            assign ap_tkeep[104] = {M_AXIS_OARG_104_WIDTH/8{1'b1}};
            assign ap_tstrb[104] = {M_AXIS_OARG_104_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 105) begin
            assign axis_clk[105] = m_axis_oarg_105_aclk;
            assign axis_rst[105] = m_axis_oarg_105_aresetn;
            assign dm_tready[105] = m_axis_oarg_105_tready;
            assign m_axis_oarg_105_tlast = dm_tlast[105];
            assign m_axis_oarg_105_tvalid = dm_tvalid[105];
            assign m_axis_oarg_105_tkeep = dm_tkeep[105][M_AXIS_OARG_105_DMWIDTH/8-1:0];
            assign m_axis_oarg_105_tstrb = dm_tstrb[105][M_AXIS_OARG_105_DMWIDTH/8-1:0];
            assign m_axis_oarg_105_tdata = dm_tdata[105][M_AXIS_OARG_105_DMWIDTH-1:0];
            assign ap_axis_oarg_105_tready = ap_tready[105];
            assign ap_tlast[105] = ap_axis_oarg_105_tlast;
            assign ap_tvalid[105] = ap_axis_oarg_105_tvalid;
            assign ap_tdata[105][M_AXIS_OARG_105_WIDTH-1:0] = ap_axis_oarg_105_tdata;
            assign ap_tkeep[105] = {M_AXIS_OARG_105_WIDTH/8{1'b1}};
            assign ap_tstrb[105] = {M_AXIS_OARG_105_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 106) begin
            assign axis_clk[106] = m_axis_oarg_106_aclk;
            assign axis_rst[106] = m_axis_oarg_106_aresetn;
            assign dm_tready[106] = m_axis_oarg_106_tready;
            assign m_axis_oarg_106_tlast = dm_tlast[106];
            assign m_axis_oarg_106_tvalid = dm_tvalid[106];
            assign m_axis_oarg_106_tkeep = dm_tkeep[106][M_AXIS_OARG_106_DMWIDTH/8-1:0];
            assign m_axis_oarg_106_tstrb = dm_tstrb[106][M_AXIS_OARG_106_DMWIDTH/8-1:0];
            assign m_axis_oarg_106_tdata = dm_tdata[106][M_AXIS_OARG_106_DMWIDTH-1:0];
            assign ap_axis_oarg_106_tready = ap_tready[106];
            assign ap_tlast[106] = ap_axis_oarg_106_tlast;
            assign ap_tvalid[106] = ap_axis_oarg_106_tvalid;
            assign ap_tdata[106][M_AXIS_OARG_106_WIDTH-1:0] = ap_axis_oarg_106_tdata;
            assign ap_tkeep[106] = {M_AXIS_OARG_106_WIDTH/8{1'b1}};
            assign ap_tstrb[106] = {M_AXIS_OARG_106_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 107) begin
            assign axis_clk[107] = m_axis_oarg_107_aclk;
            assign axis_rst[107] = m_axis_oarg_107_aresetn;
            assign dm_tready[107] = m_axis_oarg_107_tready;
            assign m_axis_oarg_107_tlast = dm_tlast[107];
            assign m_axis_oarg_107_tvalid = dm_tvalid[107];
            assign m_axis_oarg_107_tkeep = dm_tkeep[107][M_AXIS_OARG_107_DMWIDTH/8-1:0];
            assign m_axis_oarg_107_tstrb = dm_tstrb[107][M_AXIS_OARG_107_DMWIDTH/8-1:0];
            assign m_axis_oarg_107_tdata = dm_tdata[107][M_AXIS_OARG_107_DMWIDTH-1:0];
            assign ap_axis_oarg_107_tready = ap_tready[107];
            assign ap_tlast[107] = ap_axis_oarg_107_tlast;
            assign ap_tvalid[107] = ap_axis_oarg_107_tvalid;
            assign ap_tdata[107][M_AXIS_OARG_107_WIDTH-1:0] = ap_axis_oarg_107_tdata;
            assign ap_tkeep[107] = {M_AXIS_OARG_107_WIDTH/8{1'b1}};
            assign ap_tstrb[107] = {M_AXIS_OARG_107_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 108) begin
            assign axis_clk[108] = m_axis_oarg_108_aclk;
            assign axis_rst[108] = m_axis_oarg_108_aresetn;
            assign dm_tready[108] = m_axis_oarg_108_tready;
            assign m_axis_oarg_108_tlast = dm_tlast[108];
            assign m_axis_oarg_108_tvalid = dm_tvalid[108];
            assign m_axis_oarg_108_tkeep = dm_tkeep[108][M_AXIS_OARG_108_DMWIDTH/8-1:0];
            assign m_axis_oarg_108_tstrb = dm_tstrb[108][M_AXIS_OARG_108_DMWIDTH/8-1:0];
            assign m_axis_oarg_108_tdata = dm_tdata[108][M_AXIS_OARG_108_DMWIDTH-1:0];
            assign ap_axis_oarg_108_tready = ap_tready[108];
            assign ap_tlast[108] = ap_axis_oarg_108_tlast;
            assign ap_tvalid[108] = ap_axis_oarg_108_tvalid;
            assign ap_tdata[108][M_AXIS_OARG_108_WIDTH-1:0] = ap_axis_oarg_108_tdata;
            assign ap_tkeep[108] = {M_AXIS_OARG_108_WIDTH/8{1'b1}};
            assign ap_tstrb[108] = {M_AXIS_OARG_108_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 109) begin
            assign axis_clk[109] = m_axis_oarg_109_aclk;
            assign axis_rst[109] = m_axis_oarg_109_aresetn;
            assign dm_tready[109] = m_axis_oarg_109_tready;
            assign m_axis_oarg_109_tlast = dm_tlast[109];
            assign m_axis_oarg_109_tvalid = dm_tvalid[109];
            assign m_axis_oarg_109_tkeep = dm_tkeep[109][M_AXIS_OARG_109_DMWIDTH/8-1:0];
            assign m_axis_oarg_109_tstrb = dm_tstrb[109][M_AXIS_OARG_109_DMWIDTH/8-1:0];
            assign m_axis_oarg_109_tdata = dm_tdata[109][M_AXIS_OARG_109_DMWIDTH-1:0];
            assign ap_axis_oarg_109_tready = ap_tready[109];
            assign ap_tlast[109] = ap_axis_oarg_109_tlast;
            assign ap_tvalid[109] = ap_axis_oarg_109_tvalid;
            assign ap_tdata[109][M_AXIS_OARG_109_WIDTH-1:0] = ap_axis_oarg_109_tdata;
            assign ap_tkeep[109] = {M_AXIS_OARG_109_WIDTH/8{1'b1}};
            assign ap_tstrb[109] = {M_AXIS_OARG_109_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 110) begin
            assign axis_clk[110] = m_axis_oarg_110_aclk;
            assign axis_rst[110] = m_axis_oarg_110_aresetn;
            assign dm_tready[110] = m_axis_oarg_110_tready;
            assign m_axis_oarg_110_tlast = dm_tlast[110];
            assign m_axis_oarg_110_tvalid = dm_tvalid[110];
            assign m_axis_oarg_110_tkeep = dm_tkeep[110][M_AXIS_OARG_110_DMWIDTH/8-1:0];
            assign m_axis_oarg_110_tstrb = dm_tstrb[110][M_AXIS_OARG_110_DMWIDTH/8-1:0];
            assign m_axis_oarg_110_tdata = dm_tdata[110][M_AXIS_OARG_110_DMWIDTH-1:0];
            assign ap_axis_oarg_110_tready = ap_tready[110];
            assign ap_tlast[110] = ap_axis_oarg_110_tlast;
            assign ap_tvalid[110] = ap_axis_oarg_110_tvalid;
            assign ap_tdata[110][M_AXIS_OARG_110_WIDTH-1:0] = ap_axis_oarg_110_tdata;
            assign ap_tkeep[110] = {M_AXIS_OARG_110_WIDTH/8{1'b1}};
            assign ap_tstrb[110] = {M_AXIS_OARG_110_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 111) begin
            assign axis_clk[111] = m_axis_oarg_111_aclk;
            assign axis_rst[111] = m_axis_oarg_111_aresetn;
            assign dm_tready[111] = m_axis_oarg_111_tready;
            assign m_axis_oarg_111_tlast = dm_tlast[111];
            assign m_axis_oarg_111_tvalid = dm_tvalid[111];
            assign m_axis_oarg_111_tkeep = dm_tkeep[111][M_AXIS_OARG_111_DMWIDTH/8-1:0];
            assign m_axis_oarg_111_tstrb = dm_tstrb[111][M_AXIS_OARG_111_DMWIDTH/8-1:0];
            assign m_axis_oarg_111_tdata = dm_tdata[111][M_AXIS_OARG_111_DMWIDTH-1:0];
            assign ap_axis_oarg_111_tready = ap_tready[111];
            assign ap_tlast[111] = ap_axis_oarg_111_tlast;
            assign ap_tvalid[111] = ap_axis_oarg_111_tvalid;
            assign ap_tdata[111][M_AXIS_OARG_111_WIDTH-1:0] = ap_axis_oarg_111_tdata;
            assign ap_tkeep[111] = {M_AXIS_OARG_111_WIDTH/8{1'b1}};
            assign ap_tstrb[111] = {M_AXIS_OARG_111_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 112) begin
            assign axis_clk[112] = m_axis_oarg_112_aclk;
            assign axis_rst[112] = m_axis_oarg_112_aresetn;
            assign dm_tready[112] = m_axis_oarg_112_tready;
            assign m_axis_oarg_112_tlast = dm_tlast[112];
            assign m_axis_oarg_112_tvalid = dm_tvalid[112];
            assign m_axis_oarg_112_tkeep = dm_tkeep[112][M_AXIS_OARG_112_DMWIDTH/8-1:0];
            assign m_axis_oarg_112_tstrb = dm_tstrb[112][M_AXIS_OARG_112_DMWIDTH/8-1:0];
            assign m_axis_oarg_112_tdata = dm_tdata[112][M_AXIS_OARG_112_DMWIDTH-1:0];
            assign ap_axis_oarg_112_tready = ap_tready[112];
            assign ap_tlast[112] = ap_axis_oarg_112_tlast;
            assign ap_tvalid[112] = ap_axis_oarg_112_tvalid;
            assign ap_tdata[112][M_AXIS_OARG_112_WIDTH-1:0] = ap_axis_oarg_112_tdata;
            assign ap_tkeep[112] = {M_AXIS_OARG_112_WIDTH/8{1'b1}};
            assign ap_tstrb[112] = {M_AXIS_OARG_112_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 113) begin
            assign axis_clk[113] = m_axis_oarg_113_aclk;
            assign axis_rst[113] = m_axis_oarg_113_aresetn;
            assign dm_tready[113] = m_axis_oarg_113_tready;
            assign m_axis_oarg_113_tlast = dm_tlast[113];
            assign m_axis_oarg_113_tvalid = dm_tvalid[113];
            assign m_axis_oarg_113_tkeep = dm_tkeep[113][M_AXIS_OARG_113_DMWIDTH/8-1:0];
            assign m_axis_oarg_113_tstrb = dm_tstrb[113][M_AXIS_OARG_113_DMWIDTH/8-1:0];
            assign m_axis_oarg_113_tdata = dm_tdata[113][M_AXIS_OARG_113_DMWIDTH-1:0];
            assign ap_axis_oarg_113_tready = ap_tready[113];
            assign ap_tlast[113] = ap_axis_oarg_113_tlast;
            assign ap_tvalid[113] = ap_axis_oarg_113_tvalid;
            assign ap_tdata[113][M_AXIS_OARG_113_WIDTH-1:0] = ap_axis_oarg_113_tdata;
            assign ap_tkeep[113] = {M_AXIS_OARG_113_WIDTH/8{1'b1}};
            assign ap_tstrb[113] = {M_AXIS_OARG_113_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 114) begin
            assign axis_clk[114] = m_axis_oarg_114_aclk;
            assign axis_rst[114] = m_axis_oarg_114_aresetn;
            assign dm_tready[114] = m_axis_oarg_114_tready;
            assign m_axis_oarg_114_tlast = dm_tlast[114];
            assign m_axis_oarg_114_tvalid = dm_tvalid[114];
            assign m_axis_oarg_114_tkeep = dm_tkeep[114][M_AXIS_OARG_114_DMWIDTH/8-1:0];
            assign m_axis_oarg_114_tstrb = dm_tstrb[114][M_AXIS_OARG_114_DMWIDTH/8-1:0];
            assign m_axis_oarg_114_tdata = dm_tdata[114][M_AXIS_OARG_114_DMWIDTH-1:0];
            assign ap_axis_oarg_114_tready = ap_tready[114];
            assign ap_tlast[114] = ap_axis_oarg_114_tlast;
            assign ap_tvalid[114] = ap_axis_oarg_114_tvalid;
            assign ap_tdata[114][M_AXIS_OARG_114_WIDTH-1:0] = ap_axis_oarg_114_tdata;
            assign ap_tkeep[114] = {M_AXIS_OARG_114_WIDTH/8{1'b1}};
            assign ap_tstrb[114] = {M_AXIS_OARG_114_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 115) begin
            assign axis_clk[115] = m_axis_oarg_115_aclk;
            assign axis_rst[115] = m_axis_oarg_115_aresetn;
            assign dm_tready[115] = m_axis_oarg_115_tready;
            assign m_axis_oarg_115_tlast = dm_tlast[115];
            assign m_axis_oarg_115_tvalid = dm_tvalid[115];
            assign m_axis_oarg_115_tkeep = dm_tkeep[115][M_AXIS_OARG_115_DMWIDTH/8-1:0];
            assign m_axis_oarg_115_tstrb = dm_tstrb[115][M_AXIS_OARG_115_DMWIDTH/8-1:0];
            assign m_axis_oarg_115_tdata = dm_tdata[115][M_AXIS_OARG_115_DMWIDTH-1:0];
            assign ap_axis_oarg_115_tready = ap_tready[115];
            assign ap_tlast[115] = ap_axis_oarg_115_tlast;
            assign ap_tvalid[115] = ap_axis_oarg_115_tvalid;
            assign ap_tdata[115][M_AXIS_OARG_115_WIDTH-1:0] = ap_axis_oarg_115_tdata;
            assign ap_tkeep[115] = {M_AXIS_OARG_115_WIDTH/8{1'b1}};
            assign ap_tstrb[115] = {M_AXIS_OARG_115_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 116) begin
            assign axis_clk[116] = m_axis_oarg_116_aclk;
            assign axis_rst[116] = m_axis_oarg_116_aresetn;
            assign dm_tready[116] = m_axis_oarg_116_tready;
            assign m_axis_oarg_116_tlast = dm_tlast[116];
            assign m_axis_oarg_116_tvalid = dm_tvalid[116];
            assign m_axis_oarg_116_tkeep = dm_tkeep[116][M_AXIS_OARG_116_DMWIDTH/8-1:0];
            assign m_axis_oarg_116_tstrb = dm_tstrb[116][M_AXIS_OARG_116_DMWIDTH/8-1:0];
            assign m_axis_oarg_116_tdata = dm_tdata[116][M_AXIS_OARG_116_DMWIDTH-1:0];
            assign ap_axis_oarg_116_tready = ap_tready[116];
            assign ap_tlast[116] = ap_axis_oarg_116_tlast;
            assign ap_tvalid[116] = ap_axis_oarg_116_tvalid;
            assign ap_tdata[116][M_AXIS_OARG_116_WIDTH-1:0] = ap_axis_oarg_116_tdata;
            assign ap_tkeep[116] = {M_AXIS_OARG_116_WIDTH/8{1'b1}};
            assign ap_tstrb[116] = {M_AXIS_OARG_116_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 117) begin
            assign axis_clk[117] = m_axis_oarg_117_aclk;
            assign axis_rst[117] = m_axis_oarg_117_aresetn;
            assign dm_tready[117] = m_axis_oarg_117_tready;
            assign m_axis_oarg_117_tlast = dm_tlast[117];
            assign m_axis_oarg_117_tvalid = dm_tvalid[117];
            assign m_axis_oarg_117_tkeep = dm_tkeep[117][M_AXIS_OARG_117_DMWIDTH/8-1:0];
            assign m_axis_oarg_117_tstrb = dm_tstrb[117][M_AXIS_OARG_117_DMWIDTH/8-1:0];
            assign m_axis_oarg_117_tdata = dm_tdata[117][M_AXIS_OARG_117_DMWIDTH-1:0];
            assign ap_axis_oarg_117_tready = ap_tready[117];
            assign ap_tlast[117] = ap_axis_oarg_117_tlast;
            assign ap_tvalid[117] = ap_axis_oarg_117_tvalid;
            assign ap_tdata[117][M_AXIS_OARG_117_WIDTH-1:0] = ap_axis_oarg_117_tdata;
            assign ap_tkeep[117] = {M_AXIS_OARG_117_WIDTH/8{1'b1}};
            assign ap_tstrb[117] = {M_AXIS_OARG_117_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 118) begin
            assign axis_clk[118] = m_axis_oarg_118_aclk;
            assign axis_rst[118] = m_axis_oarg_118_aresetn;
            assign dm_tready[118] = m_axis_oarg_118_tready;
            assign m_axis_oarg_118_tlast = dm_tlast[118];
            assign m_axis_oarg_118_tvalid = dm_tvalid[118];
            assign m_axis_oarg_118_tkeep = dm_tkeep[118][M_AXIS_OARG_118_DMWIDTH/8-1:0];
            assign m_axis_oarg_118_tstrb = dm_tstrb[118][M_AXIS_OARG_118_DMWIDTH/8-1:0];
            assign m_axis_oarg_118_tdata = dm_tdata[118][M_AXIS_OARG_118_DMWIDTH-1:0];
            assign ap_axis_oarg_118_tready = ap_tready[118];
            assign ap_tlast[118] = ap_axis_oarg_118_tlast;
            assign ap_tvalid[118] = ap_axis_oarg_118_tvalid;
            assign ap_tdata[118][M_AXIS_OARG_118_WIDTH-1:0] = ap_axis_oarg_118_tdata;
            assign ap_tkeep[118] = {M_AXIS_OARG_118_WIDTH/8{1'b1}};
            assign ap_tstrb[118] = {M_AXIS_OARG_118_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 119) begin
            assign axis_clk[119] = m_axis_oarg_119_aclk;
            assign axis_rst[119] = m_axis_oarg_119_aresetn;
            assign dm_tready[119] = m_axis_oarg_119_tready;
            assign m_axis_oarg_119_tlast = dm_tlast[119];
            assign m_axis_oarg_119_tvalid = dm_tvalid[119];
            assign m_axis_oarg_119_tkeep = dm_tkeep[119][M_AXIS_OARG_119_DMWIDTH/8-1:0];
            assign m_axis_oarg_119_tstrb = dm_tstrb[119][M_AXIS_OARG_119_DMWIDTH/8-1:0];
            assign m_axis_oarg_119_tdata = dm_tdata[119][M_AXIS_OARG_119_DMWIDTH-1:0];
            assign ap_axis_oarg_119_tready = ap_tready[119];
            assign ap_tlast[119] = ap_axis_oarg_119_tlast;
            assign ap_tvalid[119] = ap_axis_oarg_119_tvalid;
            assign ap_tdata[119][M_AXIS_OARG_119_WIDTH-1:0] = ap_axis_oarg_119_tdata;
            assign ap_tkeep[119] = {M_AXIS_OARG_119_WIDTH/8{1'b1}};
            assign ap_tstrb[119] = {M_AXIS_OARG_119_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 120) begin
            assign axis_clk[120] = m_axis_oarg_120_aclk;
            assign axis_rst[120] = m_axis_oarg_120_aresetn;
            assign dm_tready[120] = m_axis_oarg_120_tready;
            assign m_axis_oarg_120_tlast = dm_tlast[120];
            assign m_axis_oarg_120_tvalid = dm_tvalid[120];
            assign m_axis_oarg_120_tkeep = dm_tkeep[120][M_AXIS_OARG_120_DMWIDTH/8-1:0];
            assign m_axis_oarg_120_tstrb = dm_tstrb[120][M_AXIS_OARG_120_DMWIDTH/8-1:0];
            assign m_axis_oarg_120_tdata = dm_tdata[120][M_AXIS_OARG_120_DMWIDTH-1:0];
            assign ap_axis_oarg_120_tready = ap_tready[120];
            assign ap_tlast[120] = ap_axis_oarg_120_tlast;
            assign ap_tvalid[120] = ap_axis_oarg_120_tvalid;
            assign ap_tdata[120][M_AXIS_OARG_120_WIDTH-1:0] = ap_axis_oarg_120_tdata;
            assign ap_tkeep[120] = {M_AXIS_OARG_120_WIDTH/8{1'b1}};
            assign ap_tstrb[120] = {M_AXIS_OARG_120_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 121) begin
            assign axis_clk[121] = m_axis_oarg_121_aclk;
            assign axis_rst[121] = m_axis_oarg_121_aresetn;
            assign dm_tready[121] = m_axis_oarg_121_tready;
            assign m_axis_oarg_121_tlast = dm_tlast[121];
            assign m_axis_oarg_121_tvalid = dm_tvalid[121];
            assign m_axis_oarg_121_tkeep = dm_tkeep[121][M_AXIS_OARG_121_DMWIDTH/8-1:0];
            assign m_axis_oarg_121_tstrb = dm_tstrb[121][M_AXIS_OARG_121_DMWIDTH/8-1:0];
            assign m_axis_oarg_121_tdata = dm_tdata[121][M_AXIS_OARG_121_DMWIDTH-1:0];
            assign ap_axis_oarg_121_tready = ap_tready[121];
            assign ap_tlast[121] = ap_axis_oarg_121_tlast;
            assign ap_tvalid[121] = ap_axis_oarg_121_tvalid;
            assign ap_tdata[121][M_AXIS_OARG_121_WIDTH-1:0] = ap_axis_oarg_121_tdata;
            assign ap_tkeep[121] = {M_AXIS_OARG_121_WIDTH/8{1'b1}};
            assign ap_tstrb[121] = {M_AXIS_OARG_121_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 122) begin
            assign axis_clk[122] = m_axis_oarg_122_aclk;
            assign axis_rst[122] = m_axis_oarg_122_aresetn;
            assign dm_tready[122] = m_axis_oarg_122_tready;
            assign m_axis_oarg_122_tlast = dm_tlast[122];
            assign m_axis_oarg_122_tvalid = dm_tvalid[122];
            assign m_axis_oarg_122_tkeep = dm_tkeep[122][M_AXIS_OARG_122_DMWIDTH/8-1:0];
            assign m_axis_oarg_122_tstrb = dm_tstrb[122][M_AXIS_OARG_122_DMWIDTH/8-1:0];
            assign m_axis_oarg_122_tdata = dm_tdata[122][M_AXIS_OARG_122_DMWIDTH-1:0];
            assign ap_axis_oarg_122_tready = ap_tready[122];
            assign ap_tlast[122] = ap_axis_oarg_122_tlast;
            assign ap_tvalid[122] = ap_axis_oarg_122_tvalid;
            assign ap_tdata[122][M_AXIS_OARG_122_WIDTH-1:0] = ap_axis_oarg_122_tdata;
            assign ap_tkeep[122] = {M_AXIS_OARG_122_WIDTH/8{1'b1}};
            assign ap_tstrb[122] = {M_AXIS_OARG_122_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 123) begin
            assign axis_clk[123] = m_axis_oarg_123_aclk;
            assign axis_rst[123] = m_axis_oarg_123_aresetn;
            assign dm_tready[123] = m_axis_oarg_123_tready;
            assign m_axis_oarg_123_tlast = dm_tlast[123];
            assign m_axis_oarg_123_tvalid = dm_tvalid[123];
            assign m_axis_oarg_123_tkeep = dm_tkeep[123][M_AXIS_OARG_123_DMWIDTH/8-1:0];
            assign m_axis_oarg_123_tstrb = dm_tstrb[123][M_AXIS_OARG_123_DMWIDTH/8-1:0];
            assign m_axis_oarg_123_tdata = dm_tdata[123][M_AXIS_OARG_123_DMWIDTH-1:0];
            assign ap_axis_oarg_123_tready = ap_tready[123];
            assign ap_tlast[123] = ap_axis_oarg_123_tlast;
            assign ap_tvalid[123] = ap_axis_oarg_123_tvalid;
            assign ap_tdata[123][M_AXIS_OARG_123_WIDTH-1:0] = ap_axis_oarg_123_tdata;
            assign ap_tkeep[123] = {M_AXIS_OARG_123_WIDTH/8{1'b1}};
            assign ap_tstrb[123] = {M_AXIS_OARG_123_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 124) begin
            assign axis_clk[124] = m_axis_oarg_124_aclk;
            assign axis_rst[124] = m_axis_oarg_124_aresetn;
            assign dm_tready[124] = m_axis_oarg_124_tready;
            assign m_axis_oarg_124_tlast = dm_tlast[124];
            assign m_axis_oarg_124_tvalid = dm_tvalid[124];
            assign m_axis_oarg_124_tkeep = dm_tkeep[124][M_AXIS_OARG_124_DMWIDTH/8-1:0];
            assign m_axis_oarg_124_tstrb = dm_tstrb[124][M_AXIS_OARG_124_DMWIDTH/8-1:0];
            assign m_axis_oarg_124_tdata = dm_tdata[124][M_AXIS_OARG_124_DMWIDTH-1:0];
            assign ap_axis_oarg_124_tready = ap_tready[124];
            assign ap_tlast[124] = ap_axis_oarg_124_tlast;
            assign ap_tvalid[124] = ap_axis_oarg_124_tvalid;
            assign ap_tdata[124][M_AXIS_OARG_124_WIDTH-1:0] = ap_axis_oarg_124_tdata;
            assign ap_tkeep[124] = {M_AXIS_OARG_124_WIDTH/8{1'b1}};
            assign ap_tstrb[124] = {M_AXIS_OARG_124_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 125) begin
            assign axis_clk[125] = m_axis_oarg_125_aclk;
            assign axis_rst[125] = m_axis_oarg_125_aresetn;
            assign dm_tready[125] = m_axis_oarg_125_tready;
            assign m_axis_oarg_125_tlast = dm_tlast[125];
            assign m_axis_oarg_125_tvalid = dm_tvalid[125];
            assign m_axis_oarg_125_tkeep = dm_tkeep[125][M_AXIS_OARG_125_DMWIDTH/8-1:0];
            assign m_axis_oarg_125_tstrb = dm_tstrb[125][M_AXIS_OARG_125_DMWIDTH/8-1:0];
            assign m_axis_oarg_125_tdata = dm_tdata[125][M_AXIS_OARG_125_DMWIDTH-1:0];
            assign ap_axis_oarg_125_tready = ap_tready[125];
            assign ap_tlast[125] = ap_axis_oarg_125_tlast;
            assign ap_tvalid[125] = ap_axis_oarg_125_tvalid;
            assign ap_tdata[125][M_AXIS_OARG_125_WIDTH-1:0] = ap_axis_oarg_125_tdata;
            assign ap_tkeep[125] = {M_AXIS_OARG_125_WIDTH/8{1'b1}};
            assign ap_tstrb[125] = {M_AXIS_OARG_125_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 126) begin
            assign axis_clk[126] = m_axis_oarg_126_aclk;
            assign axis_rst[126] = m_axis_oarg_126_aresetn;
            assign dm_tready[126] = m_axis_oarg_126_tready;
            assign m_axis_oarg_126_tlast = dm_tlast[126];
            assign m_axis_oarg_126_tvalid = dm_tvalid[126];
            assign m_axis_oarg_126_tkeep = dm_tkeep[126][M_AXIS_OARG_126_DMWIDTH/8-1:0];
            assign m_axis_oarg_126_tstrb = dm_tstrb[126][M_AXIS_OARG_126_DMWIDTH/8-1:0];
            assign m_axis_oarg_126_tdata = dm_tdata[126][M_AXIS_OARG_126_DMWIDTH-1:0];
            assign ap_axis_oarg_126_tready = ap_tready[126];
            assign ap_tlast[126] = ap_axis_oarg_126_tlast;
            assign ap_tvalid[126] = ap_axis_oarg_126_tvalid;
            assign ap_tdata[126][M_AXIS_OARG_126_WIDTH-1:0] = ap_axis_oarg_126_tdata;
            assign ap_tkeep[126] = {M_AXIS_OARG_126_WIDTH/8{1'b1}};
            assign ap_tstrb[126] = {M_AXIS_OARG_126_WIDTH/8{1'b1}};
        end
        if(C_NUM_OUTPUT_AXISs > 127) begin
            assign axis_clk[127] = m_axis_oarg_127_aclk;
            assign axis_rst[127] = m_axis_oarg_127_aresetn;
            assign dm_tready[127] = m_axis_oarg_127_tready;
            assign m_axis_oarg_127_tlast = dm_tlast[127];
            assign m_axis_oarg_127_tvalid = dm_tvalid[127];
            assign m_axis_oarg_127_tkeep = dm_tkeep[127][M_AXIS_OARG_127_DMWIDTH/8-1:0];
            assign m_axis_oarg_127_tstrb = dm_tstrb[127][M_AXIS_OARG_127_DMWIDTH/8-1:0];
            assign m_axis_oarg_127_tdata = dm_tdata[127][M_AXIS_OARG_127_DMWIDTH-1:0];
            assign ap_axis_oarg_127_tready = ap_tready[127];
            assign ap_tlast[127] = ap_axis_oarg_127_tlast;
            assign ap_tvalid[127] = ap_axis_oarg_127_tvalid;
            assign ap_tdata[127][M_AXIS_OARG_127_WIDTH-1:0] = ap_axis_oarg_127_tdata;
            assign ap_tkeep[127] = {M_AXIS_OARG_127_WIDTH/8{1'b1}};
            assign ap_tstrb[127] = {M_AXIS_OARG_127_WIDTH/8{1'b1}};
        end
    endgenerate    
    
    //instantiate the axis2axis modules
    genvar idx;
    generate
        for(idx=0; idx<C_NUM_OUTPUT_AXISs; idx=idx+1) begin: OUT_AXIS_GEN
            outaxis #( 
                .DATA_WIDTH(C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                .GEN_TLAST(C_GEN_TLAST_BIT_ARRAY[32*(idx+1)-1:32*idx])
            ) outaxis_i (
                .ACC_CLK(acc_clk),
                .ARESETN(acc_aresetn),
                .CTRL_ALLOW(out_axis_allow),
                .CTRL_READY(out_axis_ready[idx]),
                .CTRL_FINISHED(out_axis_finished[idx]),
                .DM_TLAST(buf_tlast[idx]),
                .DM_TVALID(buf_tvalid[idx]),
                .DM_TDATA(buf_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .DM_TREADY(buf_tready[idx]),
                .AP_TLAST(ap_tlast[idx]),
                .AP_TVALID(ap_tvalid[idx]),
                .AP_TDATA(ap_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .AP_TREADY(ap_tready[idx])
            );
            
            if(C_DEPTH_BIT_ARRAY[32*(idx+1)-1:32*idx] > 0) begin
                //use fifo
                axis_fifo #(
                    .C_DATA_WIDTH(C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_DATA_DEPTH(C_DEPTH_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_IS_ASYNC(C_IS_ASYNC_BIT_ARRAY[32*(idx+1)-1:32*idx])
                ) axis_fifo_i (
                    .aresetn(acc_aresetn),
                    .inclk(acc_clk),
                    .in_tdata(buf_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .in_tlast(buf_tlast[idx]),  
                    .in_tvalid(buf_tvalid[idx]),
                    .in_tready(buf_tready[idx]),
                    .outclk(axis_clk[idx]), 
                    .out_tdata(dwconv_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .out_tready(dwconv_tready[idx]),
                    .out_tvalid(dwconv_tvalid[idx]),
                    .out_tlast(dwconv_tlast[idx])
                );
            end
            else begin
                //if not, wire the input signals straight through
                assign dwconv_tlast[idx] = buf_tlast[idx];
                assign dwconv_tvalid[idx] = buf_tvalid[idx];
                assign buf_tready[idx] = dwconv_tready[idx];   //output
                assign dwconv_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = buf_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            end
            
            //check if data width converter is needed
            if(C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx] != C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]) begin
                 axis_dwidth_converter_v1_1_9_axis_dwidth_converter #(
                    .C_S_AXIS_TDATA_WIDTH(C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_M_AXIS_TDATA_WIDTH(C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_AXIS_TID_WIDTH(1),
                    .C_AXIS_TDEST_WIDTH(1),
                    .C_S_AXIS_TUSER_WIDTH(1),
                    .C_M_AXIS_TUSER_WIDTH(1),
                    .C_AXIS_SIGNAL_SET(32'h1F)  //Enabled: TLAST, TKEEP, TSTRB, TDATA, TREADY
                ) data_width_conv_i (
                    .aclk(axis_clk[idx]),
                    .aresetn(axis_rst[idx]),
                    .aclken(1'b1),
                    .s_axis_tvalid(dwconv_tvalid[idx]),
                    .s_axis_tready(dwconv_tready[idx]),
                    .s_axis_tdata(dwconv_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .s_axis_tstrb(ap_tstrb[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tkeep(ap_tkeep[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tlast(dwconv_tlast[idx]),
//                    .s_axis_tid(),
//                    .s_axis_tdest(),
//                    .s_axis_tuser(),
                    .m_axis_tvalid(dm_tvalid[idx]),
                    .m_axis_tready(dm_tready[idx]),
                    .m_axis_tdata(dm_tdata[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .m_axis_tstrb(dm_tstrb[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .m_axis_tkeep(dm_tkeep[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .m_axis_tlast(dm_tlast[idx])
//                    .m_axis_tid(),
//                    .m_axis_tdest(),
//                    .m_axis_tuser()
                );
            end
            else begin
                //if no data width converter, wire the input signals straight through
                assign dm_tlast[idx] = dwconv_tlast[idx];
                assign dm_tvalid[idx] = dwconv_tvalid[idx];
                assign dwconv_tready[idx] = dm_tready[idx];   //output
                assign dm_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = dwconv_tdata[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
                assign dm_tstrb[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0] = ap_tstrb[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0];
                assign dm_tkeep[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0] = ap_tkeep[idx][C_OUTAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0];
            end
        end
    endgenerate
endmodule
