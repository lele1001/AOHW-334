// (c) Copyright 2022, Advanced Micro Devices, Inc.
// 
// Permission is hereby granted, free of charge, to any person obtaining a 
// copy of this software and associated documentation files (the "Software"), 
// to deal in the Software without restriction, including without limitation 
// the rights to use, copy, modify, merge, publish, distribute, sublicense, 
// and/or sell copies of the Software, and to permit persons to whom the 
// Software is furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in 
// all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR 
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL 
// THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER 
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
// FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER 
// DEALINGS IN THE SOFTWARE.
//--------------------------------------------------------------------------

`timescale 1ps/1ps

module hw_discovery #(
   parameter integer C_NUM_PFS                     		     = 1,
   parameter [11:0]  C_CAP_BASE_ADDR               		     = 12'h600,
   parameter [11:0]  C_NEXT_CAP_ADDR           		         = 12'h0,
   parameter integer C_PF0_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter integer C_PF0_HAS_UUID_ROM	                   = 0,
   parameter integer C_PF0_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF0_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF0_HIGH_OFFSET             		     = 32'h0,
   parameter         C_PF0_UUID_ROM_INIT                   = "0",
   parameter [7:0]   C_PF0_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_13                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_14                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_14                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_14                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_14          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_14          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_14           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_14                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_15                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_15                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_15                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_15          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_15          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_15           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_15                  = 4'h0,
   parameter integer C_PF0_S_AXI_DATA_WIDTH                = 32,
   parameter integer C_PF0_S_AXI_ADDR_WIDTH                = 32,
   parameter integer C_PF1_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter         C_PF1_HAS_UUID_ROM	                   = 0,
   parameter integer C_PF1_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF1_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF1_HIGH_OFFSET             		     = 32'h0,
   parameter         C_PF1_UUID_ROM_INIT                   = "0",
   parameter [7:0]   C_PF1_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_13                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_14                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_14                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_14                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_14          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_14          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_14           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_14                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_15                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_15                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_15                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_15          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_15          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_15           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_15                  = 4'h0,
   parameter integer C_PF1_S_AXI_DATA_WIDTH                = 32,
   parameter integer C_PF1_S_AXI_ADDR_WIDTH                = 32,   
   parameter integer C_PF2_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter         C_PF2_HAS_UUID_ROM	                   = 0,
   parameter integer C_PF2_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF2_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF2_HIGH_OFFSET             		     = 32'h0,
   parameter         C_PF2_UUID_ROM_INIT                   = "0",
   parameter [7:0]   C_PF2_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_13                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_14                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_14                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_14                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_14          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_14          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_14           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_14                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_15                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_15                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_15                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_15          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_15          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_15           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_15                  = 4'h0,
   parameter integer C_PF2_S_AXI_DATA_WIDTH                = 32,
   parameter integer C_PF2_S_AXI_ADDR_WIDTH                = 32,   
   parameter integer C_PF3_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter         C_PF3_HAS_UUID_ROM	                   = 0,
   parameter integer C_PF3_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF3_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF3_HIGH_OFFSET             		     = 32'h0,
   parameter         C_PF3_UUID_ROM_INIT                   = "0",
   parameter [7:0]   C_PF3_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_13                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_14                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_14                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_14                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_14          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_14          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_14           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_14                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_15                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_15                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_15                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_15          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_15          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_15           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_15                  = 4'h0,
   parameter integer C_PF3_S_AXI_DATA_WIDTH                = 32,
   parameter integer C_PF3_S_AXI_ADDR_WIDTH                = 32,      
   parameter         C_XDEVICEFAMILY                       = "no_family" 
   )
  (
   // Clocks & Resets
   input wire                                    aclk_pcie,
   input wire                                    aresetn_pcie,
   input wire                                    aclk_ctrl,
   input wire                                    aresetn_ctrl,
   
   // slave pcie4_cfg_ext Interface (aclk_pcie)
   input  wire [7:0]                             s_pcie4_cfg_ext_function_number,
   output wire [31:0]                            s_pcie4_cfg_ext_read_data,
   output wire                                   s_pcie4_cfg_ext_read_data_valid,
   input  wire                                   s_pcie4_cfg_ext_read_received,
   input  wire [9:0]                             s_pcie4_cfg_ext_register_number,
   input  wire [3:0]                             s_pcie4_cfg_ext_write_byte_enable,
   input  wire [31:0]                            s_pcie4_cfg_ext_write_data,
   input  wire                                   s_pcie4_cfg_ext_write_received,
   
   // slave pcie4_cfg_ext Interface (aclk_pcie)
   output wire [7:0]                             m_pcie4_cfg_ext_function_number,
   input  wire [31:0]                            m_pcie4_cfg_ext_read_data,
   input  wire                                   m_pcie4_cfg_ext_read_data_valid,
   output wire                                   m_pcie4_cfg_ext_read_received,
   output wire [9:0]                             m_pcie4_cfg_ext_register_number,
   output wire [3:0]                             m_pcie4_cfg_ext_write_byte_enable,
   output wire [31:0]                            m_pcie4_cfg_ext_write_data,
   output wire                                   m_pcie4_cfg_ext_write_received,
   
   // AXI Interface (aclk_ctrl) for PF0
   input  wire [C_PF0_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf0_AWADDR,
   input  wire                                   s_axi_ctrl_pf0_AWVALID,
   output wire                                   s_axi_ctrl_pf0_AWREADY,
   input  wire [C_PF0_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf0_WDATA,
   input  wire [C_PF0_S_AXI_DATA_WIDTH/8-1:0]    s_axi_ctrl_pf0_WSTRB,
   input  wire                                   s_axi_ctrl_pf0_WVALID,
   output wire                                   s_axi_ctrl_pf0_WREADY,
   output wire [1:0]                             s_axi_ctrl_pf0_BRESP,
   output wire                                   s_axi_ctrl_pf0_BVALID,
   input  wire                                   s_axi_ctrl_pf0_BREADY,
   input  wire [C_PF0_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf0_ARADDR,
   input  wire                                   s_axi_ctrl_pf0_ARVALID,
   output wire                                   s_axi_ctrl_pf0_ARREADY,
   output wire [C_PF0_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf0_RDATA,
   output wire [1:0]                             s_axi_ctrl_pf0_RRESP,
   output wire                                   s_axi_ctrl_pf0_RVALID,
   input  wire                                   s_axi_ctrl_pf0_RREADY,
   
   // AXI Interface (aclk_ctrl) for PF1
   input  wire [C_PF1_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf1_AWADDR,
   input  wire                                   s_axi_ctrl_pf1_AWVALID,
   output wire                                   s_axi_ctrl_pf1_AWREADY,
   input  wire [C_PF1_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf1_WDATA,
   input  wire [C_PF1_S_AXI_DATA_WIDTH/8-1:0]    s_axi_ctrl_pf1_WSTRB,
   input  wire                                   s_axi_ctrl_pf1_WVALID,
   output wire                                   s_axi_ctrl_pf1_WREADY,
   output wire [1:0]                             s_axi_ctrl_pf1_BRESP,
   output wire                                   s_axi_ctrl_pf1_BVALID,
   input  wire                                   s_axi_ctrl_pf1_BREADY,
   input  wire [C_PF1_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf1_ARADDR,
   input  wire                                   s_axi_ctrl_pf1_ARVALID,
   output wire                                   s_axi_ctrl_pf1_ARREADY,
   output wire [C_PF1_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf1_RDATA,
   output wire [1:0]                             s_axi_ctrl_pf1_RRESP,
   output wire                                   s_axi_ctrl_pf1_RVALID,
   input  wire                                   s_axi_ctrl_pf1_RREADY,
   
   // AXI Interface (aclk_ctrl) for PF2
   input  wire [C_PF2_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf2_AWADDR,
   input  wire                                   s_axi_ctrl_pf2_AWVALID,
   output wire                                   s_axi_ctrl_pf2_AWREADY,
   input  wire [C_PF2_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf2_WDATA,
   input  wire [C_PF2_S_AXI_DATA_WIDTH/8-1:0]    s_axi_ctrl_pf2_WSTRB,
   input  wire                                   s_axi_ctrl_pf2_WVALID,
   output wire                                   s_axi_ctrl_pf2_WREADY,
   output wire [1:0]                             s_axi_ctrl_pf2_BRESP,
   output wire                                   s_axi_ctrl_pf2_BVALID,
   input  wire                                   s_axi_ctrl_pf2_BREADY,
   input  wire [C_PF2_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf2_ARADDR,
   input  wire                                   s_axi_ctrl_pf2_ARVALID,
   output wire                                   s_axi_ctrl_pf2_ARREADY,
   output wire [C_PF2_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf2_RDATA,
   output wire [1:0]                             s_axi_ctrl_pf2_RRESP,
   output wire                                   s_axi_ctrl_pf2_RVALID,
   input  wire                                   s_axi_ctrl_pf2_RREADY,
   
   // AXI Interface (aclk_ctrl) for PF3
   input  wire [C_PF3_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf3_AWADDR,
   input  wire                                   s_axi_ctrl_pf3_AWVALID,
   output wire                                   s_axi_ctrl_pf3_AWREADY,
   input  wire [C_PF3_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf3_WDATA,
   input  wire [C_PF3_S_AXI_DATA_WIDTH/8-1:0]    s_axi_ctrl_pf3_WSTRB,
   input  wire                                   s_axi_ctrl_pf3_WVALID,
   output wire                                   s_axi_ctrl_pf3_WREADY,
   output wire [1:0]                             s_axi_ctrl_pf3_BRESP,
   output wire                                   s_axi_ctrl_pf3_BVALID,
   input  wire                                   s_axi_ctrl_pf3_BREADY,
   input  wire [C_PF3_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf3_ARADDR,
   input  wire                                   s_axi_ctrl_pf3_ARVALID,
   output wire                                   s_axi_ctrl_pf3_ARREADY,
   output wire [C_PF3_S_AXI_DATA_WIDTH-1:0]      s_axi_ctrl_pf3_RDATA,
   output wire [1:0]                             s_axi_ctrl_pf3_RRESP,
   output wire                                   s_axi_ctrl_pf3_RVALID,
   input  wire                                   s_axi_ctrl_pf3_RREADY
  );
  
    hw_disc #(
			.C_NUM_PFS                     		    (C_NUM_PFS                     		 ),
			.C_CAP_BASE_ADDR               		    (C_CAP_BASE_ADDR               		 ),
			.C_NEXT_CAP_ADDR           		        (C_NEXT_CAP_ADDR           		     ),
			.C_PF0_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF0_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF0_HAS_UUID_ROM	                  (C_PF0_HAS_UUID_ROM	               ),
			.C_PF0_BAR_INDEX               		    (C_PF0_BAR_INDEX               		 ),
			.C_PF0_LOW_OFFSET              		    (C_PF0_LOW_OFFSET              		 ),
			.C_PF0_HIGH_OFFSET             		    (C_PF0_HIGH_OFFSET             		 ),
			.C_PF0_UUID_ROM_INIT                  (C_PF0_UUID_ROM_INIT               ),
			.C_PF0_ENTRY_TYPE_0                   (C_PF0_ENTRY_TYPE_0                ),
			.C_PF0_ENTRY_BAR_0                    (C_PF0_ENTRY_BAR_0                 ),
			.C_PF0_ENTRY_ADDR_0                   (C_PF0_ENTRY_ADDR_0                ),
			.C_PF0_ENTRY_MAJOR_VERSION_0          (C_PF0_ENTRY_MAJOR_VERSION_0       ),
			.C_PF0_ENTRY_MINOR_VERSION_0          (C_PF0_ENTRY_MINOR_VERSION_0       ),
			.C_PF0_ENTRY_VERSION_TYPE_0           (C_PF0_ENTRY_VERSION_TYPE_0        ),
			.C_PF0_ENTRY_RSVD0_0                  (C_PF0_ENTRY_RSVD0_0               ),
			.C_PF0_ENTRY_TYPE_1                   (C_PF0_ENTRY_TYPE_1                ),
			.C_PF0_ENTRY_BAR_1                    (C_PF0_ENTRY_BAR_1                 ),
			.C_PF0_ENTRY_ADDR_1                   (C_PF0_ENTRY_ADDR_1                ),
			.C_PF0_ENTRY_MAJOR_VERSION_1          (C_PF0_ENTRY_MAJOR_VERSION_1       ),
			.C_PF0_ENTRY_MINOR_VERSION_1          (C_PF0_ENTRY_MINOR_VERSION_1       ),
			.C_PF0_ENTRY_VERSION_TYPE_1           (C_PF0_ENTRY_VERSION_TYPE_1        ),
			.C_PF0_ENTRY_RSVD0_1                  (C_PF0_ENTRY_RSVD0_1               ),
			.C_PF0_ENTRY_TYPE_2                   (C_PF0_ENTRY_TYPE_2                ),
			.C_PF0_ENTRY_BAR_2                    (C_PF0_ENTRY_BAR_2                 ),
			.C_PF0_ENTRY_ADDR_2                   (C_PF0_ENTRY_ADDR_2                ),
			.C_PF0_ENTRY_MAJOR_VERSION_2          (C_PF0_ENTRY_MAJOR_VERSION_2       ),
			.C_PF0_ENTRY_MINOR_VERSION_2          (C_PF0_ENTRY_MINOR_VERSION_2       ),
			.C_PF0_ENTRY_VERSION_TYPE_2           (C_PF0_ENTRY_VERSION_TYPE_2        ),
			.C_PF0_ENTRY_RSVD0_2                  (C_PF0_ENTRY_RSVD0_2               ),
			.C_PF0_ENTRY_TYPE_3                   (C_PF0_ENTRY_TYPE_3                ),
			.C_PF0_ENTRY_BAR_3                    (C_PF0_ENTRY_BAR_3                 ),
			.C_PF0_ENTRY_ADDR_3                   (C_PF0_ENTRY_ADDR_3                ),
			.C_PF0_ENTRY_MAJOR_VERSION_3          (C_PF0_ENTRY_MAJOR_VERSION_3       ),
			.C_PF0_ENTRY_MINOR_VERSION_3          (C_PF0_ENTRY_MINOR_VERSION_3       ),
			.C_PF0_ENTRY_VERSION_TYPE_3           (C_PF0_ENTRY_VERSION_TYPE_3        ),
			.C_PF0_ENTRY_RSVD0_3                  (C_PF0_ENTRY_RSVD0_3               ),
			.C_PF0_ENTRY_TYPE_4                   (C_PF0_ENTRY_TYPE_4                ),
			.C_PF0_ENTRY_BAR_4                    (C_PF0_ENTRY_BAR_4                 ),
			.C_PF0_ENTRY_ADDR_4                   (C_PF0_ENTRY_ADDR_4                ),
			.C_PF0_ENTRY_MAJOR_VERSION_4          (C_PF0_ENTRY_MAJOR_VERSION_4       ),
			.C_PF0_ENTRY_MINOR_VERSION_4          (C_PF0_ENTRY_MINOR_VERSION_4       ),
			.C_PF0_ENTRY_VERSION_TYPE_4           (C_PF0_ENTRY_VERSION_TYPE_4        ),
			.C_PF0_ENTRY_RSVD0_4                  (C_PF0_ENTRY_RSVD0_4               ),
			.C_PF0_ENTRY_TYPE_5                   (C_PF0_ENTRY_TYPE_5                ),
			.C_PF0_ENTRY_BAR_5                    (C_PF0_ENTRY_BAR_5                 ),
			.C_PF0_ENTRY_ADDR_5                   (C_PF0_ENTRY_ADDR_5                ),
			.C_PF0_ENTRY_MAJOR_VERSION_5          (C_PF0_ENTRY_MAJOR_VERSION_5       ),
			.C_PF0_ENTRY_MINOR_VERSION_5          (C_PF0_ENTRY_MINOR_VERSION_5       ),
			.C_PF0_ENTRY_VERSION_TYPE_5           (C_PF0_ENTRY_VERSION_TYPE_5        ),
			.C_PF0_ENTRY_RSVD0_5                  (C_PF0_ENTRY_RSVD0_5               ),
			.C_PF0_ENTRY_TYPE_6                   (C_PF0_ENTRY_TYPE_6                ),
			.C_PF0_ENTRY_BAR_6                    (C_PF0_ENTRY_BAR_6                 ),
			.C_PF0_ENTRY_ADDR_6                   (C_PF0_ENTRY_ADDR_6                ),
			.C_PF0_ENTRY_MAJOR_VERSION_6          (C_PF0_ENTRY_MAJOR_VERSION_6       ),
			.C_PF0_ENTRY_MINOR_VERSION_6          (C_PF0_ENTRY_MINOR_VERSION_6       ),
			.C_PF0_ENTRY_VERSION_TYPE_6           (C_PF0_ENTRY_VERSION_TYPE_6        ),
			.C_PF0_ENTRY_RSVD0_6                  (C_PF0_ENTRY_RSVD0_6               ),
			.C_PF0_ENTRY_TYPE_7                   (C_PF0_ENTRY_TYPE_7                ),
			.C_PF0_ENTRY_BAR_7                    (C_PF0_ENTRY_BAR_7                 ),
			.C_PF0_ENTRY_ADDR_7                   (C_PF0_ENTRY_ADDR_7                ),
			.C_PF0_ENTRY_MAJOR_VERSION_7          (C_PF0_ENTRY_MAJOR_VERSION_7       ),
			.C_PF0_ENTRY_MINOR_VERSION_7          (C_PF0_ENTRY_MINOR_VERSION_7       ),
			.C_PF0_ENTRY_VERSION_TYPE_7           (C_PF0_ENTRY_VERSION_TYPE_7        ),
			.C_PF0_ENTRY_RSVD0_7                  (C_PF0_ENTRY_RSVD0_7               ),
			.C_PF0_ENTRY_TYPE_8                   (C_PF0_ENTRY_TYPE_8                ),
			.C_PF0_ENTRY_BAR_8                    (C_PF0_ENTRY_BAR_8                 ),
			.C_PF0_ENTRY_ADDR_8                   (C_PF0_ENTRY_ADDR_8                ),
			.C_PF0_ENTRY_MAJOR_VERSION_8          (C_PF0_ENTRY_MAJOR_VERSION_8       ),
			.C_PF0_ENTRY_MINOR_VERSION_8          (C_PF0_ENTRY_MINOR_VERSION_8       ),
			.C_PF0_ENTRY_VERSION_TYPE_8           (C_PF0_ENTRY_VERSION_TYPE_8        ),
			.C_PF0_ENTRY_RSVD0_8                  (C_PF0_ENTRY_RSVD0_8               ),
			.C_PF0_ENTRY_TYPE_9                   (C_PF0_ENTRY_TYPE_9                ),
			.C_PF0_ENTRY_BAR_9                    (C_PF0_ENTRY_BAR_9                 ),
			.C_PF0_ENTRY_ADDR_9                   (C_PF0_ENTRY_ADDR_9                ),
			.C_PF0_ENTRY_MAJOR_VERSION_9          (C_PF0_ENTRY_MAJOR_VERSION_9       ),
			.C_PF0_ENTRY_MINOR_VERSION_9          (C_PF0_ENTRY_MINOR_VERSION_9       ),
			.C_PF0_ENTRY_VERSION_TYPE_9           (C_PF0_ENTRY_VERSION_TYPE_9        ),
			.C_PF0_ENTRY_RSVD0_9                  (C_PF0_ENTRY_RSVD0_9               ),
			.C_PF0_ENTRY_TYPE_10                  (C_PF0_ENTRY_TYPE_10               ),
			.C_PF0_ENTRY_BAR_10                   (C_PF0_ENTRY_BAR_10                ),
			.C_PF0_ENTRY_ADDR_10                  (C_PF0_ENTRY_ADDR_10               ),
			.C_PF0_ENTRY_MAJOR_VERSION_10         (C_PF0_ENTRY_MAJOR_VERSION_10      ),
			.C_PF0_ENTRY_MINOR_VERSION_10         (C_PF0_ENTRY_MINOR_VERSION_10      ),
			.C_PF0_ENTRY_VERSION_TYPE_10          (C_PF0_ENTRY_VERSION_TYPE_10       ),
			.C_PF0_ENTRY_RSVD0_10                 (C_PF0_ENTRY_RSVD0_10              ),
			.C_PF0_ENTRY_TYPE_11                  (C_PF0_ENTRY_TYPE_11               ),
			.C_PF0_ENTRY_BAR_11                   (C_PF0_ENTRY_BAR_11                ),
			.C_PF0_ENTRY_ADDR_11                  (C_PF0_ENTRY_ADDR_11               ),
			.C_PF0_ENTRY_MAJOR_VERSION_11         (C_PF0_ENTRY_MAJOR_VERSION_11      ),
			.C_PF0_ENTRY_MINOR_VERSION_11         (C_PF0_ENTRY_MINOR_VERSION_11      ),
			.C_PF0_ENTRY_VERSION_TYPE_11          (C_PF0_ENTRY_VERSION_TYPE_11       ),
			.C_PF0_ENTRY_RSVD0_11                 (C_PF0_ENTRY_RSVD0_11              ),
			.C_PF0_ENTRY_TYPE_12                  (C_PF0_ENTRY_TYPE_12               ),
			.C_PF0_ENTRY_BAR_12                   (C_PF0_ENTRY_BAR_12                ),
			.C_PF0_ENTRY_ADDR_12                  (C_PF0_ENTRY_ADDR_12               ),
			.C_PF0_ENTRY_MAJOR_VERSION_12         (C_PF0_ENTRY_MAJOR_VERSION_12      ),
			.C_PF0_ENTRY_MINOR_VERSION_12         (C_PF0_ENTRY_MINOR_VERSION_12      ),
			.C_PF0_ENTRY_VERSION_TYPE_12          (C_PF0_ENTRY_VERSION_TYPE_12       ),
			.C_PF0_ENTRY_RSVD0_12                 (C_PF0_ENTRY_RSVD0_12              ),
			.C_PF0_ENTRY_TYPE_13                  (C_PF0_ENTRY_TYPE_13               ),
			.C_PF0_ENTRY_BAR_13                   (C_PF0_ENTRY_BAR_13                ),
			.C_PF0_ENTRY_ADDR_13                  (C_PF0_ENTRY_ADDR_13               ),
			.C_PF0_ENTRY_MAJOR_VERSION_13         (C_PF0_ENTRY_MAJOR_VERSION_13      ),
			.C_PF0_ENTRY_MINOR_VERSION_13         (C_PF0_ENTRY_MINOR_VERSION_13      ),
			.C_PF0_ENTRY_VERSION_TYPE_13          (C_PF0_ENTRY_VERSION_TYPE_13       ),
			.C_PF0_ENTRY_RSVD0_13                 (C_PF0_ENTRY_RSVD0_13              ),
			.C_PF0_ENTRY_TYPE_14                  (C_PF0_ENTRY_TYPE_14               ),
			.C_PF0_ENTRY_BAR_14                   (C_PF0_ENTRY_BAR_14                ),
			.C_PF0_ENTRY_ADDR_14                  (C_PF0_ENTRY_ADDR_14               ),
			.C_PF0_ENTRY_MAJOR_VERSION_14         (C_PF0_ENTRY_MAJOR_VERSION_14      ),
			.C_PF0_ENTRY_MINOR_VERSION_14         (C_PF0_ENTRY_MINOR_VERSION_14      ),
			.C_PF0_ENTRY_VERSION_TYPE_14          (C_PF0_ENTRY_VERSION_TYPE_14       ),
			.C_PF0_ENTRY_RSVD0_14                 (C_PF0_ENTRY_RSVD0_14              ),
			.C_PF0_ENTRY_TYPE_15                  (C_PF0_ENTRY_TYPE_15               ),
			.C_PF0_ENTRY_BAR_15                   (C_PF0_ENTRY_BAR_15                ),
			.C_PF0_ENTRY_ADDR_15                  (C_PF0_ENTRY_ADDR_15               ),
			.C_PF0_ENTRY_MAJOR_VERSION_15         (C_PF0_ENTRY_MAJOR_VERSION_15      ),
			.C_PF0_ENTRY_MINOR_VERSION_15         (C_PF0_ENTRY_MINOR_VERSION_15      ),
			.C_PF0_ENTRY_VERSION_TYPE_15          (C_PF0_ENTRY_VERSION_TYPE_15       ),
			.C_PF0_ENTRY_RSVD0_15                 (C_PF0_ENTRY_RSVD0_15              ),
			.C_PF0_S_AXI_DATA_WIDTH               (C_PF0_S_AXI_DATA_WIDTH            ),
			.C_PF0_S_AXI_ADDR_WIDTH               (C_PF0_S_AXI_ADDR_WIDTH            ),
			.C_PF1_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF1_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF1_HAS_UUID_ROM	                  (C_PF1_HAS_UUID_ROM	               ),
			.C_PF1_BAR_INDEX               		    (C_PF1_BAR_INDEX               		 ),
			.C_PF1_LOW_OFFSET              		    (C_PF1_LOW_OFFSET              		 ),
			.C_PF1_HIGH_OFFSET             		    (C_PF1_HIGH_OFFSET             		 ),
			.C_PF1_UUID_ROM_INIT                  (C_PF1_UUID_ROM_INIT               ),
			.C_PF1_ENTRY_TYPE_0                   (C_PF1_ENTRY_TYPE_0                ),
			.C_PF1_ENTRY_BAR_0                    (C_PF1_ENTRY_BAR_0                 ),
			.C_PF1_ENTRY_ADDR_0                   (C_PF1_ENTRY_ADDR_0                ),
			.C_PF1_ENTRY_MAJOR_VERSION_0          (C_PF1_ENTRY_MAJOR_VERSION_0       ),
			.C_PF1_ENTRY_MINOR_VERSION_0          (C_PF1_ENTRY_MINOR_VERSION_0       ),
			.C_PF1_ENTRY_VERSION_TYPE_0           (C_PF1_ENTRY_VERSION_TYPE_0        ),
			.C_PF1_ENTRY_RSVD0_0                  (C_PF1_ENTRY_RSVD0_0               ),
			.C_PF1_ENTRY_TYPE_1                   (C_PF1_ENTRY_TYPE_1                ),
			.C_PF1_ENTRY_BAR_1                    (C_PF1_ENTRY_BAR_1                 ),
			.C_PF1_ENTRY_ADDR_1                   (C_PF1_ENTRY_ADDR_1                ),
			.C_PF1_ENTRY_MAJOR_VERSION_1          (C_PF1_ENTRY_MAJOR_VERSION_1       ),
			.C_PF1_ENTRY_MINOR_VERSION_1          (C_PF1_ENTRY_MINOR_VERSION_1       ),
			.C_PF1_ENTRY_VERSION_TYPE_1           (C_PF1_ENTRY_VERSION_TYPE_1        ),
			.C_PF1_ENTRY_RSVD0_1                  (C_PF1_ENTRY_RSVD0_1               ),
			.C_PF1_ENTRY_TYPE_2                   (C_PF1_ENTRY_TYPE_2                ),
			.C_PF1_ENTRY_BAR_2                    (C_PF1_ENTRY_BAR_2                 ),
			.C_PF1_ENTRY_ADDR_2                   (C_PF1_ENTRY_ADDR_2                ),
			.C_PF1_ENTRY_MAJOR_VERSION_2          (C_PF1_ENTRY_MAJOR_VERSION_2       ),
			.C_PF1_ENTRY_MINOR_VERSION_2          (C_PF1_ENTRY_MINOR_VERSION_2       ),
			.C_PF1_ENTRY_VERSION_TYPE_2           (C_PF1_ENTRY_VERSION_TYPE_2        ),
			.C_PF1_ENTRY_RSVD0_2                  (C_PF1_ENTRY_RSVD0_2               ),
			.C_PF1_ENTRY_TYPE_3                   (C_PF1_ENTRY_TYPE_3                ),
			.C_PF1_ENTRY_BAR_3                    (C_PF1_ENTRY_BAR_3                 ),
			.C_PF1_ENTRY_ADDR_3                   (C_PF1_ENTRY_ADDR_3                ),
			.C_PF1_ENTRY_MAJOR_VERSION_3          (C_PF1_ENTRY_MAJOR_VERSION_3       ),
			.C_PF1_ENTRY_MINOR_VERSION_3          (C_PF1_ENTRY_MINOR_VERSION_3       ),
			.C_PF1_ENTRY_VERSION_TYPE_3           (C_PF1_ENTRY_VERSION_TYPE_3        ),
			.C_PF1_ENTRY_RSVD0_3                  (C_PF1_ENTRY_RSVD0_3               ),
			.C_PF1_ENTRY_TYPE_4                   (C_PF1_ENTRY_TYPE_4                ),
			.C_PF1_ENTRY_BAR_4                    (C_PF1_ENTRY_BAR_4                 ),
			.C_PF1_ENTRY_ADDR_4                   (C_PF1_ENTRY_ADDR_4                ),
			.C_PF1_ENTRY_MAJOR_VERSION_4          (C_PF1_ENTRY_MAJOR_VERSION_4       ),
			.C_PF1_ENTRY_MINOR_VERSION_4          (C_PF1_ENTRY_MINOR_VERSION_4       ),
			.C_PF1_ENTRY_VERSION_TYPE_4           (C_PF1_ENTRY_VERSION_TYPE_4        ),
			.C_PF1_ENTRY_RSVD0_4                  (C_PF1_ENTRY_RSVD0_4               ),
			.C_PF1_ENTRY_TYPE_5                   (C_PF1_ENTRY_TYPE_5                ),
			.C_PF1_ENTRY_BAR_5                    (C_PF1_ENTRY_BAR_5                 ),
			.C_PF1_ENTRY_ADDR_5                   (C_PF1_ENTRY_ADDR_5                ),
			.C_PF1_ENTRY_MAJOR_VERSION_5          (C_PF1_ENTRY_MAJOR_VERSION_5       ),
			.C_PF1_ENTRY_MINOR_VERSION_5          (C_PF1_ENTRY_MINOR_VERSION_5       ),
			.C_PF1_ENTRY_VERSION_TYPE_5           (C_PF1_ENTRY_VERSION_TYPE_5        ),
			.C_PF1_ENTRY_RSVD0_5                  (C_PF1_ENTRY_RSVD0_5               ),
			.C_PF1_ENTRY_TYPE_6                   (C_PF1_ENTRY_TYPE_6                ),
			.C_PF1_ENTRY_BAR_6                    (C_PF1_ENTRY_BAR_6                 ),
			.C_PF1_ENTRY_ADDR_6                   (C_PF1_ENTRY_ADDR_6                ),
			.C_PF1_ENTRY_MAJOR_VERSION_6          (C_PF1_ENTRY_MAJOR_VERSION_6       ),
			.C_PF1_ENTRY_MINOR_VERSION_6          (C_PF1_ENTRY_MINOR_VERSION_6       ),
			.C_PF1_ENTRY_VERSION_TYPE_6           (C_PF1_ENTRY_VERSION_TYPE_6        ),
			.C_PF1_ENTRY_RSVD0_6                  (C_PF1_ENTRY_RSVD0_6               ),
			.C_PF1_ENTRY_TYPE_7                   (C_PF1_ENTRY_TYPE_7                ),
			.C_PF1_ENTRY_BAR_7                    (C_PF1_ENTRY_BAR_7                 ),
			.C_PF1_ENTRY_ADDR_7                   (C_PF1_ENTRY_ADDR_7                ),
			.C_PF1_ENTRY_MAJOR_VERSION_7          (C_PF1_ENTRY_MAJOR_VERSION_7       ),
			.C_PF1_ENTRY_MINOR_VERSION_7          (C_PF1_ENTRY_MINOR_VERSION_7       ),
			.C_PF1_ENTRY_VERSION_TYPE_7           (C_PF1_ENTRY_VERSION_TYPE_7        ),
			.C_PF1_ENTRY_RSVD0_7                  (C_PF1_ENTRY_RSVD0_7               ),
			.C_PF1_ENTRY_TYPE_8                   (C_PF1_ENTRY_TYPE_8                ),
			.C_PF1_ENTRY_BAR_8                    (C_PF1_ENTRY_BAR_8                 ),
			.C_PF1_ENTRY_ADDR_8                   (C_PF1_ENTRY_ADDR_8                ),
			.C_PF1_ENTRY_MAJOR_VERSION_8          (C_PF1_ENTRY_MAJOR_VERSION_8       ),
			.C_PF1_ENTRY_MINOR_VERSION_8          (C_PF1_ENTRY_MINOR_VERSION_8       ),
			.C_PF1_ENTRY_VERSION_TYPE_8           (C_PF1_ENTRY_VERSION_TYPE_8        ),
			.C_PF1_ENTRY_RSVD0_8                  (C_PF1_ENTRY_RSVD0_8               ),
			.C_PF1_ENTRY_TYPE_9                   (C_PF1_ENTRY_TYPE_9                ),
			.C_PF1_ENTRY_BAR_9                    (C_PF1_ENTRY_BAR_9                 ),
			.C_PF1_ENTRY_ADDR_9                   (C_PF1_ENTRY_ADDR_9                ),
			.C_PF1_ENTRY_MAJOR_VERSION_9          (C_PF1_ENTRY_MAJOR_VERSION_9       ),
			.C_PF1_ENTRY_MINOR_VERSION_9          (C_PF1_ENTRY_MINOR_VERSION_9       ),
			.C_PF1_ENTRY_VERSION_TYPE_9           (C_PF1_ENTRY_VERSION_TYPE_9        ),
			.C_PF1_ENTRY_RSVD0_9                  (C_PF1_ENTRY_RSVD0_9               ),
			.C_PF1_ENTRY_TYPE_10                  (C_PF1_ENTRY_TYPE_10               ),
			.C_PF1_ENTRY_BAR_10                   (C_PF1_ENTRY_BAR_10                ),
			.C_PF1_ENTRY_ADDR_10                  (C_PF1_ENTRY_ADDR_10               ),
			.C_PF1_ENTRY_MAJOR_VERSION_10         (C_PF1_ENTRY_MAJOR_VERSION_10      ),
			.C_PF1_ENTRY_MINOR_VERSION_10         (C_PF1_ENTRY_MINOR_VERSION_10      ),
			.C_PF1_ENTRY_VERSION_TYPE_10          (C_PF1_ENTRY_VERSION_TYPE_10       ),
			.C_PF1_ENTRY_RSVD0_10                 (C_PF1_ENTRY_RSVD0_10              ),
			.C_PF1_ENTRY_TYPE_11                  (C_PF1_ENTRY_TYPE_11               ),
			.C_PF1_ENTRY_BAR_11                   (C_PF1_ENTRY_BAR_11                ),
			.C_PF1_ENTRY_ADDR_11                  (C_PF1_ENTRY_ADDR_11               ),
			.C_PF1_ENTRY_MAJOR_VERSION_11         (C_PF1_ENTRY_MAJOR_VERSION_11      ),
			.C_PF1_ENTRY_MINOR_VERSION_11         (C_PF1_ENTRY_MINOR_VERSION_11      ),
			.C_PF1_ENTRY_VERSION_TYPE_11          (C_PF1_ENTRY_VERSION_TYPE_11       ),
			.C_PF1_ENTRY_RSVD0_11                 (C_PF1_ENTRY_RSVD0_11              ),
			.C_PF1_ENTRY_TYPE_12                  (C_PF1_ENTRY_TYPE_12               ),
			.C_PF1_ENTRY_BAR_12                   (C_PF1_ENTRY_BAR_12                ),
			.C_PF1_ENTRY_ADDR_12                  (C_PF1_ENTRY_ADDR_12               ),
			.C_PF1_ENTRY_MAJOR_VERSION_12         (C_PF1_ENTRY_MAJOR_VERSION_12      ),
			.C_PF1_ENTRY_MINOR_VERSION_12         (C_PF1_ENTRY_MINOR_VERSION_12      ),
			.C_PF1_ENTRY_VERSION_TYPE_12          (C_PF1_ENTRY_VERSION_TYPE_12       ),
			.C_PF1_ENTRY_RSVD0_12                 (C_PF1_ENTRY_RSVD0_12              ),
			.C_PF1_ENTRY_TYPE_13                  (C_PF1_ENTRY_TYPE_13               ),
			.C_PF1_ENTRY_BAR_13                   (C_PF1_ENTRY_BAR_13                ),
			.C_PF1_ENTRY_ADDR_13                  (C_PF1_ENTRY_ADDR_13               ),
			.C_PF1_ENTRY_MAJOR_VERSION_13         (C_PF1_ENTRY_MAJOR_VERSION_13      ),
			.C_PF1_ENTRY_MINOR_VERSION_13         (C_PF1_ENTRY_MINOR_VERSION_13      ),
			.C_PF1_ENTRY_VERSION_TYPE_13          (C_PF1_ENTRY_VERSION_TYPE_13       ),
			.C_PF1_ENTRY_RSVD0_13                 (C_PF1_ENTRY_RSVD0_13              ),
			.C_PF1_ENTRY_TYPE_14                  (C_PF1_ENTRY_TYPE_14               ),
			.C_PF1_ENTRY_BAR_14                   (C_PF1_ENTRY_BAR_14                ),
			.C_PF1_ENTRY_ADDR_14                  (C_PF1_ENTRY_ADDR_14               ),
			.C_PF1_ENTRY_MAJOR_VERSION_14         (C_PF1_ENTRY_MAJOR_VERSION_14      ),
			.C_PF1_ENTRY_MINOR_VERSION_14         (C_PF1_ENTRY_MINOR_VERSION_14      ),
			.C_PF1_ENTRY_VERSION_TYPE_14          (C_PF1_ENTRY_VERSION_TYPE_14       ),
			.C_PF1_ENTRY_RSVD0_14                 (C_PF1_ENTRY_RSVD0_14              ),
			.C_PF1_ENTRY_TYPE_15                  (C_PF1_ENTRY_TYPE_15               ),
			.C_PF1_ENTRY_BAR_15                   (C_PF1_ENTRY_BAR_15                ),
			.C_PF1_ENTRY_ADDR_15                  (C_PF1_ENTRY_ADDR_15               ),
			.C_PF1_ENTRY_MAJOR_VERSION_15         (C_PF1_ENTRY_MAJOR_VERSION_15      ),
			.C_PF1_ENTRY_MINOR_VERSION_15         (C_PF1_ENTRY_MINOR_VERSION_15      ),
			.C_PF1_ENTRY_VERSION_TYPE_15          (C_PF1_ENTRY_VERSION_TYPE_15       ),
			.C_PF1_ENTRY_RSVD0_15                 (C_PF1_ENTRY_RSVD0_15              ),
			.C_PF1_S_AXI_DATA_WIDTH               (C_PF1_S_AXI_DATA_WIDTH            ),
			.C_PF1_S_AXI_ADDR_WIDTH               (C_PF1_S_AXI_ADDR_WIDTH            ),
			.C_PF2_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF2_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF2_HAS_UUID_ROM	                  (C_PF2_HAS_UUID_ROM	               ),
			.C_PF2_BAR_INDEX               		    (C_PF2_BAR_INDEX               		 ),
			.C_PF2_LOW_OFFSET              		    (C_PF2_LOW_OFFSET              		 ),
			.C_PF2_HIGH_OFFSET             		    (C_PF2_HIGH_OFFSET             		 ),
			.C_PF2_UUID_ROM_INIT                  (C_PF2_UUID_ROM_INIT               ),
			.C_PF2_ENTRY_TYPE_0                   (C_PF2_ENTRY_TYPE_0                ),
			.C_PF2_ENTRY_BAR_0                    (C_PF2_ENTRY_BAR_0                 ),
			.C_PF2_ENTRY_ADDR_0                   (C_PF2_ENTRY_ADDR_0                ),
			.C_PF2_ENTRY_MAJOR_VERSION_0          (C_PF2_ENTRY_MAJOR_VERSION_0       ),
			.C_PF2_ENTRY_MINOR_VERSION_0          (C_PF2_ENTRY_MINOR_VERSION_0       ),
			.C_PF2_ENTRY_VERSION_TYPE_0           (C_PF2_ENTRY_VERSION_TYPE_0        ),
			.C_PF2_ENTRY_RSVD0_0                  (C_PF2_ENTRY_RSVD0_0               ),
			.C_PF2_ENTRY_TYPE_1                   (C_PF2_ENTRY_TYPE_1                ),
			.C_PF2_ENTRY_BAR_1                    (C_PF2_ENTRY_BAR_1                 ),
			.C_PF2_ENTRY_ADDR_1                   (C_PF2_ENTRY_ADDR_1                ),
			.C_PF2_ENTRY_MAJOR_VERSION_1          (C_PF2_ENTRY_MAJOR_VERSION_1       ),
			.C_PF2_ENTRY_MINOR_VERSION_1          (C_PF2_ENTRY_MINOR_VERSION_1       ),
			.C_PF2_ENTRY_VERSION_TYPE_1           (C_PF2_ENTRY_VERSION_TYPE_1        ),
			.C_PF2_ENTRY_RSVD0_1                  (C_PF2_ENTRY_RSVD0_1               ),
			.C_PF2_ENTRY_TYPE_2                   (C_PF2_ENTRY_TYPE_2                ),
			.C_PF2_ENTRY_BAR_2                    (C_PF2_ENTRY_BAR_2                 ),
			.C_PF2_ENTRY_ADDR_2                   (C_PF2_ENTRY_ADDR_2                ),
			.C_PF2_ENTRY_MAJOR_VERSION_2          (C_PF2_ENTRY_MAJOR_VERSION_2       ),
			.C_PF2_ENTRY_MINOR_VERSION_2          (C_PF2_ENTRY_MINOR_VERSION_2       ),
			.C_PF2_ENTRY_VERSION_TYPE_2           (C_PF2_ENTRY_VERSION_TYPE_2        ),
			.C_PF2_ENTRY_RSVD0_2                  (C_PF2_ENTRY_RSVD0_2               ),
			.C_PF2_ENTRY_TYPE_3                   (C_PF2_ENTRY_TYPE_3                ),
			.C_PF2_ENTRY_BAR_3                    (C_PF2_ENTRY_BAR_3                 ),
			.C_PF2_ENTRY_ADDR_3                   (C_PF2_ENTRY_ADDR_3                ),
			.C_PF2_ENTRY_MAJOR_VERSION_3          (C_PF2_ENTRY_MAJOR_VERSION_3       ),
			.C_PF2_ENTRY_MINOR_VERSION_3          (C_PF2_ENTRY_MINOR_VERSION_3       ),
			.C_PF2_ENTRY_VERSION_TYPE_3           (C_PF2_ENTRY_VERSION_TYPE_3        ),
			.C_PF2_ENTRY_RSVD0_3                  (C_PF2_ENTRY_RSVD0_3               ),
			.C_PF2_ENTRY_TYPE_4                   (C_PF2_ENTRY_TYPE_4                ),
			.C_PF2_ENTRY_BAR_4                    (C_PF2_ENTRY_BAR_4                 ),
			.C_PF2_ENTRY_ADDR_4                   (C_PF2_ENTRY_ADDR_4                ),
			.C_PF2_ENTRY_MAJOR_VERSION_4          (C_PF2_ENTRY_MAJOR_VERSION_4       ),
			.C_PF2_ENTRY_MINOR_VERSION_4          (C_PF2_ENTRY_MINOR_VERSION_4       ),
			.C_PF2_ENTRY_VERSION_TYPE_4           (C_PF2_ENTRY_VERSION_TYPE_4        ),
			.C_PF2_ENTRY_RSVD0_4                  (C_PF2_ENTRY_RSVD0_4               ),
			.C_PF2_ENTRY_TYPE_5                   (C_PF2_ENTRY_TYPE_5                ),
			.C_PF2_ENTRY_BAR_5                    (C_PF2_ENTRY_BAR_5                 ),
			.C_PF2_ENTRY_ADDR_5                   (C_PF2_ENTRY_ADDR_5                ),
			.C_PF2_ENTRY_MAJOR_VERSION_5          (C_PF2_ENTRY_MAJOR_VERSION_5       ),
			.C_PF2_ENTRY_MINOR_VERSION_5          (C_PF2_ENTRY_MINOR_VERSION_5       ),
			.C_PF2_ENTRY_VERSION_TYPE_5           (C_PF2_ENTRY_VERSION_TYPE_5        ),
			.C_PF2_ENTRY_RSVD0_5                  (C_PF2_ENTRY_RSVD0_5               ),
			.C_PF2_ENTRY_TYPE_6                   (C_PF2_ENTRY_TYPE_6                ),
			.C_PF2_ENTRY_BAR_6                    (C_PF2_ENTRY_BAR_6                 ),
			.C_PF2_ENTRY_ADDR_6                   (C_PF2_ENTRY_ADDR_6                ),
			.C_PF2_ENTRY_MAJOR_VERSION_6          (C_PF2_ENTRY_MAJOR_VERSION_6       ),
			.C_PF2_ENTRY_MINOR_VERSION_6          (C_PF2_ENTRY_MINOR_VERSION_6       ),
			.C_PF2_ENTRY_VERSION_TYPE_6           (C_PF2_ENTRY_VERSION_TYPE_6        ),
			.C_PF2_ENTRY_RSVD0_6                  (C_PF2_ENTRY_RSVD0_6               ),
			.C_PF2_ENTRY_TYPE_7                   (C_PF2_ENTRY_TYPE_7                ),
			.C_PF2_ENTRY_BAR_7                    (C_PF2_ENTRY_BAR_7                 ),
			.C_PF2_ENTRY_ADDR_7                   (C_PF2_ENTRY_ADDR_7                ),
			.C_PF2_ENTRY_MAJOR_VERSION_7          (C_PF2_ENTRY_MAJOR_VERSION_7       ),
			.C_PF2_ENTRY_MINOR_VERSION_7          (C_PF2_ENTRY_MINOR_VERSION_7       ),
			.C_PF2_ENTRY_VERSION_TYPE_7           (C_PF2_ENTRY_VERSION_TYPE_7        ),
			.C_PF2_ENTRY_RSVD0_7                  (C_PF2_ENTRY_RSVD0_7               ),
			.C_PF2_ENTRY_TYPE_8                   (C_PF2_ENTRY_TYPE_8                ),
			.C_PF2_ENTRY_BAR_8                    (C_PF2_ENTRY_BAR_8                 ),
			.C_PF2_ENTRY_ADDR_8                   (C_PF2_ENTRY_ADDR_8                ),
			.C_PF2_ENTRY_MAJOR_VERSION_8          (C_PF2_ENTRY_MAJOR_VERSION_8       ),
			.C_PF2_ENTRY_MINOR_VERSION_8          (C_PF2_ENTRY_MINOR_VERSION_8       ),
			.C_PF2_ENTRY_VERSION_TYPE_8           (C_PF2_ENTRY_VERSION_TYPE_8        ),
			.C_PF2_ENTRY_RSVD0_8                  (C_PF2_ENTRY_RSVD0_8               ),
			.C_PF2_ENTRY_TYPE_9                   (C_PF2_ENTRY_TYPE_9                ),
			.C_PF2_ENTRY_BAR_9                    (C_PF2_ENTRY_BAR_9                 ),
			.C_PF2_ENTRY_ADDR_9                   (C_PF2_ENTRY_ADDR_9                ),
			.C_PF2_ENTRY_MAJOR_VERSION_9          (C_PF2_ENTRY_MAJOR_VERSION_9       ),
			.C_PF2_ENTRY_MINOR_VERSION_9          (C_PF2_ENTRY_MINOR_VERSION_9       ),
			.C_PF2_ENTRY_VERSION_TYPE_9           (C_PF2_ENTRY_VERSION_TYPE_9        ),
			.C_PF2_ENTRY_RSVD0_9                  (C_PF2_ENTRY_RSVD0_9               ),
			.C_PF2_ENTRY_TYPE_10                  (C_PF2_ENTRY_TYPE_10               ),
			.C_PF2_ENTRY_BAR_10                   (C_PF2_ENTRY_BAR_10                ),
			.C_PF2_ENTRY_ADDR_10                  (C_PF2_ENTRY_ADDR_10               ),
			.C_PF2_ENTRY_MAJOR_VERSION_10         (C_PF2_ENTRY_MAJOR_VERSION_10      ),
			.C_PF2_ENTRY_MINOR_VERSION_10         (C_PF2_ENTRY_MINOR_VERSION_10      ),
			.C_PF2_ENTRY_VERSION_TYPE_10          (C_PF2_ENTRY_VERSION_TYPE_10       ),
			.C_PF2_ENTRY_RSVD0_10                 (C_PF2_ENTRY_RSVD0_10              ),
			.C_PF2_ENTRY_TYPE_11                  (C_PF2_ENTRY_TYPE_11               ),
			.C_PF2_ENTRY_BAR_11                   (C_PF2_ENTRY_BAR_11                ),
			.C_PF2_ENTRY_ADDR_11                  (C_PF2_ENTRY_ADDR_11               ),
			.C_PF2_ENTRY_MAJOR_VERSION_11         (C_PF2_ENTRY_MAJOR_VERSION_11      ),
			.C_PF2_ENTRY_MINOR_VERSION_11         (C_PF2_ENTRY_MINOR_VERSION_11      ),
			.C_PF2_ENTRY_VERSION_TYPE_11          (C_PF2_ENTRY_VERSION_TYPE_11       ),
			.C_PF2_ENTRY_RSVD0_11                 (C_PF2_ENTRY_RSVD0_11              ),
			.C_PF2_ENTRY_TYPE_12                  (C_PF2_ENTRY_TYPE_12               ),
			.C_PF2_ENTRY_BAR_12                   (C_PF2_ENTRY_BAR_12                ),
			.C_PF2_ENTRY_ADDR_12                  (C_PF2_ENTRY_ADDR_12               ),
			.C_PF2_ENTRY_MAJOR_VERSION_12         (C_PF2_ENTRY_MAJOR_VERSION_12      ),
			.C_PF2_ENTRY_MINOR_VERSION_12         (C_PF2_ENTRY_MINOR_VERSION_12      ),
			.C_PF2_ENTRY_VERSION_TYPE_12          (C_PF2_ENTRY_VERSION_TYPE_12       ),
			.C_PF2_ENTRY_RSVD0_12                 (C_PF2_ENTRY_RSVD0_12              ),
			.C_PF2_ENTRY_TYPE_13                  (C_PF2_ENTRY_TYPE_13               ),
			.C_PF2_ENTRY_BAR_13                   (C_PF2_ENTRY_BAR_13                ),
			.C_PF2_ENTRY_ADDR_13                  (C_PF2_ENTRY_ADDR_13               ),
			.C_PF2_ENTRY_MAJOR_VERSION_13         (C_PF2_ENTRY_MAJOR_VERSION_13      ),
			.C_PF2_ENTRY_MINOR_VERSION_13         (C_PF2_ENTRY_MINOR_VERSION_13      ),
			.C_PF2_ENTRY_VERSION_TYPE_13          (C_PF2_ENTRY_VERSION_TYPE_13       ),
			.C_PF2_ENTRY_RSVD0_13                 (C_PF2_ENTRY_RSVD0_13              ),
			.C_PF2_ENTRY_TYPE_14                  (C_PF2_ENTRY_TYPE_14               ),
			.C_PF2_ENTRY_BAR_14                   (C_PF2_ENTRY_BAR_14                ),
			.C_PF2_ENTRY_ADDR_14                  (C_PF2_ENTRY_ADDR_14               ),
			.C_PF2_ENTRY_MAJOR_VERSION_14         (C_PF2_ENTRY_MAJOR_VERSION_14      ),
			.C_PF2_ENTRY_MINOR_VERSION_14         (C_PF2_ENTRY_MINOR_VERSION_14      ),
			.C_PF2_ENTRY_VERSION_TYPE_14          (C_PF2_ENTRY_VERSION_TYPE_14       ),
			.C_PF2_ENTRY_RSVD0_14                 (C_PF2_ENTRY_RSVD0_14              ),
			.C_PF2_ENTRY_TYPE_15                  (C_PF2_ENTRY_TYPE_15               ),
			.C_PF2_ENTRY_BAR_15                   (C_PF2_ENTRY_BAR_15                ),
			.C_PF2_ENTRY_ADDR_15                  (C_PF2_ENTRY_ADDR_15               ),
			.C_PF2_ENTRY_MAJOR_VERSION_15         (C_PF2_ENTRY_MAJOR_VERSION_15      ),
			.C_PF2_ENTRY_MINOR_VERSION_15         (C_PF2_ENTRY_MINOR_VERSION_15      ),
			.C_PF2_ENTRY_VERSION_TYPE_15          (C_PF2_ENTRY_VERSION_TYPE_15       ),
			.C_PF2_ENTRY_RSVD0_15                 (C_PF2_ENTRY_RSVD0_15              ),
			.C_PF2_S_AXI_DATA_WIDTH               (C_PF2_S_AXI_DATA_WIDTH            ),
			.C_PF2_S_AXI_ADDR_WIDTH               (C_PF2_S_AXI_ADDR_WIDTH            ),
			.C_PF3_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF3_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF3_HAS_UUID_ROM	                  (C_PF3_HAS_UUID_ROM	               ),
			.C_PF3_BAR_INDEX               		    (C_PF3_BAR_INDEX               		 ),
			.C_PF3_LOW_OFFSET              		    (C_PF3_LOW_OFFSET              		 ),
			.C_PF3_HIGH_OFFSET             		    (C_PF3_HIGH_OFFSET             		 ),
			.C_PF3_UUID_ROM_INIT                  (C_PF3_UUID_ROM_INIT               ),
			.C_PF3_ENTRY_TYPE_0                   (C_PF3_ENTRY_TYPE_0                ),
			.C_PF3_ENTRY_BAR_0                    (C_PF3_ENTRY_BAR_0                 ),
			.C_PF3_ENTRY_ADDR_0                   (C_PF3_ENTRY_ADDR_0                ),
			.C_PF3_ENTRY_MAJOR_VERSION_0          (C_PF3_ENTRY_MAJOR_VERSION_0       ),
			.C_PF3_ENTRY_MINOR_VERSION_0          (C_PF3_ENTRY_MINOR_VERSION_0       ),
			.C_PF3_ENTRY_VERSION_TYPE_0           (C_PF3_ENTRY_VERSION_TYPE_0        ),
			.C_PF3_ENTRY_RSVD0_0                  (C_PF3_ENTRY_RSVD0_0               ),
			.C_PF3_ENTRY_TYPE_1                   (C_PF3_ENTRY_TYPE_1                ),
			.C_PF3_ENTRY_BAR_1                    (C_PF3_ENTRY_BAR_1                 ),
			.C_PF3_ENTRY_ADDR_1                   (C_PF3_ENTRY_ADDR_1                ),
			.C_PF3_ENTRY_MAJOR_VERSION_1          (C_PF3_ENTRY_MAJOR_VERSION_1       ),
			.C_PF3_ENTRY_MINOR_VERSION_1          (C_PF3_ENTRY_MINOR_VERSION_1       ),
			.C_PF3_ENTRY_VERSION_TYPE_1           (C_PF3_ENTRY_VERSION_TYPE_1        ),
			.C_PF3_ENTRY_RSVD0_1                  (C_PF3_ENTRY_RSVD0_1               ),
			.C_PF3_ENTRY_TYPE_2                   (C_PF3_ENTRY_TYPE_2                ),
			.C_PF3_ENTRY_BAR_2                    (C_PF3_ENTRY_BAR_2                 ),
			.C_PF3_ENTRY_ADDR_2                   (C_PF3_ENTRY_ADDR_2                ),
			.C_PF3_ENTRY_MAJOR_VERSION_2          (C_PF3_ENTRY_MAJOR_VERSION_2       ),
			.C_PF3_ENTRY_MINOR_VERSION_2          (C_PF3_ENTRY_MINOR_VERSION_2       ),
			.C_PF3_ENTRY_VERSION_TYPE_2           (C_PF3_ENTRY_VERSION_TYPE_2        ),
			.C_PF3_ENTRY_RSVD0_2                  (C_PF3_ENTRY_RSVD0_2               ),
			.C_PF3_ENTRY_TYPE_3                   (C_PF3_ENTRY_TYPE_3                ),
			.C_PF3_ENTRY_BAR_3                    (C_PF3_ENTRY_BAR_3                 ),
			.C_PF3_ENTRY_ADDR_3                   (C_PF3_ENTRY_ADDR_3                ),
			.C_PF3_ENTRY_MAJOR_VERSION_3          (C_PF3_ENTRY_MAJOR_VERSION_3       ),
			.C_PF3_ENTRY_MINOR_VERSION_3          (C_PF3_ENTRY_MINOR_VERSION_3       ),
			.C_PF3_ENTRY_VERSION_TYPE_3           (C_PF3_ENTRY_VERSION_TYPE_3        ),
			.C_PF3_ENTRY_RSVD0_3                  (C_PF3_ENTRY_RSVD0_3               ),
			.C_PF3_ENTRY_TYPE_4                   (C_PF3_ENTRY_TYPE_4                ),
			.C_PF3_ENTRY_BAR_4                    (C_PF3_ENTRY_BAR_4                 ),
			.C_PF3_ENTRY_ADDR_4                   (C_PF3_ENTRY_ADDR_4                ),
			.C_PF3_ENTRY_MAJOR_VERSION_4          (C_PF3_ENTRY_MAJOR_VERSION_4       ),
			.C_PF3_ENTRY_MINOR_VERSION_4          (C_PF3_ENTRY_MINOR_VERSION_4       ),
			.C_PF3_ENTRY_VERSION_TYPE_4           (C_PF3_ENTRY_VERSION_TYPE_4        ),
			.C_PF3_ENTRY_RSVD0_4                  (C_PF3_ENTRY_RSVD0_4               ),
			.C_PF3_ENTRY_TYPE_5                   (C_PF3_ENTRY_TYPE_5                ),
			.C_PF3_ENTRY_BAR_5                    (C_PF3_ENTRY_BAR_5                 ),
			.C_PF3_ENTRY_ADDR_5                   (C_PF3_ENTRY_ADDR_5                ),
			.C_PF3_ENTRY_MAJOR_VERSION_5          (C_PF3_ENTRY_MAJOR_VERSION_5       ),
			.C_PF3_ENTRY_MINOR_VERSION_5          (C_PF3_ENTRY_MINOR_VERSION_5       ),
			.C_PF3_ENTRY_VERSION_TYPE_5           (C_PF3_ENTRY_VERSION_TYPE_5        ),
			.C_PF3_ENTRY_RSVD0_5                  (C_PF3_ENTRY_RSVD0_5               ),
			.C_PF3_ENTRY_TYPE_6                   (C_PF3_ENTRY_TYPE_6                ),
			.C_PF3_ENTRY_BAR_6                    (C_PF3_ENTRY_BAR_6                 ),
			.C_PF3_ENTRY_ADDR_6                   (C_PF3_ENTRY_ADDR_6                ),
			.C_PF3_ENTRY_MAJOR_VERSION_6          (C_PF3_ENTRY_MAJOR_VERSION_6       ),
			.C_PF3_ENTRY_MINOR_VERSION_6          (C_PF3_ENTRY_MINOR_VERSION_6       ),
			.C_PF3_ENTRY_VERSION_TYPE_6           (C_PF3_ENTRY_VERSION_TYPE_6        ),
			.C_PF3_ENTRY_RSVD0_6                  (C_PF3_ENTRY_RSVD0_6               ),
			.C_PF3_ENTRY_TYPE_7                   (C_PF3_ENTRY_TYPE_7                ),
			.C_PF3_ENTRY_BAR_7                    (C_PF3_ENTRY_BAR_7                 ),
			.C_PF3_ENTRY_ADDR_7                   (C_PF3_ENTRY_ADDR_7                ),
			.C_PF3_ENTRY_MAJOR_VERSION_7          (C_PF3_ENTRY_MAJOR_VERSION_7       ),
			.C_PF3_ENTRY_MINOR_VERSION_7          (C_PF3_ENTRY_MINOR_VERSION_7       ),
			.C_PF3_ENTRY_VERSION_TYPE_7           (C_PF3_ENTRY_VERSION_TYPE_7        ),
			.C_PF3_ENTRY_RSVD0_7                  (C_PF3_ENTRY_RSVD0_7               ),
			.C_PF3_ENTRY_TYPE_8                   (C_PF3_ENTRY_TYPE_8                ),
			.C_PF3_ENTRY_BAR_8                    (C_PF3_ENTRY_BAR_8                 ),
			.C_PF3_ENTRY_ADDR_8                   (C_PF3_ENTRY_ADDR_8                ),
			.C_PF3_ENTRY_MAJOR_VERSION_8          (C_PF3_ENTRY_MAJOR_VERSION_8       ),
			.C_PF3_ENTRY_MINOR_VERSION_8          (C_PF3_ENTRY_MINOR_VERSION_8       ),
			.C_PF3_ENTRY_VERSION_TYPE_8           (C_PF3_ENTRY_VERSION_TYPE_8        ),
			.C_PF3_ENTRY_RSVD0_8                  (C_PF3_ENTRY_RSVD0_8               ),
			.C_PF3_ENTRY_TYPE_9                   (C_PF3_ENTRY_TYPE_9                ),
			.C_PF3_ENTRY_BAR_9                    (C_PF3_ENTRY_BAR_9                 ),
			.C_PF3_ENTRY_ADDR_9                   (C_PF3_ENTRY_ADDR_9                ),
			.C_PF3_ENTRY_MAJOR_VERSION_9          (C_PF3_ENTRY_MAJOR_VERSION_9       ),
			.C_PF3_ENTRY_MINOR_VERSION_9          (C_PF3_ENTRY_MINOR_VERSION_9       ),
			.C_PF3_ENTRY_VERSION_TYPE_9           (C_PF3_ENTRY_VERSION_TYPE_9        ),
			.C_PF3_ENTRY_RSVD0_9                  (C_PF3_ENTRY_RSVD0_9               ),
			.C_PF3_ENTRY_TYPE_10                  (C_PF3_ENTRY_TYPE_10               ),
			.C_PF3_ENTRY_BAR_10                   (C_PF3_ENTRY_BAR_10                ),
			.C_PF3_ENTRY_ADDR_10                  (C_PF3_ENTRY_ADDR_10               ),
			.C_PF3_ENTRY_MAJOR_VERSION_10         (C_PF3_ENTRY_MAJOR_VERSION_10      ),
			.C_PF3_ENTRY_MINOR_VERSION_10         (C_PF3_ENTRY_MINOR_VERSION_10      ),
			.C_PF3_ENTRY_VERSION_TYPE_10          (C_PF3_ENTRY_VERSION_TYPE_10       ),
			.C_PF3_ENTRY_RSVD0_10                 (C_PF3_ENTRY_RSVD0_10              ),
			.C_PF3_ENTRY_TYPE_11                  (C_PF3_ENTRY_TYPE_11               ),
			.C_PF3_ENTRY_BAR_11                   (C_PF3_ENTRY_BAR_11                ),
			.C_PF3_ENTRY_ADDR_11                  (C_PF3_ENTRY_ADDR_11               ),
			.C_PF3_ENTRY_MAJOR_VERSION_11         (C_PF3_ENTRY_MAJOR_VERSION_11      ),
			.C_PF3_ENTRY_MINOR_VERSION_11         (C_PF3_ENTRY_MINOR_VERSION_11      ),
			.C_PF3_ENTRY_VERSION_TYPE_11          (C_PF3_ENTRY_VERSION_TYPE_11       ),
			.C_PF3_ENTRY_RSVD0_11                 (C_PF3_ENTRY_RSVD0_11              ),
			.C_PF3_ENTRY_TYPE_12                  (C_PF3_ENTRY_TYPE_12               ),
			.C_PF3_ENTRY_BAR_12                   (C_PF3_ENTRY_BAR_12                ),
			.C_PF3_ENTRY_ADDR_12                  (C_PF3_ENTRY_ADDR_12               ),
			.C_PF3_ENTRY_MAJOR_VERSION_12         (C_PF3_ENTRY_MAJOR_VERSION_12      ),
			.C_PF3_ENTRY_MINOR_VERSION_12         (C_PF3_ENTRY_MINOR_VERSION_12      ),
			.C_PF3_ENTRY_VERSION_TYPE_12          (C_PF3_ENTRY_VERSION_TYPE_12       ),
			.C_PF3_ENTRY_RSVD0_12                 (C_PF3_ENTRY_RSVD0_12              ),
			.C_PF3_ENTRY_TYPE_13                  (C_PF3_ENTRY_TYPE_13               ),
			.C_PF3_ENTRY_BAR_13                   (C_PF3_ENTRY_BAR_13                ),
			.C_PF3_ENTRY_ADDR_13                  (C_PF3_ENTRY_ADDR_13               ),
			.C_PF3_ENTRY_MAJOR_VERSION_13         (C_PF3_ENTRY_MAJOR_VERSION_13      ),
			.C_PF3_ENTRY_MINOR_VERSION_13         (C_PF3_ENTRY_MINOR_VERSION_13      ),
			.C_PF3_ENTRY_VERSION_TYPE_13          (C_PF3_ENTRY_VERSION_TYPE_13       ),
			.C_PF3_ENTRY_RSVD0_13                 (C_PF3_ENTRY_RSVD0_13              ),
			.C_PF3_ENTRY_TYPE_14                  (C_PF3_ENTRY_TYPE_14               ),
			.C_PF3_ENTRY_BAR_14                   (C_PF3_ENTRY_BAR_14                ),
			.C_PF3_ENTRY_ADDR_14                  (C_PF3_ENTRY_ADDR_14               ),
			.C_PF3_ENTRY_MAJOR_VERSION_14         (C_PF3_ENTRY_MAJOR_VERSION_14      ),
			.C_PF3_ENTRY_MINOR_VERSION_14         (C_PF3_ENTRY_MINOR_VERSION_14      ),
			.C_PF3_ENTRY_VERSION_TYPE_14          (C_PF3_ENTRY_VERSION_TYPE_14       ),
			.C_PF3_ENTRY_RSVD0_14                 (C_PF3_ENTRY_RSVD0_14              ),
			.C_PF3_ENTRY_TYPE_15                  (C_PF3_ENTRY_TYPE_15               ),
			.C_PF3_ENTRY_BAR_15                   (C_PF3_ENTRY_BAR_15                ),
			.C_PF3_ENTRY_ADDR_15                  (C_PF3_ENTRY_ADDR_15               ),
			.C_PF3_ENTRY_MAJOR_VERSION_15         (C_PF3_ENTRY_MAJOR_VERSION_15      ),
			.C_PF3_ENTRY_MINOR_VERSION_15         (C_PF3_ENTRY_MINOR_VERSION_15      ),
			.C_PF3_ENTRY_VERSION_TYPE_15          (C_PF3_ENTRY_VERSION_TYPE_15       ),
			.C_PF3_ENTRY_RSVD0_15                 (C_PF3_ENTRY_RSVD0_15              ),
			.C_PF3_S_AXI_DATA_WIDTH               (C_PF3_S_AXI_DATA_WIDTH            ),
			.C_PF3_S_AXI_ADDR_WIDTH               (C_PF3_S_AXI_ADDR_WIDTH            ),
			.C_XDEVICEFAMILY                      (C_XDEVICEFAMILY                   )
    ) hw_disc_inst (
      .aclk_pcie     												(aclk_pcie                         ),   
      .aresetn_pcie  												(aresetn_pcie                      ),          
      .aclk_ctrl     												(aclk_ctrl                         ),
      .aresetn_ctrl  												(aresetn_ctrl                      ),
      .s_pcie4_cfg_ext_function_number      (s_pcie4_cfg_ext_function_number   ),
      .s_pcie4_cfg_ext_read_data            (s_pcie4_cfg_ext_read_data         ),
      .s_pcie4_cfg_ext_read_data_valid      (s_pcie4_cfg_ext_read_data_valid   ),
      .s_pcie4_cfg_ext_read_received        (s_pcie4_cfg_ext_read_received     ),
      .s_pcie4_cfg_ext_register_number      (s_pcie4_cfg_ext_register_number   ),
      .s_pcie4_cfg_ext_write_byte_enable    (s_pcie4_cfg_ext_write_byte_enable ),
      .s_pcie4_cfg_ext_write_data           (s_pcie4_cfg_ext_write_data        ),
      .s_pcie4_cfg_ext_write_received       (s_pcie4_cfg_ext_write_received    ),
      .m_pcie4_cfg_ext_function_number      (m_pcie4_cfg_ext_function_number   ),
      .m_pcie4_cfg_ext_read_data            (m_pcie4_cfg_ext_read_data         ),
      .m_pcie4_cfg_ext_read_data_valid      (m_pcie4_cfg_ext_read_data_valid   ),
      .m_pcie4_cfg_ext_read_received        (m_pcie4_cfg_ext_read_received     ),
      .m_pcie4_cfg_ext_register_number      (m_pcie4_cfg_ext_register_number   ),
      .m_pcie4_cfg_ext_write_byte_enable    (m_pcie4_cfg_ext_write_byte_enable ),
      .m_pcie4_cfg_ext_write_data           (m_pcie4_cfg_ext_write_data        ),      
      .m_pcie4_cfg_ext_write_received       (m_pcie4_cfg_ext_write_received    ),
      .s_axi_ctrl_pf0_AWADDR                (s_axi_ctrl_pf0_AWADDR             ),
      .s_axi_ctrl_pf0_AWVALID               (s_axi_ctrl_pf0_AWVALID            ),
      .s_axi_ctrl_pf0_AWREADY               (s_axi_ctrl_pf0_AWREADY            ),
      .s_axi_ctrl_pf0_WDATA                 (s_axi_ctrl_pf0_WDATA              ),
      .s_axi_ctrl_pf0_WSTRB                 (s_axi_ctrl_pf0_WSTRB              ),
      .s_axi_ctrl_pf0_WVALID                (s_axi_ctrl_pf0_WVALID             ),
      .s_axi_ctrl_pf0_WREADY                (s_axi_ctrl_pf0_WREADY             ),
      .s_axi_ctrl_pf0_BRESP                 (s_axi_ctrl_pf0_BRESP              ),
      .s_axi_ctrl_pf0_BVALID                (s_axi_ctrl_pf0_BVALID             ),
      .s_axi_ctrl_pf0_BREADY                (s_axi_ctrl_pf0_BREADY             ),
      .s_axi_ctrl_pf0_ARADDR                (s_axi_ctrl_pf0_ARADDR             ),
      .s_axi_ctrl_pf0_ARVALID               (s_axi_ctrl_pf0_ARVALID            ),
      .s_axi_ctrl_pf0_ARREADY               (s_axi_ctrl_pf0_ARREADY            ),
      .s_axi_ctrl_pf0_RDATA                 (s_axi_ctrl_pf0_RDATA              ),
      .s_axi_ctrl_pf0_RRESP                 (s_axi_ctrl_pf0_RRESP              ),
      .s_axi_ctrl_pf0_RVALID                (s_axi_ctrl_pf0_RVALID             ),
      .s_axi_ctrl_pf0_RREADY                (s_axi_ctrl_pf0_RREADY             ),
      .s_axi_ctrl_pf1_AWADDR                (s_axi_ctrl_pf1_AWADDR             ),
      .s_axi_ctrl_pf1_AWVALID               (s_axi_ctrl_pf1_AWVALID            ),
      .s_axi_ctrl_pf1_AWREADY               (s_axi_ctrl_pf1_AWREADY            ),
      .s_axi_ctrl_pf1_WDATA                 (s_axi_ctrl_pf1_WDATA              ),
      .s_axi_ctrl_pf1_WSTRB                 (s_axi_ctrl_pf1_WSTRB              ),
      .s_axi_ctrl_pf1_WVALID                (s_axi_ctrl_pf1_WVALID             ),
      .s_axi_ctrl_pf1_WREADY                (s_axi_ctrl_pf1_WREADY             ),
      .s_axi_ctrl_pf1_BRESP                 (s_axi_ctrl_pf1_BRESP              ),
      .s_axi_ctrl_pf1_BVALID                (s_axi_ctrl_pf1_BVALID             ),
      .s_axi_ctrl_pf1_BREADY                (s_axi_ctrl_pf1_BREADY             ),
      .s_axi_ctrl_pf1_ARADDR                (s_axi_ctrl_pf1_ARADDR             ),
      .s_axi_ctrl_pf1_ARVALID               (s_axi_ctrl_pf1_ARVALID            ),
      .s_axi_ctrl_pf1_ARREADY               (s_axi_ctrl_pf1_ARREADY            ),
      .s_axi_ctrl_pf1_RDATA                 (s_axi_ctrl_pf1_RDATA              ),
      .s_axi_ctrl_pf1_RRESP                 (s_axi_ctrl_pf1_RRESP              ),
      .s_axi_ctrl_pf1_RVALID                (s_axi_ctrl_pf1_RVALID             ),
      .s_axi_ctrl_pf1_RREADY                (s_axi_ctrl_pf1_RREADY             ),
      .s_axi_ctrl_pf2_AWADDR                (s_axi_ctrl_pf2_AWADDR             ),
      .s_axi_ctrl_pf2_AWVALID               (s_axi_ctrl_pf2_AWVALID            ),
      .s_axi_ctrl_pf2_AWREADY               (s_axi_ctrl_pf2_AWREADY            ),
      .s_axi_ctrl_pf2_WDATA                 (s_axi_ctrl_pf2_WDATA              ),
      .s_axi_ctrl_pf2_WSTRB                 (s_axi_ctrl_pf2_WSTRB              ),
      .s_axi_ctrl_pf2_WVALID                (s_axi_ctrl_pf2_WVALID             ),
      .s_axi_ctrl_pf2_WREADY                (s_axi_ctrl_pf2_WREADY             ),
      .s_axi_ctrl_pf2_BRESP                 (s_axi_ctrl_pf2_BRESP              ),
      .s_axi_ctrl_pf2_BVALID                (s_axi_ctrl_pf2_BVALID             ),
      .s_axi_ctrl_pf2_BREADY                (s_axi_ctrl_pf2_BREADY             ),
      .s_axi_ctrl_pf2_ARADDR                (s_axi_ctrl_pf2_ARADDR             ),
      .s_axi_ctrl_pf2_ARVALID               (s_axi_ctrl_pf2_ARVALID            ),
      .s_axi_ctrl_pf2_ARREADY               (s_axi_ctrl_pf2_ARREADY            ),
      .s_axi_ctrl_pf2_RDATA                 (s_axi_ctrl_pf2_RDATA              ),
      .s_axi_ctrl_pf2_RRESP                 (s_axi_ctrl_pf2_RRESP              ),
      .s_axi_ctrl_pf2_RVALID                (s_axi_ctrl_pf2_RVALID             ),
      .s_axi_ctrl_pf2_RREADY                (s_axi_ctrl_pf2_RREADY             ),
      .s_axi_ctrl_pf3_AWADDR                (s_axi_ctrl_pf3_AWADDR             ),
      .s_axi_ctrl_pf3_AWVALID               (s_axi_ctrl_pf3_AWVALID            ),
      .s_axi_ctrl_pf3_AWREADY               (s_axi_ctrl_pf3_AWREADY            ),
      .s_axi_ctrl_pf3_WDATA                 (s_axi_ctrl_pf3_WDATA              ),
      .s_axi_ctrl_pf3_WSTRB                 (s_axi_ctrl_pf3_WSTRB              ),
      .s_axi_ctrl_pf3_WVALID                (s_axi_ctrl_pf3_WVALID             ),
      .s_axi_ctrl_pf3_WREADY                (s_axi_ctrl_pf3_WREADY             ),
      .s_axi_ctrl_pf3_BRESP                 (s_axi_ctrl_pf3_BRESP              ),
      .s_axi_ctrl_pf3_BVALID                (s_axi_ctrl_pf3_BVALID             ),
      .s_axi_ctrl_pf3_BREADY                (s_axi_ctrl_pf3_BREADY             ),
      .s_axi_ctrl_pf3_ARADDR                (s_axi_ctrl_pf3_ARADDR             ),
      .s_axi_ctrl_pf3_ARVALID               (s_axi_ctrl_pf3_ARVALID            ),
      .s_axi_ctrl_pf3_ARREADY               (s_axi_ctrl_pf3_ARREADY            ),
      .s_axi_ctrl_pf3_RDATA                 (s_axi_ctrl_pf3_RDATA              ),
      .s_axi_ctrl_pf3_RRESP                 (s_axi_ctrl_pf3_RRESP              ),
      .s_axi_ctrl_pf3_RVALID                (s_axi_ctrl_pf3_RVALID             ),
      .s_axi_ctrl_pf3_RREADY                (s_axi_ctrl_pf3_RREADY             )
    );
    
endmodule


