// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689
`timescale 1ns / 1ps

module in_fifo_args #(
    parameter C_NUM_INPUT_FIFOs = 0,
    parameter [31:0] S_AXIS_FIFO_0_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_1_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_2_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_3_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_4_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_5_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_6_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_7_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_8_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_9_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_10_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_11_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_12_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_13_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_14_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_15_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_16_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_17_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_18_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_19_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_20_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_21_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_22_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_23_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_24_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_25_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_26_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_27_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_28_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_29_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_30_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_31_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_32_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_33_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_34_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_35_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_36_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_37_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_38_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_39_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_40_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_41_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_42_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_43_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_44_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_45_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_46_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_47_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_48_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_49_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_50_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_51_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_52_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_53_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_54_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_55_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_56_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_57_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_58_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_59_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_60_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_61_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_62_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_63_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_64_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_65_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_66_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_67_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_68_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_69_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_70_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_71_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_72_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_73_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_74_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_75_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_76_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_77_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_78_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_79_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_80_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_81_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_82_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_83_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_84_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_85_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_86_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_87_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_88_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_89_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_90_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_91_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_92_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_93_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_94_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_95_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_96_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_97_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_98_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_99_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_100_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_101_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_102_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_103_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_104_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_105_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_106_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_107_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_108_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_109_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_110_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_111_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_112_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_113_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_114_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_115_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_116_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_117_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_118_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_119_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_120_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_121_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_122_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_123_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_124_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_125_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_126_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_127_WIDTH = 8,     //width of input fifo interface on the accelerator, actual
    parameter [31:0] S_AXIS_FIFO_0_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_1_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_2_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_3_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_4_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_5_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_6_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_7_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_8_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_9_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_10_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_11_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_12_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_13_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_14_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_15_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_16_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_17_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_18_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_19_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_20_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_21_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_22_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_23_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_24_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_25_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_26_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_27_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_28_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_29_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_30_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_31_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_32_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_33_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_34_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_35_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_36_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_37_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_38_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_39_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_40_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_41_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_42_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_43_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_44_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_45_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_46_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_47_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_48_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_49_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_50_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_51_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_52_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_53_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_54_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_55_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_56_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_57_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_58_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_59_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_60_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_61_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_62_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_63_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_64_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_65_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_66_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_67_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_68_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_69_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_70_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_71_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_72_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_73_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_74_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_75_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_76_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_77_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_78_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_79_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_80_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_81_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_82_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_83_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_84_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_85_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_86_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_87_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_88_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_89_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_90_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_91_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_92_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_93_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_94_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_95_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_96_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_97_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_98_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_99_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_100_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_101_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_102_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_103_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_104_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_105_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_106_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_107_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_108_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_109_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_110_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_111_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_112_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_113_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_114_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_115_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_116_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_117_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_118_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_119_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_120_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_121_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_122_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_123_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_124_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_125_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_126_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_127_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_0_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_1_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_2_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_3_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_4_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_5_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_6_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_7_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_8_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_9_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_10_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_11_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_12_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_13_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_14_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_15_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_16_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_17_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_18_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_19_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_20_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_21_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_22_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_23_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_24_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_25_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_26_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_27_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_28_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_29_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_30_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_31_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_32_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_33_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_34_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_35_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_36_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_37_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_38_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_39_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_40_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_41_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_42_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_43_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_44_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_45_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_46_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_47_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_48_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_49_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_50_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_51_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_52_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_53_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_54_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_55_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_56_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_57_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_58_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_59_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_60_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_61_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_62_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_63_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_64_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_65_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_66_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_67_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_68_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_69_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_70_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_71_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_72_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_73_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_74_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_75_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_76_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_77_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_78_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_79_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_80_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_81_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_82_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_83_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_84_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_85_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_86_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_87_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_88_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_89_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_90_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_91_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_92_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_93_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_94_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_95_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_96_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_97_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_98_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_99_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_100_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_101_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_102_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_103_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_104_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_105_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_106_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_107_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_108_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_109_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_110_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_111_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_112_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_113_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_114_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_115_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_116_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_117_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_118_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_119_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_120_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_121_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_122_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_123_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_124_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_125_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_126_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_127_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_0_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_1_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_2_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_3_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_4_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_5_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_6_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_7_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_8_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_9_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_10_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_11_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_12_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_13_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_14_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_15_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_16_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_17_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_18_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_19_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_20_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_21_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_22_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_23_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_24_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_25_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_26_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_27_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_28_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_29_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_30_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_31_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_32_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_33_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_34_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_35_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_36_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_37_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_38_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_39_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_40_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_41_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_42_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_43_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_44_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_45_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_46_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_47_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_48_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_49_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_50_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_51_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_52_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_53_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_54_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_55_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_56_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_57_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_58_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_59_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_60_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_61_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_62_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_63_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_64_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_65_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_66_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_67_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_68_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_69_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_70_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_71_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_72_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_73_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_74_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_75_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_76_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_77_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_78_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_79_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_80_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_81_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_82_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_83_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_84_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_85_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_86_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_87_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_88_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_89_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_90_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_91_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_92_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_93_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_94_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_95_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_96_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_97_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_98_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_99_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_100_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_101_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_102_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_103_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_104_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_105_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_106_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_107_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_108_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_109_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_110_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_111_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_112_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_113_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_114_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_115_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_116_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_117_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_118_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_119_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_120_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_121_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_122_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_123_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_124_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_125_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_126_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_127_BYTE_WIDTH = 8     //width of input fifo interface on the accelerator, padded
 ) (
    input acc_clk,
    input acc_aresetn,
    //control interface
    input in_fifo_allow,
    output [C_NUM_INPUT_FIFOs-1:0] in_fifo_ready,
    output [C_NUM_INPUT_FIFOs-1:0] in_fifo_finished,
    //input AXI-Stream to FIFO interface 0
    input s_axis_fifo_0_aclk,
    input s_axis_fifo_0_aresetn,
    input s_axis_fifo_0_tlast,
    input s_axis_fifo_0_tvalid,
    input [S_AXIS_FIFO_0_DMWIDTH/8-1:0] s_axis_fifo_0_tkeep,
    input [S_AXIS_FIFO_0_DMWIDTH/8-1:0] s_axis_fifo_0_tstrb,
    input [S_AXIS_FIFO_0_DMWIDTH-1:0] s_axis_fifo_0_tdata,
    output s_axis_fifo_0_tready,
    output ap_fifo_iarg_0_empty_n,
    output [S_AXIS_FIFO_0_WIDTH-1:0] ap_fifo_iarg_0_dout,
    input ap_fifo_iarg_0_read,
    //input AXI-Stream to FIFO interface 1
    input s_axis_fifo_1_aclk,
    input s_axis_fifo_1_aresetn,
    input s_axis_fifo_1_tlast,
    input s_axis_fifo_1_tvalid,
    input [S_AXIS_FIFO_1_DMWIDTH/8-1:0] s_axis_fifo_1_tkeep,
    input [S_AXIS_FIFO_1_DMWIDTH/8-1:0] s_axis_fifo_1_tstrb,
    input [S_AXIS_FIFO_1_DMWIDTH-1:0] s_axis_fifo_1_tdata,
    output s_axis_fifo_1_tready,
    output ap_fifo_iarg_1_empty_n,
    output [S_AXIS_FIFO_1_WIDTH-1:0] ap_fifo_iarg_1_dout,
    input ap_fifo_iarg_1_read,
    //input AXI-Stream to FIFO interface 2
    input s_axis_fifo_2_aclk,
    input s_axis_fifo_2_aresetn,
    input s_axis_fifo_2_tlast,
    input s_axis_fifo_2_tvalid,
    input [S_AXIS_FIFO_2_DMWIDTH/8-1:0] s_axis_fifo_2_tkeep,
    input [S_AXIS_FIFO_2_DMWIDTH/8-1:0] s_axis_fifo_2_tstrb,
    input [S_AXIS_FIFO_2_DMWIDTH-1:0] s_axis_fifo_2_tdata,
    output s_axis_fifo_2_tready,
    output ap_fifo_iarg_2_empty_n,
    output [S_AXIS_FIFO_2_WIDTH-1:0] ap_fifo_iarg_2_dout,
    input ap_fifo_iarg_2_read,
    //input AXI-Stream to FIFO interface 3
    input s_axis_fifo_3_aclk,
    input s_axis_fifo_3_aresetn,
    input s_axis_fifo_3_tlast,
    input s_axis_fifo_3_tvalid,
    input [S_AXIS_FIFO_3_DMWIDTH/8-1:0] s_axis_fifo_3_tkeep,
    input [S_AXIS_FIFO_3_DMWIDTH/8-1:0] s_axis_fifo_3_tstrb,
    input [S_AXIS_FIFO_3_DMWIDTH-1:0] s_axis_fifo_3_tdata,
    output s_axis_fifo_3_tready,
    output ap_fifo_iarg_3_empty_n,
    output [S_AXIS_FIFO_3_WIDTH-1:0] ap_fifo_iarg_3_dout,
    input ap_fifo_iarg_3_read,
    //input AXI-Stream to FIFO interface 4
    input s_axis_fifo_4_aclk,
    input s_axis_fifo_4_aresetn,
    input s_axis_fifo_4_tlast,
    input s_axis_fifo_4_tvalid,
    input [S_AXIS_FIFO_4_DMWIDTH/8-1:0] s_axis_fifo_4_tkeep,
    input [S_AXIS_FIFO_4_DMWIDTH/8-1:0] s_axis_fifo_4_tstrb,
    input [S_AXIS_FIFO_4_DMWIDTH-1:0] s_axis_fifo_4_tdata,
    output s_axis_fifo_4_tready,
    output ap_fifo_iarg_4_empty_n,
    output [S_AXIS_FIFO_4_WIDTH-1:0] ap_fifo_iarg_4_dout,
    input ap_fifo_iarg_4_read,
    //input AXI-Stream to FIFO interface 5
    input s_axis_fifo_5_aclk,
    input s_axis_fifo_5_aresetn,
    input s_axis_fifo_5_tlast,
    input s_axis_fifo_5_tvalid,
    input [S_AXIS_FIFO_5_DMWIDTH/8-1:0] s_axis_fifo_5_tkeep,
    input [S_AXIS_FIFO_5_DMWIDTH/8-1:0] s_axis_fifo_5_tstrb,
    input [S_AXIS_FIFO_5_DMWIDTH-1:0] s_axis_fifo_5_tdata,
    output s_axis_fifo_5_tready,
    output ap_fifo_iarg_5_empty_n,
    output [S_AXIS_FIFO_5_WIDTH-1:0] ap_fifo_iarg_5_dout,
    input ap_fifo_iarg_5_read,
    //input AXI-Stream to FIFO interface 6
    input s_axis_fifo_6_aclk,
    input s_axis_fifo_6_aresetn,
    input s_axis_fifo_6_tlast,
    input s_axis_fifo_6_tvalid,
    input [S_AXIS_FIFO_6_DMWIDTH/8-1:0] s_axis_fifo_6_tkeep,
    input [S_AXIS_FIFO_6_DMWIDTH/8-1:0] s_axis_fifo_6_tstrb,
    input [S_AXIS_FIFO_6_DMWIDTH-1:0] s_axis_fifo_6_tdata,
    output s_axis_fifo_6_tready,
    output ap_fifo_iarg_6_empty_n,
    output [S_AXIS_FIFO_6_WIDTH-1:0] ap_fifo_iarg_6_dout,
    input ap_fifo_iarg_6_read,
    //input AXI-Stream to FIFO interface 7
    input s_axis_fifo_7_aclk,
    input s_axis_fifo_7_aresetn,
    input s_axis_fifo_7_tlast,
    input s_axis_fifo_7_tvalid,
    input [S_AXIS_FIFO_7_DMWIDTH/8-1:0] s_axis_fifo_7_tkeep,
    input [S_AXIS_FIFO_7_DMWIDTH/8-1:0] s_axis_fifo_7_tstrb,
    input [S_AXIS_FIFO_7_DMWIDTH-1:0] s_axis_fifo_7_tdata,
    output s_axis_fifo_7_tready,
    output ap_fifo_iarg_7_empty_n,
    output [S_AXIS_FIFO_7_WIDTH-1:0] ap_fifo_iarg_7_dout,
    input ap_fifo_iarg_7_read,
    //input AXI-Stream to FIFO interface 8
    input s_axis_fifo_8_aclk,
    input s_axis_fifo_8_aresetn,
    input s_axis_fifo_8_tlast,
    input s_axis_fifo_8_tvalid,
    input [S_AXIS_FIFO_8_DMWIDTH/8-1:0] s_axis_fifo_8_tkeep,
    input [S_AXIS_FIFO_8_DMWIDTH/8-1:0] s_axis_fifo_8_tstrb,
    input [S_AXIS_FIFO_8_DMWIDTH-1:0] s_axis_fifo_8_tdata,
    output s_axis_fifo_8_tready,
    output ap_fifo_iarg_8_empty_n,
    output [S_AXIS_FIFO_8_WIDTH-1:0] ap_fifo_iarg_8_dout,
    input ap_fifo_iarg_8_read,
    //input AXI-Stream to FIFO interface 9
    input s_axis_fifo_9_aclk,
    input s_axis_fifo_9_aresetn,
    input s_axis_fifo_9_tlast,
    input s_axis_fifo_9_tvalid,
    input [S_AXIS_FIFO_9_DMWIDTH/8-1:0] s_axis_fifo_9_tkeep,
    input [S_AXIS_FIFO_9_DMWIDTH/8-1:0] s_axis_fifo_9_tstrb,
    input [S_AXIS_FIFO_9_DMWIDTH-1:0] s_axis_fifo_9_tdata,
    output s_axis_fifo_9_tready,
    output ap_fifo_iarg_9_empty_n,
    output [S_AXIS_FIFO_9_WIDTH-1:0] ap_fifo_iarg_9_dout,
    input ap_fifo_iarg_9_read,
    //input AXI-Stream to FIFO interface 10
    input s_axis_fifo_10_aclk,
    input s_axis_fifo_10_aresetn,
    input s_axis_fifo_10_tlast,
    input s_axis_fifo_10_tvalid,
    input [S_AXIS_FIFO_10_DMWIDTH/8-1:0] s_axis_fifo_10_tkeep,
    input [S_AXIS_FIFO_10_DMWIDTH/8-1:0] s_axis_fifo_10_tstrb,
    input [S_AXIS_FIFO_10_DMWIDTH-1:0] s_axis_fifo_10_tdata,
    output s_axis_fifo_10_tready,
    output ap_fifo_iarg_10_empty_n,
    output [S_AXIS_FIFO_10_WIDTH-1:0] ap_fifo_iarg_10_dout,
    input ap_fifo_iarg_10_read,
    //input AXI-Stream to FIFO interface 11
    input s_axis_fifo_11_aclk,
    input s_axis_fifo_11_aresetn,
    input s_axis_fifo_11_tlast,
    input s_axis_fifo_11_tvalid,
    input [S_AXIS_FIFO_11_DMWIDTH/8-1:0] s_axis_fifo_11_tkeep,
    input [S_AXIS_FIFO_11_DMWIDTH/8-1:0] s_axis_fifo_11_tstrb,
    input [S_AXIS_FIFO_11_DMWIDTH-1:0] s_axis_fifo_11_tdata,
    output s_axis_fifo_11_tready,
    output ap_fifo_iarg_11_empty_n,
    output [S_AXIS_FIFO_11_WIDTH-1:0] ap_fifo_iarg_11_dout,
    input ap_fifo_iarg_11_read,
    //input AXI-Stream to FIFO interface 12
    input s_axis_fifo_12_aclk,
    input s_axis_fifo_12_aresetn,
    input s_axis_fifo_12_tlast,
    input s_axis_fifo_12_tvalid,
    input [S_AXIS_FIFO_12_DMWIDTH/8-1:0] s_axis_fifo_12_tkeep,
    input [S_AXIS_FIFO_12_DMWIDTH/8-1:0] s_axis_fifo_12_tstrb,
    input [S_AXIS_FIFO_12_DMWIDTH-1:0] s_axis_fifo_12_tdata,
    output s_axis_fifo_12_tready,
    output ap_fifo_iarg_12_empty_n,
    output [S_AXIS_FIFO_12_WIDTH-1:0] ap_fifo_iarg_12_dout,
    input ap_fifo_iarg_12_read,
    //input AXI-Stream to FIFO interface 13
    input s_axis_fifo_13_aclk,
    input s_axis_fifo_13_aresetn,
    input s_axis_fifo_13_tlast,
    input s_axis_fifo_13_tvalid,
    input [S_AXIS_FIFO_13_DMWIDTH/8-1:0] s_axis_fifo_13_tkeep,
    input [S_AXIS_FIFO_13_DMWIDTH/8-1:0] s_axis_fifo_13_tstrb,
    input [S_AXIS_FIFO_13_DMWIDTH-1:0] s_axis_fifo_13_tdata,
    output s_axis_fifo_13_tready,
    output ap_fifo_iarg_13_empty_n,
    output [S_AXIS_FIFO_13_WIDTH-1:0] ap_fifo_iarg_13_dout,
    input ap_fifo_iarg_13_read,
    //input AXI-Stream to FIFO interface 14
    input s_axis_fifo_14_aclk,
    input s_axis_fifo_14_aresetn,
    input s_axis_fifo_14_tlast,
    input s_axis_fifo_14_tvalid,
    input [S_AXIS_FIFO_14_DMWIDTH/8-1:0] s_axis_fifo_14_tkeep,
    input [S_AXIS_FIFO_14_DMWIDTH/8-1:0] s_axis_fifo_14_tstrb,
    input [S_AXIS_FIFO_14_DMWIDTH-1:0] s_axis_fifo_14_tdata,
    output s_axis_fifo_14_tready,
    output ap_fifo_iarg_14_empty_n,
    output [S_AXIS_FIFO_14_WIDTH-1:0] ap_fifo_iarg_14_dout,
    input ap_fifo_iarg_14_read,
    //input AXI-Stream to FIFO interface 15
    input s_axis_fifo_15_aclk,
    input s_axis_fifo_15_aresetn,
    input s_axis_fifo_15_tlast,
    input s_axis_fifo_15_tvalid,
    input [S_AXIS_FIFO_15_DMWIDTH/8-1:0] s_axis_fifo_15_tkeep,
    input [S_AXIS_FIFO_15_DMWIDTH/8-1:0] s_axis_fifo_15_tstrb,
    input [S_AXIS_FIFO_15_DMWIDTH-1:0] s_axis_fifo_15_tdata,
    output s_axis_fifo_15_tready,
    output ap_fifo_iarg_15_empty_n,
    output [S_AXIS_FIFO_15_WIDTH-1:0] ap_fifo_iarg_15_dout,
    input ap_fifo_iarg_15_read,
    //input AXI-Stream to FIFO interface 16
    input s_axis_fifo_16_aclk,
    input s_axis_fifo_16_aresetn,
    input s_axis_fifo_16_tlast,
    input s_axis_fifo_16_tvalid,
    input [S_AXIS_FIFO_16_DMWIDTH/8-1:0] s_axis_fifo_16_tkeep,
    input [S_AXIS_FIFO_16_DMWIDTH/8-1:0] s_axis_fifo_16_tstrb,
    input [S_AXIS_FIFO_16_DMWIDTH-1:0] s_axis_fifo_16_tdata,
    output s_axis_fifo_16_tready,
    output ap_fifo_iarg_16_empty_n,
    output [S_AXIS_FIFO_16_WIDTH-1:0] ap_fifo_iarg_16_dout,
    input ap_fifo_iarg_16_read,
    //input AXI-Stream to FIFO interface 17
    input s_axis_fifo_17_aclk,
    input s_axis_fifo_17_aresetn,
    input s_axis_fifo_17_tlast,
    input s_axis_fifo_17_tvalid,
    input [S_AXIS_FIFO_17_DMWIDTH/8-1:0] s_axis_fifo_17_tkeep,
    input [S_AXIS_FIFO_17_DMWIDTH/8-1:0] s_axis_fifo_17_tstrb,
    input [S_AXIS_FIFO_17_DMWIDTH-1:0] s_axis_fifo_17_tdata,
    output s_axis_fifo_17_tready,
    output ap_fifo_iarg_17_empty_n,
    output [S_AXIS_FIFO_17_WIDTH-1:0] ap_fifo_iarg_17_dout,
    input ap_fifo_iarg_17_read,
    //input AXI-Stream to FIFO interface 18
    input s_axis_fifo_18_aclk,
    input s_axis_fifo_18_aresetn,
    input s_axis_fifo_18_tlast,
    input s_axis_fifo_18_tvalid,
    input [S_AXIS_FIFO_18_DMWIDTH/8-1:0] s_axis_fifo_18_tkeep,
    input [S_AXIS_FIFO_18_DMWIDTH/8-1:0] s_axis_fifo_18_tstrb,
    input [S_AXIS_FIFO_18_DMWIDTH-1:0] s_axis_fifo_18_tdata,
    output s_axis_fifo_18_tready,
    output ap_fifo_iarg_18_empty_n,
    output [S_AXIS_FIFO_18_WIDTH-1:0] ap_fifo_iarg_18_dout,
    input ap_fifo_iarg_18_read,
    //input AXI-Stream to FIFO interface 19
    input s_axis_fifo_19_aclk,
    input s_axis_fifo_19_aresetn,
    input s_axis_fifo_19_tlast,
    input s_axis_fifo_19_tvalid,
    input [S_AXIS_FIFO_19_DMWIDTH/8-1:0] s_axis_fifo_19_tkeep,
    input [S_AXIS_FIFO_19_DMWIDTH/8-1:0] s_axis_fifo_19_tstrb,
    input [S_AXIS_FIFO_19_DMWIDTH-1:0] s_axis_fifo_19_tdata,
    output s_axis_fifo_19_tready,
    output ap_fifo_iarg_19_empty_n,
    output [S_AXIS_FIFO_19_WIDTH-1:0] ap_fifo_iarg_19_dout,
    input ap_fifo_iarg_19_read,
    //input AXI-Stream to FIFO interface 20
    input s_axis_fifo_20_aclk,
    input s_axis_fifo_20_aresetn,
    input s_axis_fifo_20_tlast,
    input s_axis_fifo_20_tvalid,
    input [S_AXIS_FIFO_20_DMWIDTH/8-1:0] s_axis_fifo_20_tkeep,
    input [S_AXIS_FIFO_20_DMWIDTH/8-1:0] s_axis_fifo_20_tstrb,
    input [S_AXIS_FIFO_20_DMWIDTH-1:0] s_axis_fifo_20_tdata,
    output s_axis_fifo_20_tready,
    output ap_fifo_iarg_20_empty_n,
    output [S_AXIS_FIFO_20_WIDTH-1:0] ap_fifo_iarg_20_dout,
    input ap_fifo_iarg_20_read,
    //input AXI-Stream to FIFO interface 21
    input s_axis_fifo_21_aclk,
    input s_axis_fifo_21_aresetn,
    input s_axis_fifo_21_tlast,
    input s_axis_fifo_21_tvalid,
    input [S_AXIS_FIFO_21_DMWIDTH/8-1:0] s_axis_fifo_21_tkeep,
    input [S_AXIS_FIFO_21_DMWIDTH/8-1:0] s_axis_fifo_21_tstrb,
    input [S_AXIS_FIFO_21_DMWIDTH-1:0] s_axis_fifo_21_tdata,
    output s_axis_fifo_21_tready,
    output ap_fifo_iarg_21_empty_n,
    output [S_AXIS_FIFO_21_WIDTH-1:0] ap_fifo_iarg_21_dout,
    input ap_fifo_iarg_21_read,
    //input AXI-Stream to FIFO interface 22
    input s_axis_fifo_22_aclk,
    input s_axis_fifo_22_aresetn,
    input s_axis_fifo_22_tlast,
    input s_axis_fifo_22_tvalid,
    input [S_AXIS_FIFO_22_DMWIDTH/8-1:0] s_axis_fifo_22_tkeep,
    input [S_AXIS_FIFO_22_DMWIDTH/8-1:0] s_axis_fifo_22_tstrb,
    input [S_AXIS_FIFO_22_DMWIDTH-1:0] s_axis_fifo_22_tdata,
    output s_axis_fifo_22_tready,
    output ap_fifo_iarg_22_empty_n,
    output [S_AXIS_FIFO_22_WIDTH-1:0] ap_fifo_iarg_22_dout,
    input ap_fifo_iarg_22_read,
    //input AXI-Stream to FIFO interface 23
    input s_axis_fifo_23_aclk,
    input s_axis_fifo_23_aresetn,
    input s_axis_fifo_23_tlast,
    input s_axis_fifo_23_tvalid,
    input [S_AXIS_FIFO_23_DMWIDTH/8-1:0] s_axis_fifo_23_tkeep,
    input [S_AXIS_FIFO_23_DMWIDTH/8-1:0] s_axis_fifo_23_tstrb,
    input [S_AXIS_FIFO_23_DMWIDTH-1:0] s_axis_fifo_23_tdata,
    output s_axis_fifo_23_tready,
    output ap_fifo_iarg_23_empty_n,
    output [S_AXIS_FIFO_23_WIDTH-1:0] ap_fifo_iarg_23_dout,
    input ap_fifo_iarg_23_read,
    //input AXI-Stream to FIFO interface 24
    input s_axis_fifo_24_aclk,
    input s_axis_fifo_24_aresetn,
    input s_axis_fifo_24_tlast,
    input s_axis_fifo_24_tvalid,
    input [S_AXIS_FIFO_24_DMWIDTH/8-1:0] s_axis_fifo_24_tkeep,
    input [S_AXIS_FIFO_24_DMWIDTH/8-1:0] s_axis_fifo_24_tstrb,
    input [S_AXIS_FIFO_24_DMWIDTH-1:0] s_axis_fifo_24_tdata,
    output s_axis_fifo_24_tready,
    output ap_fifo_iarg_24_empty_n,
    output [S_AXIS_FIFO_24_WIDTH-1:0] ap_fifo_iarg_24_dout,
    input ap_fifo_iarg_24_read,
    //input AXI-Stream to FIFO interface 25
    input s_axis_fifo_25_aclk,
    input s_axis_fifo_25_aresetn,
    input s_axis_fifo_25_tlast,
    input s_axis_fifo_25_tvalid,
    input [S_AXIS_FIFO_25_DMWIDTH/8-1:0] s_axis_fifo_25_tkeep,
    input [S_AXIS_FIFO_25_DMWIDTH/8-1:0] s_axis_fifo_25_tstrb,
    input [S_AXIS_FIFO_25_DMWIDTH-1:0] s_axis_fifo_25_tdata,
    output s_axis_fifo_25_tready,
    output ap_fifo_iarg_25_empty_n,
    output [S_AXIS_FIFO_25_WIDTH-1:0] ap_fifo_iarg_25_dout,
    input ap_fifo_iarg_25_read,
    //input AXI-Stream to FIFO interface 26
    input s_axis_fifo_26_aclk,
    input s_axis_fifo_26_aresetn,
    input s_axis_fifo_26_tlast,
    input s_axis_fifo_26_tvalid,
    input [S_AXIS_FIFO_26_DMWIDTH/8-1:0] s_axis_fifo_26_tkeep,
    input [S_AXIS_FIFO_26_DMWIDTH/8-1:0] s_axis_fifo_26_tstrb,
    input [S_AXIS_FIFO_26_DMWIDTH-1:0] s_axis_fifo_26_tdata,
    output s_axis_fifo_26_tready,
    output ap_fifo_iarg_26_empty_n,
    output [S_AXIS_FIFO_26_WIDTH-1:0] ap_fifo_iarg_26_dout,
    input ap_fifo_iarg_26_read,
    //input AXI-Stream to FIFO interface 27
    input s_axis_fifo_27_aclk,
    input s_axis_fifo_27_aresetn,
    input s_axis_fifo_27_tlast,
    input s_axis_fifo_27_tvalid,
    input [S_AXIS_FIFO_27_DMWIDTH/8-1:0] s_axis_fifo_27_tkeep,
    input [S_AXIS_FIFO_27_DMWIDTH/8-1:0] s_axis_fifo_27_tstrb,
    input [S_AXIS_FIFO_27_DMWIDTH-1:0] s_axis_fifo_27_tdata,
    output s_axis_fifo_27_tready,
    output ap_fifo_iarg_27_empty_n,
    output [S_AXIS_FIFO_27_WIDTH-1:0] ap_fifo_iarg_27_dout,
    input ap_fifo_iarg_27_read,
    //input AXI-Stream to FIFO interface 28
    input s_axis_fifo_28_aclk,
    input s_axis_fifo_28_aresetn,
    input s_axis_fifo_28_tlast,
    input s_axis_fifo_28_tvalid,
    input [S_AXIS_FIFO_28_DMWIDTH/8-1:0] s_axis_fifo_28_tkeep,
    input [S_AXIS_FIFO_28_DMWIDTH/8-1:0] s_axis_fifo_28_tstrb,
    input [S_AXIS_FIFO_28_DMWIDTH-1:0] s_axis_fifo_28_tdata,
    output s_axis_fifo_28_tready,
    output ap_fifo_iarg_28_empty_n,
    output [S_AXIS_FIFO_28_WIDTH-1:0] ap_fifo_iarg_28_dout,
    input ap_fifo_iarg_28_read,
    //input AXI-Stream to FIFO interface 29
    input s_axis_fifo_29_aclk,
    input s_axis_fifo_29_aresetn,
    input s_axis_fifo_29_tlast,
    input s_axis_fifo_29_tvalid,
    input [S_AXIS_FIFO_29_DMWIDTH/8-1:0] s_axis_fifo_29_tkeep,
    input [S_AXIS_FIFO_29_DMWIDTH/8-1:0] s_axis_fifo_29_tstrb,
    input [S_AXIS_FIFO_29_DMWIDTH-1:0] s_axis_fifo_29_tdata,
    output s_axis_fifo_29_tready,
    output ap_fifo_iarg_29_empty_n,
    output [S_AXIS_FIFO_29_WIDTH-1:0] ap_fifo_iarg_29_dout,
    input ap_fifo_iarg_29_read,
    //input AXI-Stream to FIFO interface 30
    input s_axis_fifo_30_aclk,
    input s_axis_fifo_30_aresetn,
    input s_axis_fifo_30_tlast,
    input s_axis_fifo_30_tvalid,
    input [S_AXIS_FIFO_30_DMWIDTH/8-1:0] s_axis_fifo_30_tkeep,
    input [S_AXIS_FIFO_30_DMWIDTH/8-1:0] s_axis_fifo_30_tstrb,
    input [S_AXIS_FIFO_30_DMWIDTH-1:0] s_axis_fifo_30_tdata,
    output s_axis_fifo_30_tready,
    output ap_fifo_iarg_30_empty_n,
    output [S_AXIS_FIFO_30_WIDTH-1:0] ap_fifo_iarg_30_dout,
    input ap_fifo_iarg_30_read,
    //input AXI-Stream to FIFO interface 31
    input s_axis_fifo_31_aclk,
    input s_axis_fifo_31_aresetn,
    input s_axis_fifo_31_tlast,
    input s_axis_fifo_31_tvalid,
    input [S_AXIS_FIFO_31_DMWIDTH/8-1:0] s_axis_fifo_31_tkeep,
    input [S_AXIS_FIFO_31_DMWIDTH/8-1:0] s_axis_fifo_31_tstrb,
    input [S_AXIS_FIFO_31_DMWIDTH-1:0] s_axis_fifo_31_tdata,
    output s_axis_fifo_31_tready,
    output ap_fifo_iarg_31_empty_n,
    output [S_AXIS_FIFO_31_WIDTH-1:0] ap_fifo_iarg_31_dout,
    input ap_fifo_iarg_31_read,
    //input AXI-Stream to FIFO interface 32
    input s_axis_fifo_32_aclk,
    input s_axis_fifo_32_aresetn,
    input s_axis_fifo_32_tlast,
    input s_axis_fifo_32_tvalid,
    input [S_AXIS_FIFO_32_DMWIDTH/8-1:0] s_axis_fifo_32_tkeep,
    input [S_AXIS_FIFO_32_DMWIDTH/8-1:0] s_axis_fifo_32_tstrb,
    input [S_AXIS_FIFO_32_DMWIDTH-1:0] s_axis_fifo_32_tdata,
    output s_axis_fifo_32_tready,
    output ap_fifo_iarg_32_empty_n,
    output [S_AXIS_FIFO_32_WIDTH-1:0] ap_fifo_iarg_32_dout,
    input ap_fifo_iarg_32_read,
    //input AXI-Stream to FIFO interface 33
    input s_axis_fifo_33_aclk,
    input s_axis_fifo_33_aresetn,
    input s_axis_fifo_33_tlast,
    input s_axis_fifo_33_tvalid,
    input [S_AXIS_FIFO_33_DMWIDTH/8-1:0] s_axis_fifo_33_tkeep,
    input [S_AXIS_FIFO_33_DMWIDTH/8-1:0] s_axis_fifo_33_tstrb,
    input [S_AXIS_FIFO_33_DMWIDTH-1:0] s_axis_fifo_33_tdata,
    output s_axis_fifo_33_tready,
    output ap_fifo_iarg_33_empty_n,
    output [S_AXIS_FIFO_33_WIDTH-1:0] ap_fifo_iarg_33_dout,
    input ap_fifo_iarg_33_read,
    //input AXI-Stream to FIFO interface 34
    input s_axis_fifo_34_aclk,
    input s_axis_fifo_34_aresetn,
    input s_axis_fifo_34_tlast,
    input s_axis_fifo_34_tvalid,
    input [S_AXIS_FIFO_34_DMWIDTH/8-1:0] s_axis_fifo_34_tkeep,
    input [S_AXIS_FIFO_34_DMWIDTH/8-1:0] s_axis_fifo_34_tstrb,
    input [S_AXIS_FIFO_34_DMWIDTH-1:0] s_axis_fifo_34_tdata,
    output s_axis_fifo_34_tready,
    output ap_fifo_iarg_34_empty_n,
    output [S_AXIS_FIFO_34_WIDTH-1:0] ap_fifo_iarg_34_dout,
    input ap_fifo_iarg_34_read,
    //input AXI-Stream to FIFO interface 35
    input s_axis_fifo_35_aclk,
    input s_axis_fifo_35_aresetn,
    input s_axis_fifo_35_tlast,
    input s_axis_fifo_35_tvalid,
    input [S_AXIS_FIFO_35_DMWIDTH/8-1:0] s_axis_fifo_35_tkeep,
    input [S_AXIS_FIFO_35_DMWIDTH/8-1:0] s_axis_fifo_35_tstrb,
    input [S_AXIS_FIFO_35_DMWIDTH-1:0] s_axis_fifo_35_tdata,
    output s_axis_fifo_35_tready,
    output ap_fifo_iarg_35_empty_n,
    output [S_AXIS_FIFO_35_WIDTH-1:0] ap_fifo_iarg_35_dout,
    input ap_fifo_iarg_35_read,
    //input AXI-Stream to FIFO interface 36
    input s_axis_fifo_36_aclk,
    input s_axis_fifo_36_aresetn,
    input s_axis_fifo_36_tlast,
    input s_axis_fifo_36_tvalid,
    input [S_AXIS_FIFO_36_DMWIDTH/8-1:0] s_axis_fifo_36_tkeep,
    input [S_AXIS_FIFO_36_DMWIDTH/8-1:0] s_axis_fifo_36_tstrb,
    input [S_AXIS_FIFO_36_DMWIDTH-1:0] s_axis_fifo_36_tdata,
    output s_axis_fifo_36_tready,
    output ap_fifo_iarg_36_empty_n,
    output [S_AXIS_FIFO_36_WIDTH-1:0] ap_fifo_iarg_36_dout,
    input ap_fifo_iarg_36_read,
    //input AXI-Stream to FIFO interface 37
    input s_axis_fifo_37_aclk,
    input s_axis_fifo_37_aresetn,
    input s_axis_fifo_37_tlast,
    input s_axis_fifo_37_tvalid,
    input [S_AXIS_FIFO_37_DMWIDTH/8-1:0] s_axis_fifo_37_tkeep,
    input [S_AXIS_FIFO_37_DMWIDTH/8-1:0] s_axis_fifo_37_tstrb,
    input [S_AXIS_FIFO_37_DMWIDTH-1:0] s_axis_fifo_37_tdata,
    output s_axis_fifo_37_tready,
    output ap_fifo_iarg_37_empty_n,
    output [S_AXIS_FIFO_37_WIDTH-1:0] ap_fifo_iarg_37_dout,
    input ap_fifo_iarg_37_read,
    //input AXI-Stream to FIFO interface 38
    input s_axis_fifo_38_aclk,
    input s_axis_fifo_38_aresetn,
    input s_axis_fifo_38_tlast,
    input s_axis_fifo_38_tvalid,
    input [S_AXIS_FIFO_38_DMWIDTH/8-1:0] s_axis_fifo_38_tkeep,
    input [S_AXIS_FIFO_38_DMWIDTH/8-1:0] s_axis_fifo_38_tstrb,
    input [S_AXIS_FIFO_38_DMWIDTH-1:0] s_axis_fifo_38_tdata,
    output s_axis_fifo_38_tready,
    output ap_fifo_iarg_38_empty_n,
    output [S_AXIS_FIFO_38_WIDTH-1:0] ap_fifo_iarg_38_dout,
    input ap_fifo_iarg_38_read,
    //input AXI-Stream to FIFO interface 39
    input s_axis_fifo_39_aclk,
    input s_axis_fifo_39_aresetn,
    input s_axis_fifo_39_tlast,
    input s_axis_fifo_39_tvalid,
    input [S_AXIS_FIFO_39_DMWIDTH/8-1:0] s_axis_fifo_39_tkeep,
    input [S_AXIS_FIFO_39_DMWIDTH/8-1:0] s_axis_fifo_39_tstrb,
    input [S_AXIS_FIFO_39_DMWIDTH-1:0] s_axis_fifo_39_tdata,
    output s_axis_fifo_39_tready,
    output ap_fifo_iarg_39_empty_n,
    output [S_AXIS_FIFO_39_WIDTH-1:0] ap_fifo_iarg_39_dout,
    input ap_fifo_iarg_39_read,
    //input AXI-Stream to FIFO interface 40
    input s_axis_fifo_40_aclk,
    input s_axis_fifo_40_aresetn,
    input s_axis_fifo_40_tlast,
    input s_axis_fifo_40_tvalid,
    input [S_AXIS_FIFO_40_DMWIDTH/8-1:0] s_axis_fifo_40_tkeep,
    input [S_AXIS_FIFO_40_DMWIDTH/8-1:0] s_axis_fifo_40_tstrb,
    input [S_AXIS_FIFO_40_DMWIDTH-1:0] s_axis_fifo_40_tdata,
    output s_axis_fifo_40_tready,
    output ap_fifo_iarg_40_empty_n,
    output [S_AXIS_FIFO_40_WIDTH-1:0] ap_fifo_iarg_40_dout,
    input ap_fifo_iarg_40_read,
    //input AXI-Stream to FIFO interface 41
    input s_axis_fifo_41_aclk,
    input s_axis_fifo_41_aresetn,
    input s_axis_fifo_41_tlast,
    input s_axis_fifo_41_tvalid,
    input [S_AXIS_FIFO_41_DMWIDTH/8-1:0] s_axis_fifo_41_tkeep,
    input [S_AXIS_FIFO_41_DMWIDTH/8-1:0] s_axis_fifo_41_tstrb,
    input [S_AXIS_FIFO_41_DMWIDTH-1:0] s_axis_fifo_41_tdata,
    output s_axis_fifo_41_tready,
    output ap_fifo_iarg_41_empty_n,
    output [S_AXIS_FIFO_41_WIDTH-1:0] ap_fifo_iarg_41_dout,
    input ap_fifo_iarg_41_read,
    //input AXI-Stream to FIFO interface 42
    input s_axis_fifo_42_aclk,
    input s_axis_fifo_42_aresetn,
    input s_axis_fifo_42_tlast,
    input s_axis_fifo_42_tvalid,
    input [S_AXIS_FIFO_42_DMWIDTH/8-1:0] s_axis_fifo_42_tkeep,
    input [S_AXIS_FIFO_42_DMWIDTH/8-1:0] s_axis_fifo_42_tstrb,
    input [S_AXIS_FIFO_42_DMWIDTH-1:0] s_axis_fifo_42_tdata,
    output s_axis_fifo_42_tready,
    output ap_fifo_iarg_42_empty_n,
    output [S_AXIS_FIFO_42_WIDTH-1:0] ap_fifo_iarg_42_dout,
    input ap_fifo_iarg_42_read,
    //input AXI-Stream to FIFO interface 43
    input s_axis_fifo_43_aclk,
    input s_axis_fifo_43_aresetn,
    input s_axis_fifo_43_tlast,
    input s_axis_fifo_43_tvalid,
    input [S_AXIS_FIFO_43_DMWIDTH/8-1:0] s_axis_fifo_43_tkeep,
    input [S_AXIS_FIFO_43_DMWIDTH/8-1:0] s_axis_fifo_43_tstrb,
    input [S_AXIS_FIFO_43_DMWIDTH-1:0] s_axis_fifo_43_tdata,
    output s_axis_fifo_43_tready,
    output ap_fifo_iarg_43_empty_n,
    output [S_AXIS_FIFO_43_WIDTH-1:0] ap_fifo_iarg_43_dout,
    input ap_fifo_iarg_43_read,
    //input AXI-Stream to FIFO interface 44
    input s_axis_fifo_44_aclk,
    input s_axis_fifo_44_aresetn,
    input s_axis_fifo_44_tlast,
    input s_axis_fifo_44_tvalid,
    input [S_AXIS_FIFO_44_DMWIDTH/8-1:0] s_axis_fifo_44_tkeep,
    input [S_AXIS_FIFO_44_DMWIDTH/8-1:0] s_axis_fifo_44_tstrb,
    input [S_AXIS_FIFO_44_DMWIDTH-1:0] s_axis_fifo_44_tdata,
    output s_axis_fifo_44_tready,
    output ap_fifo_iarg_44_empty_n,
    output [S_AXIS_FIFO_44_WIDTH-1:0] ap_fifo_iarg_44_dout,
    input ap_fifo_iarg_44_read,
    //input AXI-Stream to FIFO interface 45
    input s_axis_fifo_45_aclk,
    input s_axis_fifo_45_aresetn,
    input s_axis_fifo_45_tlast,
    input s_axis_fifo_45_tvalid,
    input [S_AXIS_FIFO_45_DMWIDTH/8-1:0] s_axis_fifo_45_tkeep,
    input [S_AXIS_FIFO_45_DMWIDTH/8-1:0] s_axis_fifo_45_tstrb,
    input [S_AXIS_FIFO_45_DMWIDTH-1:0] s_axis_fifo_45_tdata,
    output s_axis_fifo_45_tready,
    output ap_fifo_iarg_45_empty_n,
    output [S_AXIS_FIFO_45_WIDTH-1:0] ap_fifo_iarg_45_dout,
    input ap_fifo_iarg_45_read,
    //input AXI-Stream to FIFO interface 46
    input s_axis_fifo_46_aclk,
    input s_axis_fifo_46_aresetn,
    input s_axis_fifo_46_tlast,
    input s_axis_fifo_46_tvalid,
    input [S_AXIS_FIFO_46_DMWIDTH/8-1:0] s_axis_fifo_46_tkeep,
    input [S_AXIS_FIFO_46_DMWIDTH/8-1:0] s_axis_fifo_46_tstrb,
    input [S_AXIS_FIFO_46_DMWIDTH-1:0] s_axis_fifo_46_tdata,
    output s_axis_fifo_46_tready,
    output ap_fifo_iarg_46_empty_n,
    output [S_AXIS_FIFO_46_WIDTH-1:0] ap_fifo_iarg_46_dout,
    input ap_fifo_iarg_46_read,
    //input AXI-Stream to FIFO interface 47
    input s_axis_fifo_47_aclk,
    input s_axis_fifo_47_aresetn,
    input s_axis_fifo_47_tlast,
    input s_axis_fifo_47_tvalid,
    input [S_AXIS_FIFO_47_DMWIDTH/8-1:0] s_axis_fifo_47_tkeep,
    input [S_AXIS_FIFO_47_DMWIDTH/8-1:0] s_axis_fifo_47_tstrb,
    input [S_AXIS_FIFO_47_DMWIDTH-1:0] s_axis_fifo_47_tdata,
    output s_axis_fifo_47_tready,
    output ap_fifo_iarg_47_empty_n,
    output [S_AXIS_FIFO_47_WIDTH-1:0] ap_fifo_iarg_47_dout,
    input ap_fifo_iarg_47_read,
    //input AXI-Stream to FIFO interface 48
    input s_axis_fifo_48_aclk,
    input s_axis_fifo_48_aresetn,
    input s_axis_fifo_48_tlast,
    input s_axis_fifo_48_tvalid,
    input [S_AXIS_FIFO_48_DMWIDTH/8-1:0] s_axis_fifo_48_tkeep,
    input [S_AXIS_FIFO_48_DMWIDTH/8-1:0] s_axis_fifo_48_tstrb,
    input [S_AXIS_FIFO_48_DMWIDTH-1:0] s_axis_fifo_48_tdata,
    output s_axis_fifo_48_tready,
    output ap_fifo_iarg_48_empty_n,
    output [S_AXIS_FIFO_48_WIDTH-1:0] ap_fifo_iarg_48_dout,
    input ap_fifo_iarg_48_read,
    //input AXI-Stream to FIFO interface 49
    input s_axis_fifo_49_aclk,
    input s_axis_fifo_49_aresetn,
    input s_axis_fifo_49_tlast,
    input s_axis_fifo_49_tvalid,
    input [S_AXIS_FIFO_49_DMWIDTH/8-1:0] s_axis_fifo_49_tkeep,
    input [S_AXIS_FIFO_49_DMWIDTH/8-1:0] s_axis_fifo_49_tstrb,
    input [S_AXIS_FIFO_49_DMWIDTH-1:0] s_axis_fifo_49_tdata,
    output s_axis_fifo_49_tready,
    output ap_fifo_iarg_49_empty_n,
    output [S_AXIS_FIFO_49_WIDTH-1:0] ap_fifo_iarg_49_dout,
    input ap_fifo_iarg_49_read,
    //input AXI-Stream to FIFO interface 50
    input s_axis_fifo_50_aclk,
    input s_axis_fifo_50_aresetn,
    input s_axis_fifo_50_tlast,
    input s_axis_fifo_50_tvalid,
    input [S_AXIS_FIFO_50_DMWIDTH/8-1:0] s_axis_fifo_50_tkeep,
    input [S_AXIS_FIFO_50_DMWIDTH/8-1:0] s_axis_fifo_50_tstrb,
    input [S_AXIS_FIFO_50_DMWIDTH-1:0] s_axis_fifo_50_tdata,
    output s_axis_fifo_50_tready,
    output ap_fifo_iarg_50_empty_n,
    output [S_AXIS_FIFO_50_WIDTH-1:0] ap_fifo_iarg_50_dout,
    input ap_fifo_iarg_50_read,
    //input AXI-Stream to FIFO interface 51
    input s_axis_fifo_51_aclk,
    input s_axis_fifo_51_aresetn,
    input s_axis_fifo_51_tlast,
    input s_axis_fifo_51_tvalid,
    input [S_AXIS_FIFO_51_DMWIDTH/8-1:0] s_axis_fifo_51_tkeep,
    input [S_AXIS_FIFO_51_DMWIDTH/8-1:0] s_axis_fifo_51_tstrb,
    input [S_AXIS_FIFO_51_DMWIDTH-1:0] s_axis_fifo_51_tdata,
    output s_axis_fifo_51_tready,
    output ap_fifo_iarg_51_empty_n,
    output [S_AXIS_FIFO_51_WIDTH-1:0] ap_fifo_iarg_51_dout,
    input ap_fifo_iarg_51_read,
    //input AXI-Stream to FIFO interface 52
    input s_axis_fifo_52_aclk,
    input s_axis_fifo_52_aresetn,
    input s_axis_fifo_52_tlast,
    input s_axis_fifo_52_tvalid,
    input [S_AXIS_FIFO_52_DMWIDTH/8-1:0] s_axis_fifo_52_tkeep,
    input [S_AXIS_FIFO_52_DMWIDTH/8-1:0] s_axis_fifo_52_tstrb,
    input [S_AXIS_FIFO_52_DMWIDTH-1:0] s_axis_fifo_52_tdata,
    output s_axis_fifo_52_tready,
    output ap_fifo_iarg_52_empty_n,
    output [S_AXIS_FIFO_52_WIDTH-1:0] ap_fifo_iarg_52_dout,
    input ap_fifo_iarg_52_read,
    //input AXI-Stream to FIFO interface 53
    input s_axis_fifo_53_aclk,
    input s_axis_fifo_53_aresetn,
    input s_axis_fifo_53_tlast,
    input s_axis_fifo_53_tvalid,
    input [S_AXIS_FIFO_53_DMWIDTH/8-1:0] s_axis_fifo_53_tkeep,
    input [S_AXIS_FIFO_53_DMWIDTH/8-1:0] s_axis_fifo_53_tstrb,
    input [S_AXIS_FIFO_53_DMWIDTH-1:0] s_axis_fifo_53_tdata,
    output s_axis_fifo_53_tready,
    output ap_fifo_iarg_53_empty_n,
    output [S_AXIS_FIFO_53_WIDTH-1:0] ap_fifo_iarg_53_dout,
    input ap_fifo_iarg_53_read,
    //input AXI-Stream to FIFO interface 54
    input s_axis_fifo_54_aclk,
    input s_axis_fifo_54_aresetn,
    input s_axis_fifo_54_tlast,
    input s_axis_fifo_54_tvalid,
    input [S_AXIS_FIFO_54_DMWIDTH/8-1:0] s_axis_fifo_54_tkeep,
    input [S_AXIS_FIFO_54_DMWIDTH/8-1:0] s_axis_fifo_54_tstrb,
    input [S_AXIS_FIFO_54_DMWIDTH-1:0] s_axis_fifo_54_tdata,
    output s_axis_fifo_54_tready,
    output ap_fifo_iarg_54_empty_n,
    output [S_AXIS_FIFO_54_WIDTH-1:0] ap_fifo_iarg_54_dout,
    input ap_fifo_iarg_54_read,
    //input AXI-Stream to FIFO interface 55
    input s_axis_fifo_55_aclk,
    input s_axis_fifo_55_aresetn,
    input s_axis_fifo_55_tlast,
    input s_axis_fifo_55_tvalid,
    input [S_AXIS_FIFO_55_DMWIDTH/8-1:0] s_axis_fifo_55_tkeep,
    input [S_AXIS_FIFO_55_DMWIDTH/8-1:0] s_axis_fifo_55_tstrb,
    input [S_AXIS_FIFO_55_DMWIDTH-1:0] s_axis_fifo_55_tdata,
    output s_axis_fifo_55_tready,
    output ap_fifo_iarg_55_empty_n,
    output [S_AXIS_FIFO_55_WIDTH-1:0] ap_fifo_iarg_55_dout,
    input ap_fifo_iarg_55_read,
    //input AXI-Stream to FIFO interface 56
    input s_axis_fifo_56_aclk,
    input s_axis_fifo_56_aresetn,
    input s_axis_fifo_56_tlast,
    input s_axis_fifo_56_tvalid,
    input [S_AXIS_FIFO_56_DMWIDTH/8-1:0] s_axis_fifo_56_tkeep,
    input [S_AXIS_FIFO_56_DMWIDTH/8-1:0] s_axis_fifo_56_tstrb,
    input [S_AXIS_FIFO_56_DMWIDTH-1:0] s_axis_fifo_56_tdata,
    output s_axis_fifo_56_tready,
    output ap_fifo_iarg_56_empty_n,
    output [S_AXIS_FIFO_56_WIDTH-1:0] ap_fifo_iarg_56_dout,
    input ap_fifo_iarg_56_read,
    //input AXI-Stream to FIFO interface 57
    input s_axis_fifo_57_aclk,
    input s_axis_fifo_57_aresetn,
    input s_axis_fifo_57_tlast,
    input s_axis_fifo_57_tvalid,
    input [S_AXIS_FIFO_57_DMWIDTH/8-1:0] s_axis_fifo_57_tkeep,
    input [S_AXIS_FIFO_57_DMWIDTH/8-1:0] s_axis_fifo_57_tstrb,
    input [S_AXIS_FIFO_57_DMWIDTH-1:0] s_axis_fifo_57_tdata,
    output s_axis_fifo_57_tready,
    output ap_fifo_iarg_57_empty_n,
    output [S_AXIS_FIFO_57_WIDTH-1:0] ap_fifo_iarg_57_dout,
    input ap_fifo_iarg_57_read,
    //input AXI-Stream to FIFO interface 58
    input s_axis_fifo_58_aclk,
    input s_axis_fifo_58_aresetn,
    input s_axis_fifo_58_tlast,
    input s_axis_fifo_58_tvalid,
    input [S_AXIS_FIFO_58_DMWIDTH/8-1:0] s_axis_fifo_58_tkeep,
    input [S_AXIS_FIFO_58_DMWIDTH/8-1:0] s_axis_fifo_58_tstrb,
    input [S_AXIS_FIFO_58_DMWIDTH-1:0] s_axis_fifo_58_tdata,
    output s_axis_fifo_58_tready,
    output ap_fifo_iarg_58_empty_n,
    output [S_AXIS_FIFO_58_WIDTH-1:0] ap_fifo_iarg_58_dout,
    input ap_fifo_iarg_58_read,
    //input AXI-Stream to FIFO interface 59
    input s_axis_fifo_59_aclk,
    input s_axis_fifo_59_aresetn,
    input s_axis_fifo_59_tlast,
    input s_axis_fifo_59_tvalid,
    input [S_AXIS_FIFO_59_DMWIDTH/8-1:0] s_axis_fifo_59_tkeep,
    input [S_AXIS_FIFO_59_DMWIDTH/8-1:0] s_axis_fifo_59_tstrb,
    input [S_AXIS_FIFO_59_DMWIDTH-1:0] s_axis_fifo_59_tdata,
    output s_axis_fifo_59_tready,
    output ap_fifo_iarg_59_empty_n,
    output [S_AXIS_FIFO_59_WIDTH-1:0] ap_fifo_iarg_59_dout,
    input ap_fifo_iarg_59_read,
    //input AXI-Stream to FIFO interface 60
    input s_axis_fifo_60_aclk,
    input s_axis_fifo_60_aresetn,
    input s_axis_fifo_60_tlast,
    input s_axis_fifo_60_tvalid,
    input [S_AXIS_FIFO_60_DMWIDTH/8-1:0] s_axis_fifo_60_tkeep,
    input [S_AXIS_FIFO_60_DMWIDTH/8-1:0] s_axis_fifo_60_tstrb,
    input [S_AXIS_FIFO_60_DMWIDTH-1:0] s_axis_fifo_60_tdata,
    output s_axis_fifo_60_tready,
    output ap_fifo_iarg_60_empty_n,
    output [S_AXIS_FIFO_60_WIDTH-1:0] ap_fifo_iarg_60_dout,
    input ap_fifo_iarg_60_read,
    //input AXI-Stream to FIFO interface 61
    input s_axis_fifo_61_aclk,
    input s_axis_fifo_61_aresetn,
    input s_axis_fifo_61_tlast,
    input s_axis_fifo_61_tvalid,
    input [S_AXIS_FIFO_61_DMWIDTH/8-1:0] s_axis_fifo_61_tkeep,
    input [S_AXIS_FIFO_61_DMWIDTH/8-1:0] s_axis_fifo_61_tstrb,
    input [S_AXIS_FIFO_61_DMWIDTH-1:0] s_axis_fifo_61_tdata,
    output s_axis_fifo_61_tready,
    output ap_fifo_iarg_61_empty_n,
    output [S_AXIS_FIFO_61_WIDTH-1:0] ap_fifo_iarg_61_dout,
    input ap_fifo_iarg_61_read,
    //input AXI-Stream to FIFO interface 62
    input s_axis_fifo_62_aclk,
    input s_axis_fifo_62_aresetn,
    input s_axis_fifo_62_tlast,
    input s_axis_fifo_62_tvalid,
    input [S_AXIS_FIFO_62_DMWIDTH/8-1:0] s_axis_fifo_62_tkeep,
    input [S_AXIS_FIFO_62_DMWIDTH/8-1:0] s_axis_fifo_62_tstrb,
    input [S_AXIS_FIFO_62_DMWIDTH-1:0] s_axis_fifo_62_tdata,
    output s_axis_fifo_62_tready,
    output ap_fifo_iarg_62_empty_n,
    output [S_AXIS_FIFO_62_WIDTH-1:0] ap_fifo_iarg_62_dout,
    input ap_fifo_iarg_62_read,
    //input AXI-Stream to FIFO interface 63
    input s_axis_fifo_63_aclk,
    input s_axis_fifo_63_aresetn,
    input s_axis_fifo_63_tlast,
    input s_axis_fifo_63_tvalid,
    input [S_AXIS_FIFO_63_DMWIDTH/8-1:0] s_axis_fifo_63_tkeep,
    input [S_AXIS_FIFO_63_DMWIDTH/8-1:0] s_axis_fifo_63_tstrb,
    input [S_AXIS_FIFO_63_DMWIDTH-1:0] s_axis_fifo_63_tdata,
    output s_axis_fifo_63_tready,
    output ap_fifo_iarg_63_empty_n,
    output [S_AXIS_FIFO_63_WIDTH-1:0] ap_fifo_iarg_63_dout,
    input ap_fifo_iarg_63_read,
    //input AXI-Stream to FIFO interface 64
    input s_axis_fifo_64_aclk,
    input s_axis_fifo_64_aresetn,
    input s_axis_fifo_64_tlast,
    input s_axis_fifo_64_tvalid,
    input [S_AXIS_FIFO_64_DMWIDTH/8-1:0] s_axis_fifo_64_tkeep,
    input [S_AXIS_FIFO_64_DMWIDTH/8-1:0] s_axis_fifo_64_tstrb,
    input [S_AXIS_FIFO_64_DMWIDTH-1:0] s_axis_fifo_64_tdata,
    output s_axis_fifo_64_tready,
    output ap_fifo_iarg_64_empty_n,
    output [S_AXIS_FIFO_64_WIDTH-1:0] ap_fifo_iarg_64_dout,
    input ap_fifo_iarg_64_read,
    //input AXI-Stream to FIFO interface 65
    input s_axis_fifo_65_aclk,
    input s_axis_fifo_65_aresetn,
    input s_axis_fifo_65_tlast,
    input s_axis_fifo_65_tvalid,
    input [S_AXIS_FIFO_65_DMWIDTH/8-1:0] s_axis_fifo_65_tkeep,
    input [S_AXIS_FIFO_65_DMWIDTH/8-1:0] s_axis_fifo_65_tstrb,
    input [S_AXIS_FIFO_65_DMWIDTH-1:0] s_axis_fifo_65_tdata,
    output s_axis_fifo_65_tready,
    output ap_fifo_iarg_65_empty_n,
    output [S_AXIS_FIFO_65_WIDTH-1:0] ap_fifo_iarg_65_dout,
    input ap_fifo_iarg_65_read,
    //input AXI-Stream to FIFO interface 66
    input s_axis_fifo_66_aclk,
    input s_axis_fifo_66_aresetn,
    input s_axis_fifo_66_tlast,
    input s_axis_fifo_66_tvalid,
    input [S_AXIS_FIFO_66_DMWIDTH/8-1:0] s_axis_fifo_66_tkeep,
    input [S_AXIS_FIFO_66_DMWIDTH/8-1:0] s_axis_fifo_66_tstrb,
    input [S_AXIS_FIFO_66_DMWIDTH-1:0] s_axis_fifo_66_tdata,
    output s_axis_fifo_66_tready,
    output ap_fifo_iarg_66_empty_n,
    output [S_AXIS_FIFO_66_WIDTH-1:0] ap_fifo_iarg_66_dout,
    input ap_fifo_iarg_66_read,
    //input AXI-Stream to FIFO interface 67
    input s_axis_fifo_67_aclk,
    input s_axis_fifo_67_aresetn,
    input s_axis_fifo_67_tlast,
    input s_axis_fifo_67_tvalid,
    input [S_AXIS_FIFO_67_DMWIDTH/8-1:0] s_axis_fifo_67_tkeep,
    input [S_AXIS_FIFO_67_DMWIDTH/8-1:0] s_axis_fifo_67_tstrb,
    input [S_AXIS_FIFO_67_DMWIDTH-1:0] s_axis_fifo_67_tdata,
    output s_axis_fifo_67_tready,
    output ap_fifo_iarg_67_empty_n,
    output [S_AXIS_FIFO_67_WIDTH-1:0] ap_fifo_iarg_67_dout,
    input ap_fifo_iarg_67_read,
    //input AXI-Stream to FIFO interface 68
    input s_axis_fifo_68_aclk,
    input s_axis_fifo_68_aresetn,
    input s_axis_fifo_68_tlast,
    input s_axis_fifo_68_tvalid,
    input [S_AXIS_FIFO_68_DMWIDTH/8-1:0] s_axis_fifo_68_tkeep,
    input [S_AXIS_FIFO_68_DMWIDTH/8-1:0] s_axis_fifo_68_tstrb,
    input [S_AXIS_FIFO_68_DMWIDTH-1:0] s_axis_fifo_68_tdata,
    output s_axis_fifo_68_tready,
    output ap_fifo_iarg_68_empty_n,
    output [S_AXIS_FIFO_68_WIDTH-1:0] ap_fifo_iarg_68_dout,
    input ap_fifo_iarg_68_read,
    //input AXI-Stream to FIFO interface 69
    input s_axis_fifo_69_aclk,
    input s_axis_fifo_69_aresetn,
    input s_axis_fifo_69_tlast,
    input s_axis_fifo_69_tvalid,
    input [S_AXIS_FIFO_69_DMWIDTH/8-1:0] s_axis_fifo_69_tkeep,
    input [S_AXIS_FIFO_69_DMWIDTH/8-1:0] s_axis_fifo_69_tstrb,
    input [S_AXIS_FIFO_69_DMWIDTH-1:0] s_axis_fifo_69_tdata,
    output s_axis_fifo_69_tready,
    output ap_fifo_iarg_69_empty_n,
    output [S_AXIS_FIFO_69_WIDTH-1:0] ap_fifo_iarg_69_dout,
    input ap_fifo_iarg_69_read,
    //input AXI-Stream to FIFO interface 70
    input s_axis_fifo_70_aclk,
    input s_axis_fifo_70_aresetn,
    input s_axis_fifo_70_tlast,
    input s_axis_fifo_70_tvalid,
    input [S_AXIS_FIFO_70_DMWIDTH/8-1:0] s_axis_fifo_70_tkeep,
    input [S_AXIS_FIFO_70_DMWIDTH/8-1:0] s_axis_fifo_70_tstrb,
    input [S_AXIS_FIFO_70_DMWIDTH-1:0] s_axis_fifo_70_tdata,
    output s_axis_fifo_70_tready,
    output ap_fifo_iarg_70_empty_n,
    output [S_AXIS_FIFO_70_WIDTH-1:0] ap_fifo_iarg_70_dout,
    input ap_fifo_iarg_70_read,
    //input AXI-Stream to FIFO interface 71
    input s_axis_fifo_71_aclk,
    input s_axis_fifo_71_aresetn,
    input s_axis_fifo_71_tlast,
    input s_axis_fifo_71_tvalid,
    input [S_AXIS_FIFO_71_DMWIDTH/8-1:0] s_axis_fifo_71_tkeep,
    input [S_AXIS_FIFO_71_DMWIDTH/8-1:0] s_axis_fifo_71_tstrb,
    input [S_AXIS_FIFO_71_DMWIDTH-1:0] s_axis_fifo_71_tdata,
    output s_axis_fifo_71_tready,
    output ap_fifo_iarg_71_empty_n,
    output [S_AXIS_FIFO_71_WIDTH-1:0] ap_fifo_iarg_71_dout,
    input ap_fifo_iarg_71_read,
    //input AXI-Stream to FIFO interface 72
    input s_axis_fifo_72_aclk,
    input s_axis_fifo_72_aresetn,
    input s_axis_fifo_72_tlast,
    input s_axis_fifo_72_tvalid,
    input [S_AXIS_FIFO_72_DMWIDTH/8-1:0] s_axis_fifo_72_tkeep,
    input [S_AXIS_FIFO_72_DMWIDTH/8-1:0] s_axis_fifo_72_tstrb,
    input [S_AXIS_FIFO_72_DMWIDTH-1:0] s_axis_fifo_72_tdata,
    output s_axis_fifo_72_tready,
    output ap_fifo_iarg_72_empty_n,
    output [S_AXIS_FIFO_72_WIDTH-1:0] ap_fifo_iarg_72_dout,
    input ap_fifo_iarg_72_read,
    //input AXI-Stream to FIFO interface 73
    input s_axis_fifo_73_aclk,
    input s_axis_fifo_73_aresetn,
    input s_axis_fifo_73_tlast,
    input s_axis_fifo_73_tvalid,
    input [S_AXIS_FIFO_73_DMWIDTH/8-1:0] s_axis_fifo_73_tkeep,
    input [S_AXIS_FIFO_73_DMWIDTH/8-1:0] s_axis_fifo_73_tstrb,
    input [S_AXIS_FIFO_73_DMWIDTH-1:0] s_axis_fifo_73_tdata,
    output s_axis_fifo_73_tready,
    output ap_fifo_iarg_73_empty_n,
    output [S_AXIS_FIFO_73_WIDTH-1:0] ap_fifo_iarg_73_dout,
    input ap_fifo_iarg_73_read,
    //input AXI-Stream to FIFO interface 74
    input s_axis_fifo_74_aclk,
    input s_axis_fifo_74_aresetn,
    input s_axis_fifo_74_tlast,
    input s_axis_fifo_74_tvalid,
    input [S_AXIS_FIFO_74_DMWIDTH/8-1:0] s_axis_fifo_74_tkeep,
    input [S_AXIS_FIFO_74_DMWIDTH/8-1:0] s_axis_fifo_74_tstrb,
    input [S_AXIS_FIFO_74_DMWIDTH-1:0] s_axis_fifo_74_tdata,
    output s_axis_fifo_74_tready,
    output ap_fifo_iarg_74_empty_n,
    output [S_AXIS_FIFO_74_WIDTH-1:0] ap_fifo_iarg_74_dout,
    input ap_fifo_iarg_74_read,
    //input AXI-Stream to FIFO interface 75
    input s_axis_fifo_75_aclk,
    input s_axis_fifo_75_aresetn,
    input s_axis_fifo_75_tlast,
    input s_axis_fifo_75_tvalid,
    input [S_AXIS_FIFO_75_DMWIDTH/8-1:0] s_axis_fifo_75_tkeep,
    input [S_AXIS_FIFO_75_DMWIDTH/8-1:0] s_axis_fifo_75_tstrb,
    input [S_AXIS_FIFO_75_DMWIDTH-1:0] s_axis_fifo_75_tdata,
    output s_axis_fifo_75_tready,
    output ap_fifo_iarg_75_empty_n,
    output [S_AXIS_FIFO_75_WIDTH-1:0] ap_fifo_iarg_75_dout,
    input ap_fifo_iarg_75_read,
    //input AXI-Stream to FIFO interface 76
    input s_axis_fifo_76_aclk,
    input s_axis_fifo_76_aresetn,
    input s_axis_fifo_76_tlast,
    input s_axis_fifo_76_tvalid,
    input [S_AXIS_FIFO_76_DMWIDTH/8-1:0] s_axis_fifo_76_tkeep,
    input [S_AXIS_FIFO_76_DMWIDTH/8-1:0] s_axis_fifo_76_tstrb,
    input [S_AXIS_FIFO_76_DMWIDTH-1:0] s_axis_fifo_76_tdata,
    output s_axis_fifo_76_tready,
    output ap_fifo_iarg_76_empty_n,
    output [S_AXIS_FIFO_76_WIDTH-1:0] ap_fifo_iarg_76_dout,
    input ap_fifo_iarg_76_read,
    //input AXI-Stream to FIFO interface 77
    input s_axis_fifo_77_aclk,
    input s_axis_fifo_77_aresetn,
    input s_axis_fifo_77_tlast,
    input s_axis_fifo_77_tvalid,
    input [S_AXIS_FIFO_77_DMWIDTH/8-1:0] s_axis_fifo_77_tkeep,
    input [S_AXIS_FIFO_77_DMWIDTH/8-1:0] s_axis_fifo_77_tstrb,
    input [S_AXIS_FIFO_77_DMWIDTH-1:0] s_axis_fifo_77_tdata,
    output s_axis_fifo_77_tready,
    output ap_fifo_iarg_77_empty_n,
    output [S_AXIS_FIFO_77_WIDTH-1:0] ap_fifo_iarg_77_dout,
    input ap_fifo_iarg_77_read,
    //input AXI-Stream to FIFO interface 78
    input s_axis_fifo_78_aclk,
    input s_axis_fifo_78_aresetn,
    input s_axis_fifo_78_tlast,
    input s_axis_fifo_78_tvalid,
    input [S_AXIS_FIFO_78_DMWIDTH/8-1:0] s_axis_fifo_78_tkeep,
    input [S_AXIS_FIFO_78_DMWIDTH/8-1:0] s_axis_fifo_78_tstrb,
    input [S_AXIS_FIFO_78_DMWIDTH-1:0] s_axis_fifo_78_tdata,
    output s_axis_fifo_78_tready,
    output ap_fifo_iarg_78_empty_n,
    output [S_AXIS_FIFO_78_WIDTH-1:0] ap_fifo_iarg_78_dout,
    input ap_fifo_iarg_78_read,
    //input AXI-Stream to FIFO interface 79
    input s_axis_fifo_79_aclk,
    input s_axis_fifo_79_aresetn,
    input s_axis_fifo_79_tlast,
    input s_axis_fifo_79_tvalid,
    input [S_AXIS_FIFO_79_DMWIDTH/8-1:0] s_axis_fifo_79_tkeep,
    input [S_AXIS_FIFO_79_DMWIDTH/8-1:0] s_axis_fifo_79_tstrb,
    input [S_AXIS_FIFO_79_DMWIDTH-1:0] s_axis_fifo_79_tdata,
    output s_axis_fifo_79_tready,
    output ap_fifo_iarg_79_empty_n,
    output [S_AXIS_FIFO_79_WIDTH-1:0] ap_fifo_iarg_79_dout,
    input ap_fifo_iarg_79_read,
    //input AXI-Stream to FIFO interface 80
    input s_axis_fifo_80_aclk,
    input s_axis_fifo_80_aresetn,
    input s_axis_fifo_80_tlast,
    input s_axis_fifo_80_tvalid,
    input [S_AXIS_FIFO_80_DMWIDTH/8-1:0] s_axis_fifo_80_tkeep,
    input [S_AXIS_FIFO_80_DMWIDTH/8-1:0] s_axis_fifo_80_tstrb,
    input [S_AXIS_FIFO_80_DMWIDTH-1:0] s_axis_fifo_80_tdata,
    output s_axis_fifo_80_tready,
    output ap_fifo_iarg_80_empty_n,
    output [S_AXIS_FIFO_80_WIDTH-1:0] ap_fifo_iarg_80_dout,
    input ap_fifo_iarg_80_read,
    //input AXI-Stream to FIFO interface 81
    input s_axis_fifo_81_aclk,
    input s_axis_fifo_81_aresetn,
    input s_axis_fifo_81_tlast,
    input s_axis_fifo_81_tvalid,
    input [S_AXIS_FIFO_81_DMWIDTH/8-1:0] s_axis_fifo_81_tkeep,
    input [S_AXIS_FIFO_81_DMWIDTH/8-1:0] s_axis_fifo_81_tstrb,
    input [S_AXIS_FIFO_81_DMWIDTH-1:0] s_axis_fifo_81_tdata,
    output s_axis_fifo_81_tready,
    output ap_fifo_iarg_81_empty_n,
    output [S_AXIS_FIFO_81_WIDTH-1:0] ap_fifo_iarg_81_dout,
    input ap_fifo_iarg_81_read,
    //input AXI-Stream to FIFO interface 82
    input s_axis_fifo_82_aclk,
    input s_axis_fifo_82_aresetn,
    input s_axis_fifo_82_tlast,
    input s_axis_fifo_82_tvalid,
    input [S_AXIS_FIFO_82_DMWIDTH/8-1:0] s_axis_fifo_82_tkeep,
    input [S_AXIS_FIFO_82_DMWIDTH/8-1:0] s_axis_fifo_82_tstrb,
    input [S_AXIS_FIFO_82_DMWIDTH-1:0] s_axis_fifo_82_tdata,
    output s_axis_fifo_82_tready,
    output ap_fifo_iarg_82_empty_n,
    output [S_AXIS_FIFO_82_WIDTH-1:0] ap_fifo_iarg_82_dout,
    input ap_fifo_iarg_82_read,
    //input AXI-Stream to FIFO interface 83
    input s_axis_fifo_83_aclk,
    input s_axis_fifo_83_aresetn,
    input s_axis_fifo_83_tlast,
    input s_axis_fifo_83_tvalid,
    input [S_AXIS_FIFO_83_DMWIDTH/8-1:0] s_axis_fifo_83_tkeep,
    input [S_AXIS_FIFO_83_DMWIDTH/8-1:0] s_axis_fifo_83_tstrb,
    input [S_AXIS_FIFO_83_DMWIDTH-1:0] s_axis_fifo_83_tdata,
    output s_axis_fifo_83_tready,
    output ap_fifo_iarg_83_empty_n,
    output [S_AXIS_FIFO_83_WIDTH-1:0] ap_fifo_iarg_83_dout,
    input ap_fifo_iarg_83_read,
    //input AXI-Stream to FIFO interface 84
    input s_axis_fifo_84_aclk,
    input s_axis_fifo_84_aresetn,
    input s_axis_fifo_84_tlast,
    input s_axis_fifo_84_tvalid,
    input [S_AXIS_FIFO_84_DMWIDTH/8-1:0] s_axis_fifo_84_tkeep,
    input [S_AXIS_FIFO_84_DMWIDTH/8-1:0] s_axis_fifo_84_tstrb,
    input [S_AXIS_FIFO_84_DMWIDTH-1:0] s_axis_fifo_84_tdata,
    output s_axis_fifo_84_tready,
    output ap_fifo_iarg_84_empty_n,
    output [S_AXIS_FIFO_84_WIDTH-1:0] ap_fifo_iarg_84_dout,
    input ap_fifo_iarg_84_read,
    //input AXI-Stream to FIFO interface 85
    input s_axis_fifo_85_aclk,
    input s_axis_fifo_85_aresetn,
    input s_axis_fifo_85_tlast,
    input s_axis_fifo_85_tvalid,
    input [S_AXIS_FIFO_85_DMWIDTH/8-1:0] s_axis_fifo_85_tkeep,
    input [S_AXIS_FIFO_85_DMWIDTH/8-1:0] s_axis_fifo_85_tstrb,
    input [S_AXIS_FIFO_85_DMWIDTH-1:0] s_axis_fifo_85_tdata,
    output s_axis_fifo_85_tready,
    output ap_fifo_iarg_85_empty_n,
    output [S_AXIS_FIFO_85_WIDTH-1:0] ap_fifo_iarg_85_dout,
    input ap_fifo_iarg_85_read,
    //input AXI-Stream to FIFO interface 86
    input s_axis_fifo_86_aclk,
    input s_axis_fifo_86_aresetn,
    input s_axis_fifo_86_tlast,
    input s_axis_fifo_86_tvalid,
    input [S_AXIS_FIFO_86_DMWIDTH/8-1:0] s_axis_fifo_86_tkeep,
    input [S_AXIS_FIFO_86_DMWIDTH/8-1:0] s_axis_fifo_86_tstrb,
    input [S_AXIS_FIFO_86_DMWIDTH-1:0] s_axis_fifo_86_tdata,
    output s_axis_fifo_86_tready,
    output ap_fifo_iarg_86_empty_n,
    output [S_AXIS_FIFO_86_WIDTH-1:0] ap_fifo_iarg_86_dout,
    input ap_fifo_iarg_86_read,
    //input AXI-Stream to FIFO interface 87
    input s_axis_fifo_87_aclk,
    input s_axis_fifo_87_aresetn,
    input s_axis_fifo_87_tlast,
    input s_axis_fifo_87_tvalid,
    input [S_AXIS_FIFO_87_DMWIDTH/8-1:0] s_axis_fifo_87_tkeep,
    input [S_AXIS_FIFO_87_DMWIDTH/8-1:0] s_axis_fifo_87_tstrb,
    input [S_AXIS_FIFO_87_DMWIDTH-1:0] s_axis_fifo_87_tdata,
    output s_axis_fifo_87_tready,
    output ap_fifo_iarg_87_empty_n,
    output [S_AXIS_FIFO_87_WIDTH-1:0] ap_fifo_iarg_87_dout,
    input ap_fifo_iarg_87_read,
    //input AXI-Stream to FIFO interface 88
    input s_axis_fifo_88_aclk,
    input s_axis_fifo_88_aresetn,
    input s_axis_fifo_88_tlast,
    input s_axis_fifo_88_tvalid,
    input [S_AXIS_FIFO_88_DMWIDTH/8-1:0] s_axis_fifo_88_tkeep,
    input [S_AXIS_FIFO_88_DMWIDTH/8-1:0] s_axis_fifo_88_tstrb,
    input [S_AXIS_FIFO_88_DMWIDTH-1:0] s_axis_fifo_88_tdata,
    output s_axis_fifo_88_tready,
    output ap_fifo_iarg_88_empty_n,
    output [S_AXIS_FIFO_88_WIDTH-1:0] ap_fifo_iarg_88_dout,
    input ap_fifo_iarg_88_read,
    //input AXI-Stream to FIFO interface 89
    input s_axis_fifo_89_aclk,
    input s_axis_fifo_89_aresetn,
    input s_axis_fifo_89_tlast,
    input s_axis_fifo_89_tvalid,
    input [S_AXIS_FIFO_89_DMWIDTH/8-1:0] s_axis_fifo_89_tkeep,
    input [S_AXIS_FIFO_89_DMWIDTH/8-1:0] s_axis_fifo_89_tstrb,
    input [S_AXIS_FIFO_89_DMWIDTH-1:0] s_axis_fifo_89_tdata,
    output s_axis_fifo_89_tready,
    output ap_fifo_iarg_89_empty_n,
    output [S_AXIS_FIFO_89_WIDTH-1:0] ap_fifo_iarg_89_dout,
    input ap_fifo_iarg_89_read,
    //input AXI-Stream to FIFO interface 90
    input s_axis_fifo_90_aclk,
    input s_axis_fifo_90_aresetn,
    input s_axis_fifo_90_tlast,
    input s_axis_fifo_90_tvalid,
    input [S_AXIS_FIFO_90_DMWIDTH/8-1:0] s_axis_fifo_90_tkeep,
    input [S_AXIS_FIFO_90_DMWIDTH/8-1:0] s_axis_fifo_90_tstrb,
    input [S_AXIS_FIFO_90_DMWIDTH-1:0] s_axis_fifo_90_tdata,
    output s_axis_fifo_90_tready,
    output ap_fifo_iarg_90_empty_n,
    output [S_AXIS_FIFO_90_WIDTH-1:0] ap_fifo_iarg_90_dout,
    input ap_fifo_iarg_90_read,
    //input AXI-Stream to FIFO interface 91
    input s_axis_fifo_91_aclk,
    input s_axis_fifo_91_aresetn,
    input s_axis_fifo_91_tlast,
    input s_axis_fifo_91_tvalid,
    input [S_AXIS_FIFO_91_DMWIDTH/8-1:0] s_axis_fifo_91_tkeep,
    input [S_AXIS_FIFO_91_DMWIDTH/8-1:0] s_axis_fifo_91_tstrb,
    input [S_AXIS_FIFO_91_DMWIDTH-1:0] s_axis_fifo_91_tdata,
    output s_axis_fifo_91_tready,
    output ap_fifo_iarg_91_empty_n,
    output [S_AXIS_FIFO_91_WIDTH-1:0] ap_fifo_iarg_91_dout,
    input ap_fifo_iarg_91_read,
    //input AXI-Stream to FIFO interface 92
    input s_axis_fifo_92_aclk,
    input s_axis_fifo_92_aresetn,
    input s_axis_fifo_92_tlast,
    input s_axis_fifo_92_tvalid,
    input [S_AXIS_FIFO_92_DMWIDTH/8-1:0] s_axis_fifo_92_tkeep,
    input [S_AXIS_FIFO_92_DMWIDTH/8-1:0] s_axis_fifo_92_tstrb,
    input [S_AXIS_FIFO_92_DMWIDTH-1:0] s_axis_fifo_92_tdata,
    output s_axis_fifo_92_tready,
    output ap_fifo_iarg_92_empty_n,
    output [S_AXIS_FIFO_92_WIDTH-1:0] ap_fifo_iarg_92_dout,
    input ap_fifo_iarg_92_read,
    //input AXI-Stream to FIFO interface 93
    input s_axis_fifo_93_aclk,
    input s_axis_fifo_93_aresetn,
    input s_axis_fifo_93_tlast,
    input s_axis_fifo_93_tvalid,
    input [S_AXIS_FIFO_93_DMWIDTH/8-1:0] s_axis_fifo_93_tkeep,
    input [S_AXIS_FIFO_93_DMWIDTH/8-1:0] s_axis_fifo_93_tstrb,
    input [S_AXIS_FIFO_93_DMWIDTH-1:0] s_axis_fifo_93_tdata,
    output s_axis_fifo_93_tready,
    output ap_fifo_iarg_93_empty_n,
    output [S_AXIS_FIFO_93_WIDTH-1:0] ap_fifo_iarg_93_dout,
    input ap_fifo_iarg_93_read,
    //input AXI-Stream to FIFO interface 94
    input s_axis_fifo_94_aclk,
    input s_axis_fifo_94_aresetn,
    input s_axis_fifo_94_tlast,
    input s_axis_fifo_94_tvalid,
    input [S_AXIS_FIFO_94_DMWIDTH/8-1:0] s_axis_fifo_94_tkeep,
    input [S_AXIS_FIFO_94_DMWIDTH/8-1:0] s_axis_fifo_94_tstrb,
    input [S_AXIS_FIFO_94_DMWIDTH-1:0] s_axis_fifo_94_tdata,
    output s_axis_fifo_94_tready,
    output ap_fifo_iarg_94_empty_n,
    output [S_AXIS_FIFO_94_WIDTH-1:0] ap_fifo_iarg_94_dout,
    input ap_fifo_iarg_94_read,
    //input AXI-Stream to FIFO interface 95
    input s_axis_fifo_95_aclk,
    input s_axis_fifo_95_aresetn,
    input s_axis_fifo_95_tlast,
    input s_axis_fifo_95_tvalid,
    input [S_AXIS_FIFO_95_DMWIDTH/8-1:0] s_axis_fifo_95_tkeep,
    input [S_AXIS_FIFO_95_DMWIDTH/8-1:0] s_axis_fifo_95_tstrb,
    input [S_AXIS_FIFO_95_DMWIDTH-1:0] s_axis_fifo_95_tdata,
    output s_axis_fifo_95_tready,
    output ap_fifo_iarg_95_empty_n,
    output [S_AXIS_FIFO_95_WIDTH-1:0] ap_fifo_iarg_95_dout,
    input ap_fifo_iarg_95_read,
    //input AXI-Stream to FIFO interface 96
    input s_axis_fifo_96_aclk,
    input s_axis_fifo_96_aresetn,
    input s_axis_fifo_96_tlast,
    input s_axis_fifo_96_tvalid,
    input [S_AXIS_FIFO_96_DMWIDTH/8-1:0] s_axis_fifo_96_tkeep,
    input [S_AXIS_FIFO_96_DMWIDTH/8-1:0] s_axis_fifo_96_tstrb,
    input [S_AXIS_FIFO_96_DMWIDTH-1:0] s_axis_fifo_96_tdata,
    output s_axis_fifo_96_tready,
    output ap_fifo_iarg_96_empty_n,
    output [S_AXIS_FIFO_96_WIDTH-1:0] ap_fifo_iarg_96_dout,
    input ap_fifo_iarg_96_read,
    //input AXI-Stream to FIFO interface 97
    input s_axis_fifo_97_aclk,
    input s_axis_fifo_97_aresetn,
    input s_axis_fifo_97_tlast,
    input s_axis_fifo_97_tvalid,
    input [S_AXIS_FIFO_97_DMWIDTH/8-1:0] s_axis_fifo_97_tkeep,
    input [S_AXIS_FIFO_97_DMWIDTH/8-1:0] s_axis_fifo_97_tstrb,
    input [S_AXIS_FIFO_97_DMWIDTH-1:0] s_axis_fifo_97_tdata,
    output s_axis_fifo_97_tready,
    output ap_fifo_iarg_97_empty_n,
    output [S_AXIS_FIFO_97_WIDTH-1:0] ap_fifo_iarg_97_dout,
    input ap_fifo_iarg_97_read,
    //input AXI-Stream to FIFO interface 98
    input s_axis_fifo_98_aclk,
    input s_axis_fifo_98_aresetn,
    input s_axis_fifo_98_tlast,
    input s_axis_fifo_98_tvalid,
    input [S_AXIS_FIFO_98_DMWIDTH/8-1:0] s_axis_fifo_98_tkeep,
    input [S_AXIS_FIFO_98_DMWIDTH/8-1:0] s_axis_fifo_98_tstrb,
    input [S_AXIS_FIFO_98_DMWIDTH-1:0] s_axis_fifo_98_tdata,
    output s_axis_fifo_98_tready,
    output ap_fifo_iarg_98_empty_n,
    output [S_AXIS_FIFO_98_WIDTH-1:0] ap_fifo_iarg_98_dout,
    input ap_fifo_iarg_98_read,
    //input AXI-Stream to FIFO interface 99
    input s_axis_fifo_99_aclk,
    input s_axis_fifo_99_aresetn,
    input s_axis_fifo_99_tlast,
    input s_axis_fifo_99_tvalid,
    input [S_AXIS_FIFO_99_DMWIDTH/8-1:0] s_axis_fifo_99_tkeep,
    input [S_AXIS_FIFO_99_DMWIDTH/8-1:0] s_axis_fifo_99_tstrb,
    input [S_AXIS_FIFO_99_DMWIDTH-1:0] s_axis_fifo_99_tdata,
    output s_axis_fifo_99_tready,
    output ap_fifo_iarg_99_empty_n,
    output [S_AXIS_FIFO_99_WIDTH-1:0] ap_fifo_iarg_99_dout,
    input ap_fifo_iarg_99_read,
    //input AXI-Stream to FIFO interface 100
    input s_axis_fifo_100_aclk,
    input s_axis_fifo_100_aresetn,
    input s_axis_fifo_100_tlast,
    input s_axis_fifo_100_tvalid,
    input [S_AXIS_FIFO_100_DMWIDTH/8-1:0] s_axis_fifo_100_tkeep,
    input [S_AXIS_FIFO_100_DMWIDTH/8-1:0] s_axis_fifo_100_tstrb,
    input [S_AXIS_FIFO_100_DMWIDTH-1:0] s_axis_fifo_100_tdata,
    output s_axis_fifo_100_tready,
    output ap_fifo_iarg_100_empty_n,
    output [S_AXIS_FIFO_100_WIDTH-1:0] ap_fifo_iarg_100_dout,
    input ap_fifo_iarg_100_read,
    //input AXI-Stream to FIFO interface 101
    input s_axis_fifo_101_aclk,
    input s_axis_fifo_101_aresetn,
    input s_axis_fifo_101_tlast,
    input s_axis_fifo_101_tvalid,
    input [S_AXIS_FIFO_101_DMWIDTH/8-1:0] s_axis_fifo_101_tkeep,
    input [S_AXIS_FIFO_101_DMWIDTH/8-1:0] s_axis_fifo_101_tstrb,
    input [S_AXIS_FIFO_101_DMWIDTH-1:0] s_axis_fifo_101_tdata,
    output s_axis_fifo_101_tready,
    output ap_fifo_iarg_101_empty_n,
    output [S_AXIS_FIFO_101_WIDTH-1:0] ap_fifo_iarg_101_dout,
    input ap_fifo_iarg_101_read,
    //input AXI-Stream to FIFO interface 102
    input s_axis_fifo_102_aclk,
    input s_axis_fifo_102_aresetn,
    input s_axis_fifo_102_tlast,
    input s_axis_fifo_102_tvalid,
    input [S_AXIS_FIFO_102_DMWIDTH/8-1:0] s_axis_fifo_102_tkeep,
    input [S_AXIS_FIFO_102_DMWIDTH/8-1:0] s_axis_fifo_102_tstrb,
    input [S_AXIS_FIFO_102_DMWIDTH-1:0] s_axis_fifo_102_tdata,
    output s_axis_fifo_102_tready,
    output ap_fifo_iarg_102_empty_n,
    output [S_AXIS_FIFO_102_WIDTH-1:0] ap_fifo_iarg_102_dout,
    input ap_fifo_iarg_102_read,
    //input AXI-Stream to FIFO interface 103
    input s_axis_fifo_103_aclk,
    input s_axis_fifo_103_aresetn,
    input s_axis_fifo_103_tlast,
    input s_axis_fifo_103_tvalid,
    input [S_AXIS_FIFO_103_DMWIDTH/8-1:0] s_axis_fifo_103_tkeep,
    input [S_AXIS_FIFO_103_DMWIDTH/8-1:0] s_axis_fifo_103_tstrb,
    input [S_AXIS_FIFO_103_DMWIDTH-1:0] s_axis_fifo_103_tdata,
    output s_axis_fifo_103_tready,
    output ap_fifo_iarg_103_empty_n,
    output [S_AXIS_FIFO_103_WIDTH-1:0] ap_fifo_iarg_103_dout,
    input ap_fifo_iarg_103_read,
    //input AXI-Stream to FIFO interface 104
    input s_axis_fifo_104_aclk,
    input s_axis_fifo_104_aresetn,
    input s_axis_fifo_104_tlast,
    input s_axis_fifo_104_tvalid,
    input [S_AXIS_FIFO_104_DMWIDTH/8-1:0] s_axis_fifo_104_tkeep,
    input [S_AXIS_FIFO_104_DMWIDTH/8-1:0] s_axis_fifo_104_tstrb,
    input [S_AXIS_FIFO_104_DMWIDTH-1:0] s_axis_fifo_104_tdata,
    output s_axis_fifo_104_tready,
    output ap_fifo_iarg_104_empty_n,
    output [S_AXIS_FIFO_104_WIDTH-1:0] ap_fifo_iarg_104_dout,
    input ap_fifo_iarg_104_read,
    //input AXI-Stream to FIFO interface 105
    input s_axis_fifo_105_aclk,
    input s_axis_fifo_105_aresetn,
    input s_axis_fifo_105_tlast,
    input s_axis_fifo_105_tvalid,
    input [S_AXIS_FIFO_105_DMWIDTH/8-1:0] s_axis_fifo_105_tkeep,
    input [S_AXIS_FIFO_105_DMWIDTH/8-1:0] s_axis_fifo_105_tstrb,
    input [S_AXIS_FIFO_105_DMWIDTH-1:0] s_axis_fifo_105_tdata,
    output s_axis_fifo_105_tready,
    output ap_fifo_iarg_105_empty_n,
    output [S_AXIS_FIFO_105_WIDTH-1:0] ap_fifo_iarg_105_dout,
    input ap_fifo_iarg_105_read,
    //input AXI-Stream to FIFO interface 106
    input s_axis_fifo_106_aclk,
    input s_axis_fifo_106_aresetn,
    input s_axis_fifo_106_tlast,
    input s_axis_fifo_106_tvalid,
    input [S_AXIS_FIFO_106_DMWIDTH/8-1:0] s_axis_fifo_106_tkeep,
    input [S_AXIS_FIFO_106_DMWIDTH/8-1:0] s_axis_fifo_106_tstrb,
    input [S_AXIS_FIFO_106_DMWIDTH-1:0] s_axis_fifo_106_tdata,
    output s_axis_fifo_106_tready,
    output ap_fifo_iarg_106_empty_n,
    output [S_AXIS_FIFO_106_WIDTH-1:0] ap_fifo_iarg_106_dout,
    input ap_fifo_iarg_106_read,
    //input AXI-Stream to FIFO interface 107
    input s_axis_fifo_107_aclk,
    input s_axis_fifo_107_aresetn,
    input s_axis_fifo_107_tlast,
    input s_axis_fifo_107_tvalid,
    input [S_AXIS_FIFO_107_DMWIDTH/8-1:0] s_axis_fifo_107_tkeep,
    input [S_AXIS_FIFO_107_DMWIDTH/8-1:0] s_axis_fifo_107_tstrb,
    input [S_AXIS_FIFO_107_DMWIDTH-1:0] s_axis_fifo_107_tdata,
    output s_axis_fifo_107_tready,
    output ap_fifo_iarg_107_empty_n,
    output [S_AXIS_FIFO_107_WIDTH-1:0] ap_fifo_iarg_107_dout,
    input ap_fifo_iarg_107_read,
    //input AXI-Stream to FIFO interface 108
    input s_axis_fifo_108_aclk,
    input s_axis_fifo_108_aresetn,
    input s_axis_fifo_108_tlast,
    input s_axis_fifo_108_tvalid,
    input [S_AXIS_FIFO_108_DMWIDTH/8-1:0] s_axis_fifo_108_tkeep,
    input [S_AXIS_FIFO_108_DMWIDTH/8-1:0] s_axis_fifo_108_tstrb,
    input [S_AXIS_FIFO_108_DMWIDTH-1:0] s_axis_fifo_108_tdata,
    output s_axis_fifo_108_tready,
    output ap_fifo_iarg_108_empty_n,
    output [S_AXIS_FIFO_108_WIDTH-1:0] ap_fifo_iarg_108_dout,
    input ap_fifo_iarg_108_read,
    //input AXI-Stream to FIFO interface 109
    input s_axis_fifo_109_aclk,
    input s_axis_fifo_109_aresetn,
    input s_axis_fifo_109_tlast,
    input s_axis_fifo_109_tvalid,
    input [S_AXIS_FIFO_109_DMWIDTH/8-1:0] s_axis_fifo_109_tkeep,
    input [S_AXIS_FIFO_109_DMWIDTH/8-1:0] s_axis_fifo_109_tstrb,
    input [S_AXIS_FIFO_109_DMWIDTH-1:0] s_axis_fifo_109_tdata,
    output s_axis_fifo_109_tready,
    output ap_fifo_iarg_109_empty_n,
    output [S_AXIS_FIFO_109_WIDTH-1:0] ap_fifo_iarg_109_dout,
    input ap_fifo_iarg_109_read,
    //input AXI-Stream to FIFO interface 110
    input s_axis_fifo_110_aclk,
    input s_axis_fifo_110_aresetn,
    input s_axis_fifo_110_tlast,
    input s_axis_fifo_110_tvalid,
    input [S_AXIS_FIFO_110_DMWIDTH/8-1:0] s_axis_fifo_110_tkeep,
    input [S_AXIS_FIFO_110_DMWIDTH/8-1:0] s_axis_fifo_110_tstrb,
    input [S_AXIS_FIFO_110_DMWIDTH-1:0] s_axis_fifo_110_tdata,
    output s_axis_fifo_110_tready,
    output ap_fifo_iarg_110_empty_n,
    output [S_AXIS_FIFO_110_WIDTH-1:0] ap_fifo_iarg_110_dout,
    input ap_fifo_iarg_110_read,
    //input AXI-Stream to FIFO interface 111
    input s_axis_fifo_111_aclk,
    input s_axis_fifo_111_aresetn,
    input s_axis_fifo_111_tlast,
    input s_axis_fifo_111_tvalid,
    input [S_AXIS_FIFO_111_DMWIDTH/8-1:0] s_axis_fifo_111_tkeep,
    input [S_AXIS_FIFO_111_DMWIDTH/8-1:0] s_axis_fifo_111_tstrb,
    input [S_AXIS_FIFO_111_DMWIDTH-1:0] s_axis_fifo_111_tdata,
    output s_axis_fifo_111_tready,
    output ap_fifo_iarg_111_empty_n,
    output [S_AXIS_FIFO_111_WIDTH-1:0] ap_fifo_iarg_111_dout,
    input ap_fifo_iarg_111_read,
    //input AXI-Stream to FIFO interface 112
    input s_axis_fifo_112_aclk,
    input s_axis_fifo_112_aresetn,
    input s_axis_fifo_112_tlast,
    input s_axis_fifo_112_tvalid,
    input [S_AXIS_FIFO_112_DMWIDTH/8-1:0] s_axis_fifo_112_tkeep,
    input [S_AXIS_FIFO_112_DMWIDTH/8-1:0] s_axis_fifo_112_tstrb,
    input [S_AXIS_FIFO_112_DMWIDTH-1:0] s_axis_fifo_112_tdata,
    output s_axis_fifo_112_tready,
    output ap_fifo_iarg_112_empty_n,
    output [S_AXIS_FIFO_112_WIDTH-1:0] ap_fifo_iarg_112_dout,
    input ap_fifo_iarg_112_read,
    //input AXI-Stream to FIFO interface 113
    input s_axis_fifo_113_aclk,
    input s_axis_fifo_113_aresetn,
    input s_axis_fifo_113_tlast,
    input s_axis_fifo_113_tvalid,
    input [S_AXIS_FIFO_113_DMWIDTH/8-1:0] s_axis_fifo_113_tkeep,
    input [S_AXIS_FIFO_113_DMWIDTH/8-1:0] s_axis_fifo_113_tstrb,
    input [S_AXIS_FIFO_113_DMWIDTH-1:0] s_axis_fifo_113_tdata,
    output s_axis_fifo_113_tready,
    output ap_fifo_iarg_113_empty_n,
    output [S_AXIS_FIFO_113_WIDTH-1:0] ap_fifo_iarg_113_dout,
    input ap_fifo_iarg_113_read,
    //input AXI-Stream to FIFO interface 114
    input s_axis_fifo_114_aclk,
    input s_axis_fifo_114_aresetn,
    input s_axis_fifo_114_tlast,
    input s_axis_fifo_114_tvalid,
    input [S_AXIS_FIFO_114_DMWIDTH/8-1:0] s_axis_fifo_114_tkeep,
    input [S_AXIS_FIFO_114_DMWIDTH/8-1:0] s_axis_fifo_114_tstrb,
    input [S_AXIS_FIFO_114_DMWIDTH-1:0] s_axis_fifo_114_tdata,
    output s_axis_fifo_114_tready,
    output ap_fifo_iarg_114_empty_n,
    output [S_AXIS_FIFO_114_WIDTH-1:0] ap_fifo_iarg_114_dout,
    input ap_fifo_iarg_114_read,
    //input AXI-Stream to FIFO interface 115
    input s_axis_fifo_115_aclk,
    input s_axis_fifo_115_aresetn,
    input s_axis_fifo_115_tlast,
    input s_axis_fifo_115_tvalid,
    input [S_AXIS_FIFO_115_DMWIDTH/8-1:0] s_axis_fifo_115_tkeep,
    input [S_AXIS_FIFO_115_DMWIDTH/8-1:0] s_axis_fifo_115_tstrb,
    input [S_AXIS_FIFO_115_DMWIDTH-1:0] s_axis_fifo_115_tdata,
    output s_axis_fifo_115_tready,
    output ap_fifo_iarg_115_empty_n,
    output [S_AXIS_FIFO_115_WIDTH-1:0] ap_fifo_iarg_115_dout,
    input ap_fifo_iarg_115_read,
    //input AXI-Stream to FIFO interface 116
    input s_axis_fifo_116_aclk,
    input s_axis_fifo_116_aresetn,
    input s_axis_fifo_116_tlast,
    input s_axis_fifo_116_tvalid,
    input [S_AXIS_FIFO_116_DMWIDTH/8-1:0] s_axis_fifo_116_tkeep,
    input [S_AXIS_FIFO_116_DMWIDTH/8-1:0] s_axis_fifo_116_tstrb,
    input [S_AXIS_FIFO_116_DMWIDTH-1:0] s_axis_fifo_116_tdata,
    output s_axis_fifo_116_tready,
    output ap_fifo_iarg_116_empty_n,
    output [S_AXIS_FIFO_116_WIDTH-1:0] ap_fifo_iarg_116_dout,
    input ap_fifo_iarg_116_read,
    //input AXI-Stream to FIFO interface 117
    input s_axis_fifo_117_aclk,
    input s_axis_fifo_117_aresetn,
    input s_axis_fifo_117_tlast,
    input s_axis_fifo_117_tvalid,
    input [S_AXIS_FIFO_117_DMWIDTH/8-1:0] s_axis_fifo_117_tkeep,
    input [S_AXIS_FIFO_117_DMWIDTH/8-1:0] s_axis_fifo_117_tstrb,
    input [S_AXIS_FIFO_117_DMWIDTH-1:0] s_axis_fifo_117_tdata,
    output s_axis_fifo_117_tready,
    output ap_fifo_iarg_117_empty_n,
    output [S_AXIS_FIFO_117_WIDTH-1:0] ap_fifo_iarg_117_dout,
    input ap_fifo_iarg_117_read,
    //input AXI-Stream to FIFO interface 118
    input s_axis_fifo_118_aclk,
    input s_axis_fifo_118_aresetn,
    input s_axis_fifo_118_tlast,
    input s_axis_fifo_118_tvalid,
    input [S_AXIS_FIFO_118_DMWIDTH/8-1:0] s_axis_fifo_118_tkeep,
    input [S_AXIS_FIFO_118_DMWIDTH/8-1:0] s_axis_fifo_118_tstrb,
    input [S_AXIS_FIFO_118_DMWIDTH-1:0] s_axis_fifo_118_tdata,
    output s_axis_fifo_118_tready,
    output ap_fifo_iarg_118_empty_n,
    output [S_AXIS_FIFO_118_WIDTH-1:0] ap_fifo_iarg_118_dout,
    input ap_fifo_iarg_118_read,
    //input AXI-Stream to FIFO interface 119
    input s_axis_fifo_119_aclk,
    input s_axis_fifo_119_aresetn,
    input s_axis_fifo_119_tlast,
    input s_axis_fifo_119_tvalid,
    input [S_AXIS_FIFO_119_DMWIDTH/8-1:0] s_axis_fifo_119_tkeep,
    input [S_AXIS_FIFO_119_DMWIDTH/8-1:0] s_axis_fifo_119_tstrb,
    input [S_AXIS_FIFO_119_DMWIDTH-1:0] s_axis_fifo_119_tdata,
    output s_axis_fifo_119_tready,
    output ap_fifo_iarg_119_empty_n,
    output [S_AXIS_FIFO_119_WIDTH-1:0] ap_fifo_iarg_119_dout,
    input ap_fifo_iarg_119_read,
    //input AXI-Stream to FIFO interface 120
    input s_axis_fifo_120_aclk,
    input s_axis_fifo_120_aresetn,
    input s_axis_fifo_120_tlast,
    input s_axis_fifo_120_tvalid,
    input [S_AXIS_FIFO_120_DMWIDTH/8-1:0] s_axis_fifo_120_tkeep,
    input [S_AXIS_FIFO_120_DMWIDTH/8-1:0] s_axis_fifo_120_tstrb,
    input [S_AXIS_FIFO_120_DMWIDTH-1:0] s_axis_fifo_120_tdata,
    output s_axis_fifo_120_tready,
    output ap_fifo_iarg_120_empty_n,
    output [S_AXIS_FIFO_120_WIDTH-1:0] ap_fifo_iarg_120_dout,
    input ap_fifo_iarg_120_read,
    //input AXI-Stream to FIFO interface 121
    input s_axis_fifo_121_aclk,
    input s_axis_fifo_121_aresetn,
    input s_axis_fifo_121_tlast,
    input s_axis_fifo_121_tvalid,
    input [S_AXIS_FIFO_121_DMWIDTH/8-1:0] s_axis_fifo_121_tkeep,
    input [S_AXIS_FIFO_121_DMWIDTH/8-1:0] s_axis_fifo_121_tstrb,
    input [S_AXIS_FIFO_121_DMWIDTH-1:0] s_axis_fifo_121_tdata,
    output s_axis_fifo_121_tready,
    output ap_fifo_iarg_121_empty_n,
    output [S_AXIS_FIFO_121_WIDTH-1:0] ap_fifo_iarg_121_dout,
    input ap_fifo_iarg_121_read,
    //input AXI-Stream to FIFO interface 122
    input s_axis_fifo_122_aclk,
    input s_axis_fifo_122_aresetn,
    input s_axis_fifo_122_tlast,
    input s_axis_fifo_122_tvalid,
    input [S_AXIS_FIFO_122_DMWIDTH/8-1:0] s_axis_fifo_122_tkeep,
    input [S_AXIS_FIFO_122_DMWIDTH/8-1:0] s_axis_fifo_122_tstrb,
    input [S_AXIS_FIFO_122_DMWIDTH-1:0] s_axis_fifo_122_tdata,
    output s_axis_fifo_122_tready,
    output ap_fifo_iarg_122_empty_n,
    output [S_AXIS_FIFO_122_WIDTH-1:0] ap_fifo_iarg_122_dout,
    input ap_fifo_iarg_122_read,
    //input AXI-Stream to FIFO interface 123
    input s_axis_fifo_123_aclk,
    input s_axis_fifo_123_aresetn,
    input s_axis_fifo_123_tlast,
    input s_axis_fifo_123_tvalid,
    input [S_AXIS_FIFO_123_DMWIDTH/8-1:0] s_axis_fifo_123_tkeep,
    input [S_AXIS_FIFO_123_DMWIDTH/8-1:0] s_axis_fifo_123_tstrb,
    input [S_AXIS_FIFO_123_DMWIDTH-1:0] s_axis_fifo_123_tdata,
    output s_axis_fifo_123_tready,
    output ap_fifo_iarg_123_empty_n,
    output [S_AXIS_FIFO_123_WIDTH-1:0] ap_fifo_iarg_123_dout,
    input ap_fifo_iarg_123_read,
    //input AXI-Stream to FIFO interface 124
    input s_axis_fifo_124_aclk,
    input s_axis_fifo_124_aresetn,
    input s_axis_fifo_124_tlast,
    input s_axis_fifo_124_tvalid,
    input [S_AXIS_FIFO_124_DMWIDTH/8-1:0] s_axis_fifo_124_tkeep,
    input [S_AXIS_FIFO_124_DMWIDTH/8-1:0] s_axis_fifo_124_tstrb,
    input [S_AXIS_FIFO_124_DMWIDTH-1:0] s_axis_fifo_124_tdata,
    output s_axis_fifo_124_tready,
    output ap_fifo_iarg_124_empty_n,
    output [S_AXIS_FIFO_124_WIDTH-1:0] ap_fifo_iarg_124_dout,
    input ap_fifo_iarg_124_read,
    //input AXI-Stream to FIFO interface 125
    input s_axis_fifo_125_aclk,
    input s_axis_fifo_125_aresetn,
    input s_axis_fifo_125_tlast,
    input s_axis_fifo_125_tvalid,
    input [S_AXIS_FIFO_125_DMWIDTH/8-1:0] s_axis_fifo_125_tkeep,
    input [S_AXIS_FIFO_125_DMWIDTH/8-1:0] s_axis_fifo_125_tstrb,
    input [S_AXIS_FIFO_125_DMWIDTH-1:0] s_axis_fifo_125_tdata,
    output s_axis_fifo_125_tready,
    output ap_fifo_iarg_125_empty_n,
    output [S_AXIS_FIFO_125_WIDTH-1:0] ap_fifo_iarg_125_dout,
    input ap_fifo_iarg_125_read,
    //input AXI-Stream to FIFO interface 126
    input s_axis_fifo_126_aclk,
    input s_axis_fifo_126_aresetn,
    input s_axis_fifo_126_tlast,
    input s_axis_fifo_126_tvalid,
    input [S_AXIS_FIFO_126_DMWIDTH/8-1:0] s_axis_fifo_126_tkeep,
    input [S_AXIS_FIFO_126_DMWIDTH/8-1:0] s_axis_fifo_126_tstrb,
    input [S_AXIS_FIFO_126_DMWIDTH-1:0] s_axis_fifo_126_tdata,
    output s_axis_fifo_126_tready,
    output ap_fifo_iarg_126_empty_n,
    output [S_AXIS_FIFO_126_WIDTH-1:0] ap_fifo_iarg_126_dout,
    input ap_fifo_iarg_126_read,
    //input AXI-Stream to FIFO interface 127
    input s_axis_fifo_127_aclk,
    input s_axis_fifo_127_aresetn,
    input s_axis_fifo_127_tlast,
    input s_axis_fifo_127_tvalid,
    input [S_AXIS_FIFO_127_DMWIDTH/8-1:0] s_axis_fifo_127_tkeep,
    input [S_AXIS_FIFO_127_DMWIDTH/8-1:0] s_axis_fifo_127_tstrb,
    input [S_AXIS_FIFO_127_DMWIDTH-1:0] s_axis_fifo_127_tdata,
    output s_axis_fifo_127_tready,
    output ap_fifo_iarg_127_empty_n,
    output [S_AXIS_FIFO_127_WIDTH-1:0] ap_fifo_iarg_127_dout,
    input ap_fifo_iarg_127_read
    );
    
// function called round8 rounds value upto next power of 8 if needed
function integer round8 (input integer val);
begin
    for(round8=0; round8<val; round8=round8+8)
        round8=round8;
    end
endfunction
    

    localparam C_MAX_INPUT_FIFOs = 128;
    localparam C_MAX_BIT_WIDTH = 1024;
    localparam [(C_MAX_INPUT_FIFOs*32)-1:0] C_INFIFO_BIT_ARRAY = {S_AXIS_FIFO_127_BYTE_WIDTH,S_AXIS_FIFO_126_BYTE_WIDTH,S_AXIS_FIFO_125_BYTE_WIDTH,S_AXIS_FIFO_124_BYTE_WIDTH,S_AXIS_FIFO_123_BYTE_WIDTH,S_AXIS_FIFO_122_BYTE_WIDTH,S_AXIS_FIFO_121_BYTE_WIDTH,S_AXIS_FIFO_120_BYTE_WIDTH,S_AXIS_FIFO_119_BYTE_WIDTH,S_AXIS_FIFO_118_BYTE_WIDTH,S_AXIS_FIFO_117_BYTE_WIDTH,S_AXIS_FIFO_116_BYTE_WIDTH,S_AXIS_FIFO_115_BYTE_WIDTH,S_AXIS_FIFO_114_BYTE_WIDTH,S_AXIS_FIFO_113_BYTE_WIDTH,S_AXIS_FIFO_112_BYTE_WIDTH,S_AXIS_FIFO_111_BYTE_WIDTH,S_AXIS_FIFO_110_BYTE_WIDTH,S_AXIS_FIFO_109_BYTE_WIDTH,S_AXIS_FIFO_108_BYTE_WIDTH,S_AXIS_FIFO_107_BYTE_WIDTH,S_AXIS_FIFO_106_BYTE_WIDTH,S_AXIS_FIFO_105_BYTE_WIDTH,S_AXIS_FIFO_104_BYTE_WIDTH,S_AXIS_FIFO_103_BYTE_WIDTH,S_AXIS_FIFO_102_BYTE_WIDTH,S_AXIS_FIFO_101_BYTE_WIDTH,S_AXIS_FIFO_100_BYTE_WIDTH,S_AXIS_FIFO_99_BYTE_WIDTH,S_AXIS_FIFO_98_BYTE_WIDTH,S_AXIS_FIFO_97_BYTE_WIDTH,S_AXIS_FIFO_96_BYTE_WIDTH,S_AXIS_FIFO_95_BYTE_WIDTH,S_AXIS_FIFO_94_BYTE_WIDTH,S_AXIS_FIFO_93_BYTE_WIDTH,S_AXIS_FIFO_92_BYTE_WIDTH,S_AXIS_FIFO_91_BYTE_WIDTH,S_AXIS_FIFO_90_BYTE_WIDTH,S_AXIS_FIFO_89_BYTE_WIDTH,S_AXIS_FIFO_88_BYTE_WIDTH,S_AXIS_FIFO_87_BYTE_WIDTH,S_AXIS_FIFO_86_BYTE_WIDTH,S_AXIS_FIFO_85_BYTE_WIDTH,S_AXIS_FIFO_84_BYTE_WIDTH,S_AXIS_FIFO_83_BYTE_WIDTH,S_AXIS_FIFO_82_BYTE_WIDTH,S_AXIS_FIFO_81_BYTE_WIDTH,S_AXIS_FIFO_80_BYTE_WIDTH,S_AXIS_FIFO_79_BYTE_WIDTH,S_AXIS_FIFO_78_BYTE_WIDTH,S_AXIS_FIFO_77_BYTE_WIDTH,S_AXIS_FIFO_76_BYTE_WIDTH,S_AXIS_FIFO_75_BYTE_WIDTH,S_AXIS_FIFO_74_BYTE_WIDTH,S_AXIS_FIFO_73_BYTE_WIDTH,S_AXIS_FIFO_72_BYTE_WIDTH,S_AXIS_FIFO_71_BYTE_WIDTH,S_AXIS_FIFO_70_BYTE_WIDTH,S_AXIS_FIFO_69_BYTE_WIDTH,S_AXIS_FIFO_68_BYTE_WIDTH,S_AXIS_FIFO_67_BYTE_WIDTH,S_AXIS_FIFO_66_BYTE_WIDTH,S_AXIS_FIFO_65_BYTE_WIDTH,S_AXIS_FIFO_64_BYTE_WIDTH,S_AXIS_FIFO_63_BYTE_WIDTH,S_AXIS_FIFO_62_BYTE_WIDTH,S_AXIS_FIFO_61_BYTE_WIDTH,S_AXIS_FIFO_60_BYTE_WIDTH,S_AXIS_FIFO_59_BYTE_WIDTH,S_AXIS_FIFO_58_BYTE_WIDTH,S_AXIS_FIFO_57_BYTE_WIDTH,S_AXIS_FIFO_56_BYTE_WIDTH,S_AXIS_FIFO_55_BYTE_WIDTH,S_AXIS_FIFO_54_BYTE_WIDTH,S_AXIS_FIFO_53_BYTE_WIDTH,S_AXIS_FIFO_52_BYTE_WIDTH,S_AXIS_FIFO_51_BYTE_WIDTH,S_AXIS_FIFO_50_BYTE_WIDTH,S_AXIS_FIFO_49_BYTE_WIDTH,S_AXIS_FIFO_48_BYTE_WIDTH,S_AXIS_FIFO_47_BYTE_WIDTH,S_AXIS_FIFO_46_BYTE_WIDTH,S_AXIS_FIFO_45_BYTE_WIDTH,S_AXIS_FIFO_44_BYTE_WIDTH,S_AXIS_FIFO_43_BYTE_WIDTH,S_AXIS_FIFO_42_BYTE_WIDTH,S_AXIS_FIFO_41_BYTE_WIDTH,S_AXIS_FIFO_40_BYTE_WIDTH,S_AXIS_FIFO_39_BYTE_WIDTH,S_AXIS_FIFO_38_BYTE_WIDTH,S_AXIS_FIFO_37_BYTE_WIDTH,S_AXIS_FIFO_36_BYTE_WIDTH,S_AXIS_FIFO_35_BYTE_WIDTH,S_AXIS_FIFO_34_BYTE_WIDTH,S_AXIS_FIFO_33_BYTE_WIDTH,S_AXIS_FIFO_32_BYTE_WIDTH,S_AXIS_FIFO_31_BYTE_WIDTH,S_AXIS_FIFO_30_BYTE_WIDTH,S_AXIS_FIFO_29_BYTE_WIDTH,S_AXIS_FIFO_28_BYTE_WIDTH,S_AXIS_FIFO_27_BYTE_WIDTH,S_AXIS_FIFO_26_BYTE_WIDTH,S_AXIS_FIFO_25_BYTE_WIDTH,S_AXIS_FIFO_24_BYTE_WIDTH,S_AXIS_FIFO_23_BYTE_WIDTH,S_AXIS_FIFO_22_BYTE_WIDTH,S_AXIS_FIFO_21_BYTE_WIDTH,S_AXIS_FIFO_20_BYTE_WIDTH,S_AXIS_FIFO_19_BYTE_WIDTH,S_AXIS_FIFO_18_BYTE_WIDTH,S_AXIS_FIFO_17_BYTE_WIDTH,S_AXIS_FIFO_16_BYTE_WIDTH,S_AXIS_FIFO_15_BYTE_WIDTH,S_AXIS_FIFO_14_BYTE_WIDTH,S_AXIS_FIFO_13_BYTE_WIDTH,S_AXIS_FIFO_12_BYTE_WIDTH,S_AXIS_FIFO_11_BYTE_WIDTH,S_AXIS_FIFO_10_BYTE_WIDTH,S_AXIS_FIFO_9_BYTE_WIDTH,S_AXIS_FIFO_8_BYTE_WIDTH,S_AXIS_FIFO_7_BYTE_WIDTH,S_AXIS_FIFO_6_BYTE_WIDTH,S_AXIS_FIFO_5_BYTE_WIDTH,S_AXIS_FIFO_4_BYTE_WIDTH,S_AXIS_FIFO_3_BYTE_WIDTH,S_AXIS_FIFO_2_BYTE_WIDTH,S_AXIS_FIFO_1_BYTE_WIDTH,S_AXIS_FIFO_0_BYTE_WIDTH};
    localparam [(C_MAX_INPUT_FIFOs*32)-1:0] C_INFIFO_REAL_ARRAY = {S_AXIS_FIFO_127_WIDTH,S_AXIS_FIFO_126_WIDTH,S_AXIS_FIFO_125_WIDTH,S_AXIS_FIFO_124_WIDTH,S_AXIS_FIFO_123_WIDTH,S_AXIS_FIFO_122_WIDTH,S_AXIS_FIFO_121_WIDTH,S_AXIS_FIFO_120_WIDTH,S_AXIS_FIFO_119_WIDTH,S_AXIS_FIFO_118_WIDTH,S_AXIS_FIFO_117_WIDTH,S_AXIS_FIFO_116_WIDTH,S_AXIS_FIFO_115_WIDTH,S_AXIS_FIFO_114_WIDTH,S_AXIS_FIFO_113_WIDTH,S_AXIS_FIFO_112_WIDTH,S_AXIS_FIFO_111_WIDTH,S_AXIS_FIFO_110_WIDTH,S_AXIS_FIFO_109_WIDTH,S_AXIS_FIFO_108_WIDTH,S_AXIS_FIFO_107_WIDTH,S_AXIS_FIFO_106_WIDTH,S_AXIS_FIFO_105_WIDTH,S_AXIS_FIFO_104_WIDTH,S_AXIS_FIFO_103_WIDTH,S_AXIS_FIFO_102_WIDTH,S_AXIS_FIFO_101_WIDTH,S_AXIS_FIFO_100_WIDTH,S_AXIS_FIFO_99_WIDTH,S_AXIS_FIFO_98_WIDTH,S_AXIS_FIFO_97_WIDTH,S_AXIS_FIFO_96_WIDTH,S_AXIS_FIFO_95_WIDTH,S_AXIS_FIFO_94_WIDTH,S_AXIS_FIFO_93_WIDTH,S_AXIS_FIFO_92_WIDTH,S_AXIS_FIFO_91_WIDTH,S_AXIS_FIFO_90_WIDTH,S_AXIS_FIFO_89_WIDTH,S_AXIS_FIFO_88_WIDTH,S_AXIS_FIFO_87_WIDTH,S_AXIS_FIFO_86_WIDTH,S_AXIS_FIFO_85_WIDTH,S_AXIS_FIFO_84_WIDTH,S_AXIS_FIFO_83_WIDTH,S_AXIS_FIFO_82_WIDTH,S_AXIS_FIFO_81_WIDTH,S_AXIS_FIFO_80_WIDTH,S_AXIS_FIFO_79_WIDTH,S_AXIS_FIFO_78_WIDTH,S_AXIS_FIFO_77_WIDTH,S_AXIS_FIFO_76_WIDTH,S_AXIS_FIFO_75_WIDTH,S_AXIS_FIFO_74_WIDTH,S_AXIS_FIFO_73_WIDTH,S_AXIS_FIFO_72_WIDTH,S_AXIS_FIFO_71_WIDTH,S_AXIS_FIFO_70_WIDTH,S_AXIS_FIFO_69_WIDTH,S_AXIS_FIFO_68_WIDTH,S_AXIS_FIFO_67_WIDTH,S_AXIS_FIFO_66_WIDTH,S_AXIS_FIFO_65_WIDTH,S_AXIS_FIFO_64_WIDTH,S_AXIS_FIFO_63_WIDTH,S_AXIS_FIFO_62_WIDTH,S_AXIS_FIFO_61_WIDTH,S_AXIS_FIFO_60_WIDTH,S_AXIS_FIFO_59_WIDTH,S_AXIS_FIFO_58_WIDTH,S_AXIS_FIFO_57_WIDTH,S_AXIS_FIFO_56_WIDTH,S_AXIS_FIFO_55_WIDTH,S_AXIS_FIFO_54_WIDTH,S_AXIS_FIFO_53_WIDTH,S_AXIS_FIFO_52_WIDTH,S_AXIS_FIFO_51_WIDTH,S_AXIS_FIFO_50_WIDTH,S_AXIS_FIFO_49_WIDTH,S_AXIS_FIFO_48_WIDTH,S_AXIS_FIFO_47_WIDTH,S_AXIS_FIFO_46_WIDTH,S_AXIS_FIFO_45_WIDTH,S_AXIS_FIFO_44_WIDTH,S_AXIS_FIFO_43_WIDTH,S_AXIS_FIFO_42_WIDTH,S_AXIS_FIFO_41_WIDTH,S_AXIS_FIFO_40_WIDTH,S_AXIS_FIFO_39_WIDTH,S_AXIS_FIFO_38_WIDTH,S_AXIS_FIFO_37_WIDTH,S_AXIS_FIFO_36_WIDTH,S_AXIS_FIFO_35_WIDTH,S_AXIS_FIFO_34_WIDTH,S_AXIS_FIFO_33_WIDTH,S_AXIS_FIFO_32_WIDTH,S_AXIS_FIFO_31_WIDTH,S_AXIS_FIFO_30_WIDTH,S_AXIS_FIFO_29_WIDTH,S_AXIS_FIFO_28_WIDTH,S_AXIS_FIFO_27_WIDTH,S_AXIS_FIFO_26_WIDTH,S_AXIS_FIFO_25_WIDTH,S_AXIS_FIFO_24_WIDTH,S_AXIS_FIFO_23_WIDTH,S_AXIS_FIFO_22_WIDTH,S_AXIS_FIFO_21_WIDTH,S_AXIS_FIFO_20_WIDTH,S_AXIS_FIFO_19_WIDTH,S_AXIS_FIFO_18_WIDTH,S_AXIS_FIFO_17_WIDTH,S_AXIS_FIFO_16_WIDTH,S_AXIS_FIFO_15_WIDTH,S_AXIS_FIFO_14_WIDTH,S_AXIS_FIFO_13_WIDTH,S_AXIS_FIFO_12_WIDTH,S_AXIS_FIFO_11_WIDTH,S_AXIS_FIFO_10_WIDTH,S_AXIS_FIFO_9_WIDTH,S_AXIS_FIFO_8_WIDTH,S_AXIS_FIFO_7_WIDTH,S_AXIS_FIFO_6_WIDTH,S_AXIS_FIFO_5_WIDTH,S_AXIS_FIFO_4_WIDTH,S_AXIS_FIFO_3_WIDTH,S_AXIS_FIFO_2_WIDTH,S_AXIS_FIFO_1_WIDTH,S_AXIS_FIFO_0_WIDTH};
    localparam [(C_MAX_INPUT_FIFOs*32)-1:0] C_DEPTH_BIT_ARRAY = {S_AXIS_FIFO_127_DEPTH,S_AXIS_FIFO_126_DEPTH,S_AXIS_FIFO_125_DEPTH,S_AXIS_FIFO_124_DEPTH,S_AXIS_FIFO_123_DEPTH,S_AXIS_FIFO_122_DEPTH,S_AXIS_FIFO_121_DEPTH,S_AXIS_FIFO_120_DEPTH,S_AXIS_FIFO_119_DEPTH,S_AXIS_FIFO_118_DEPTH,S_AXIS_FIFO_117_DEPTH,S_AXIS_FIFO_116_DEPTH,S_AXIS_FIFO_115_DEPTH,S_AXIS_FIFO_114_DEPTH,S_AXIS_FIFO_113_DEPTH,S_AXIS_FIFO_112_DEPTH,S_AXIS_FIFO_111_DEPTH,S_AXIS_FIFO_110_DEPTH,S_AXIS_FIFO_109_DEPTH,S_AXIS_FIFO_108_DEPTH,S_AXIS_FIFO_107_DEPTH,S_AXIS_FIFO_106_DEPTH,S_AXIS_FIFO_105_DEPTH,S_AXIS_FIFO_104_DEPTH,S_AXIS_FIFO_103_DEPTH,S_AXIS_FIFO_102_DEPTH,S_AXIS_FIFO_101_DEPTH,S_AXIS_FIFO_100_DEPTH,S_AXIS_FIFO_99_DEPTH,S_AXIS_FIFO_98_DEPTH,S_AXIS_FIFO_97_DEPTH,S_AXIS_FIFO_96_DEPTH,S_AXIS_FIFO_95_DEPTH,S_AXIS_FIFO_94_DEPTH,S_AXIS_FIFO_93_DEPTH,S_AXIS_FIFO_92_DEPTH,S_AXIS_FIFO_91_DEPTH,S_AXIS_FIFO_90_DEPTH,S_AXIS_FIFO_89_DEPTH,S_AXIS_FIFO_88_DEPTH,S_AXIS_FIFO_87_DEPTH,S_AXIS_FIFO_86_DEPTH,S_AXIS_FIFO_85_DEPTH,S_AXIS_FIFO_84_DEPTH,S_AXIS_FIFO_83_DEPTH,S_AXIS_FIFO_82_DEPTH,S_AXIS_FIFO_81_DEPTH,S_AXIS_FIFO_80_DEPTH,S_AXIS_FIFO_79_DEPTH,S_AXIS_FIFO_78_DEPTH,S_AXIS_FIFO_77_DEPTH,S_AXIS_FIFO_76_DEPTH,S_AXIS_FIFO_75_DEPTH,S_AXIS_FIFO_74_DEPTH,S_AXIS_FIFO_73_DEPTH,S_AXIS_FIFO_72_DEPTH,S_AXIS_FIFO_71_DEPTH,S_AXIS_FIFO_70_DEPTH,S_AXIS_FIFO_69_DEPTH,S_AXIS_FIFO_68_DEPTH,S_AXIS_FIFO_67_DEPTH,S_AXIS_FIFO_66_DEPTH,S_AXIS_FIFO_65_DEPTH,S_AXIS_FIFO_64_DEPTH,S_AXIS_FIFO_63_DEPTH,S_AXIS_FIFO_62_DEPTH,S_AXIS_FIFO_61_DEPTH,S_AXIS_FIFO_60_DEPTH,S_AXIS_FIFO_59_DEPTH,S_AXIS_FIFO_58_DEPTH,S_AXIS_FIFO_57_DEPTH,S_AXIS_FIFO_56_DEPTH,S_AXIS_FIFO_55_DEPTH,S_AXIS_FIFO_54_DEPTH,S_AXIS_FIFO_53_DEPTH,S_AXIS_FIFO_52_DEPTH,S_AXIS_FIFO_51_DEPTH,S_AXIS_FIFO_50_DEPTH,S_AXIS_FIFO_49_DEPTH,S_AXIS_FIFO_48_DEPTH,S_AXIS_FIFO_47_DEPTH,S_AXIS_FIFO_46_DEPTH,S_AXIS_FIFO_45_DEPTH,S_AXIS_FIFO_44_DEPTH,S_AXIS_FIFO_43_DEPTH,S_AXIS_FIFO_42_DEPTH,S_AXIS_FIFO_41_DEPTH,S_AXIS_FIFO_40_DEPTH,S_AXIS_FIFO_39_DEPTH,S_AXIS_FIFO_38_DEPTH,S_AXIS_FIFO_37_DEPTH,S_AXIS_FIFO_36_DEPTH,S_AXIS_FIFO_35_DEPTH,S_AXIS_FIFO_34_DEPTH,S_AXIS_FIFO_33_DEPTH,S_AXIS_FIFO_32_DEPTH,S_AXIS_FIFO_31_DEPTH,S_AXIS_FIFO_30_DEPTH,S_AXIS_FIFO_29_DEPTH,S_AXIS_FIFO_28_DEPTH,S_AXIS_FIFO_27_DEPTH,S_AXIS_FIFO_26_DEPTH,S_AXIS_FIFO_25_DEPTH,S_AXIS_FIFO_24_DEPTH,S_AXIS_FIFO_23_DEPTH,S_AXIS_FIFO_22_DEPTH,S_AXIS_FIFO_21_DEPTH,S_AXIS_FIFO_20_DEPTH,S_AXIS_FIFO_19_DEPTH,S_AXIS_FIFO_18_DEPTH,S_AXIS_FIFO_17_DEPTH,S_AXIS_FIFO_16_DEPTH,S_AXIS_FIFO_15_DEPTH,S_AXIS_FIFO_14_DEPTH,S_AXIS_FIFO_13_DEPTH,S_AXIS_FIFO_12_DEPTH,S_AXIS_FIFO_11_DEPTH,S_AXIS_FIFO_10_DEPTH,S_AXIS_FIFO_9_DEPTH,S_AXIS_FIFO_8_DEPTH,S_AXIS_FIFO_7_DEPTH,S_AXIS_FIFO_6_DEPTH,S_AXIS_FIFO_5_DEPTH,S_AXIS_FIFO_4_DEPTH,S_AXIS_FIFO_3_DEPTH,S_AXIS_FIFO_2_DEPTH,S_AXIS_FIFO_1_DEPTH,S_AXIS_FIFO_0_DEPTH};
    localparam [(C_MAX_INPUT_FIFOs*32)-1:0] C_DMWIDTH_BIT_ARRAY = {S_AXIS_FIFO_127_DMWIDTH,S_AXIS_FIFO_126_DMWIDTH,S_AXIS_FIFO_125_DMWIDTH,S_AXIS_FIFO_124_DMWIDTH,S_AXIS_FIFO_123_DMWIDTH,S_AXIS_FIFO_122_DMWIDTH,S_AXIS_FIFO_121_DMWIDTH,S_AXIS_FIFO_120_DMWIDTH,S_AXIS_FIFO_119_DMWIDTH,S_AXIS_FIFO_118_DMWIDTH,S_AXIS_FIFO_117_DMWIDTH,S_AXIS_FIFO_116_DMWIDTH,S_AXIS_FIFO_115_DMWIDTH,S_AXIS_FIFO_114_DMWIDTH,S_AXIS_FIFO_113_DMWIDTH,S_AXIS_FIFO_112_DMWIDTH,S_AXIS_FIFO_111_DMWIDTH,S_AXIS_FIFO_110_DMWIDTH,S_AXIS_FIFO_109_DMWIDTH,S_AXIS_FIFO_108_DMWIDTH,S_AXIS_FIFO_107_DMWIDTH,S_AXIS_FIFO_106_DMWIDTH,S_AXIS_FIFO_105_DMWIDTH,S_AXIS_FIFO_104_DMWIDTH,S_AXIS_FIFO_103_DMWIDTH,S_AXIS_FIFO_102_DMWIDTH,S_AXIS_FIFO_101_DMWIDTH,S_AXIS_FIFO_100_DMWIDTH,S_AXIS_FIFO_99_DMWIDTH,S_AXIS_FIFO_98_DMWIDTH,S_AXIS_FIFO_97_DMWIDTH,S_AXIS_FIFO_96_DMWIDTH,S_AXIS_FIFO_95_DMWIDTH,S_AXIS_FIFO_94_DMWIDTH,S_AXIS_FIFO_93_DMWIDTH,S_AXIS_FIFO_92_DMWIDTH,S_AXIS_FIFO_91_DMWIDTH,S_AXIS_FIFO_90_DMWIDTH,S_AXIS_FIFO_89_DMWIDTH,S_AXIS_FIFO_88_DMWIDTH,S_AXIS_FIFO_87_DMWIDTH,S_AXIS_FIFO_86_DMWIDTH,S_AXIS_FIFO_85_DMWIDTH,S_AXIS_FIFO_84_DMWIDTH,S_AXIS_FIFO_83_DMWIDTH,S_AXIS_FIFO_82_DMWIDTH,S_AXIS_FIFO_81_DMWIDTH,S_AXIS_FIFO_80_DMWIDTH,S_AXIS_FIFO_79_DMWIDTH,S_AXIS_FIFO_78_DMWIDTH,S_AXIS_FIFO_77_DMWIDTH,S_AXIS_FIFO_76_DMWIDTH,S_AXIS_FIFO_75_DMWIDTH,S_AXIS_FIFO_74_DMWIDTH,S_AXIS_FIFO_73_DMWIDTH,S_AXIS_FIFO_72_DMWIDTH,S_AXIS_FIFO_71_DMWIDTH,S_AXIS_FIFO_70_DMWIDTH,S_AXIS_FIFO_69_DMWIDTH,S_AXIS_FIFO_68_DMWIDTH,S_AXIS_FIFO_67_DMWIDTH,S_AXIS_FIFO_66_DMWIDTH,S_AXIS_FIFO_65_DMWIDTH,S_AXIS_FIFO_64_DMWIDTH,S_AXIS_FIFO_63_DMWIDTH,S_AXIS_FIFO_62_DMWIDTH,S_AXIS_FIFO_61_DMWIDTH,S_AXIS_FIFO_60_DMWIDTH,S_AXIS_FIFO_59_DMWIDTH,S_AXIS_FIFO_58_DMWIDTH,S_AXIS_FIFO_57_DMWIDTH,S_AXIS_FIFO_56_DMWIDTH,S_AXIS_FIFO_55_DMWIDTH,S_AXIS_FIFO_54_DMWIDTH,S_AXIS_FIFO_53_DMWIDTH,S_AXIS_FIFO_52_DMWIDTH,S_AXIS_FIFO_51_DMWIDTH,S_AXIS_FIFO_50_DMWIDTH,S_AXIS_FIFO_49_DMWIDTH,S_AXIS_FIFO_48_DMWIDTH,S_AXIS_FIFO_47_DMWIDTH,S_AXIS_FIFO_46_DMWIDTH,S_AXIS_FIFO_45_DMWIDTH,S_AXIS_FIFO_44_DMWIDTH,S_AXIS_FIFO_43_DMWIDTH,S_AXIS_FIFO_42_DMWIDTH,S_AXIS_FIFO_41_DMWIDTH,S_AXIS_FIFO_40_DMWIDTH,S_AXIS_FIFO_39_DMWIDTH,S_AXIS_FIFO_38_DMWIDTH,S_AXIS_FIFO_37_DMWIDTH,S_AXIS_FIFO_36_DMWIDTH,S_AXIS_FIFO_35_DMWIDTH,S_AXIS_FIFO_34_DMWIDTH,S_AXIS_FIFO_33_DMWIDTH,S_AXIS_FIFO_32_DMWIDTH,S_AXIS_FIFO_31_DMWIDTH,S_AXIS_FIFO_30_DMWIDTH,S_AXIS_FIFO_29_DMWIDTH,S_AXIS_FIFO_28_DMWIDTH,S_AXIS_FIFO_27_DMWIDTH,S_AXIS_FIFO_26_DMWIDTH,S_AXIS_FIFO_25_DMWIDTH,S_AXIS_FIFO_24_DMWIDTH,S_AXIS_FIFO_23_DMWIDTH,S_AXIS_FIFO_22_DMWIDTH,S_AXIS_FIFO_21_DMWIDTH,S_AXIS_FIFO_20_DMWIDTH,S_AXIS_FIFO_19_DMWIDTH,S_AXIS_FIFO_18_DMWIDTH,S_AXIS_FIFO_17_DMWIDTH,S_AXIS_FIFO_16_DMWIDTH,S_AXIS_FIFO_15_DMWIDTH,S_AXIS_FIFO_14_DMWIDTH,S_AXIS_FIFO_13_DMWIDTH,S_AXIS_FIFO_12_DMWIDTH,S_AXIS_FIFO_11_DMWIDTH,S_AXIS_FIFO_10_DMWIDTH,S_AXIS_FIFO_9_DMWIDTH,S_AXIS_FIFO_8_DMWIDTH,S_AXIS_FIFO_7_DMWIDTH,S_AXIS_FIFO_6_DMWIDTH,S_AXIS_FIFO_5_DMWIDTH,S_AXIS_FIFO_4_DMWIDTH,S_AXIS_FIFO_3_DMWIDTH,S_AXIS_FIFO_2_DMWIDTH,S_AXIS_FIFO_1_DMWIDTH,S_AXIS_FIFO_0_DMWIDTH};
    localparam [(C_MAX_INPUT_FIFOs*32)-1:0] C_IS_ASYNC_BIT_ARRAY = {S_AXIS_FIFO_127_IS_ASYNC,S_AXIS_FIFO_126_IS_ASYNC,S_AXIS_FIFO_125_IS_ASYNC,S_AXIS_FIFO_124_IS_ASYNC,S_AXIS_FIFO_123_IS_ASYNC,S_AXIS_FIFO_122_IS_ASYNC,S_AXIS_FIFO_121_IS_ASYNC,S_AXIS_FIFO_120_IS_ASYNC,S_AXIS_FIFO_119_IS_ASYNC,S_AXIS_FIFO_118_IS_ASYNC,S_AXIS_FIFO_117_IS_ASYNC,S_AXIS_FIFO_116_IS_ASYNC,S_AXIS_FIFO_115_IS_ASYNC,S_AXIS_FIFO_114_IS_ASYNC,S_AXIS_FIFO_113_IS_ASYNC,S_AXIS_FIFO_112_IS_ASYNC,S_AXIS_FIFO_111_IS_ASYNC,S_AXIS_FIFO_110_IS_ASYNC,S_AXIS_FIFO_109_IS_ASYNC,S_AXIS_FIFO_108_IS_ASYNC,S_AXIS_FIFO_107_IS_ASYNC,S_AXIS_FIFO_106_IS_ASYNC,S_AXIS_FIFO_105_IS_ASYNC,S_AXIS_FIFO_104_IS_ASYNC,S_AXIS_FIFO_103_IS_ASYNC,S_AXIS_FIFO_102_IS_ASYNC,S_AXIS_FIFO_101_IS_ASYNC,S_AXIS_FIFO_100_IS_ASYNC,S_AXIS_FIFO_99_IS_ASYNC,S_AXIS_FIFO_98_IS_ASYNC,S_AXIS_FIFO_97_IS_ASYNC,S_AXIS_FIFO_96_IS_ASYNC,S_AXIS_FIFO_95_IS_ASYNC,S_AXIS_FIFO_94_IS_ASYNC,S_AXIS_FIFO_93_IS_ASYNC,S_AXIS_FIFO_92_IS_ASYNC,S_AXIS_FIFO_91_IS_ASYNC,S_AXIS_FIFO_90_IS_ASYNC,S_AXIS_FIFO_89_IS_ASYNC,S_AXIS_FIFO_88_IS_ASYNC,S_AXIS_FIFO_87_IS_ASYNC,S_AXIS_FIFO_86_IS_ASYNC,S_AXIS_FIFO_85_IS_ASYNC,S_AXIS_FIFO_84_IS_ASYNC,S_AXIS_FIFO_83_IS_ASYNC,S_AXIS_FIFO_82_IS_ASYNC,S_AXIS_FIFO_81_IS_ASYNC,S_AXIS_FIFO_80_IS_ASYNC,S_AXIS_FIFO_79_IS_ASYNC,S_AXIS_FIFO_78_IS_ASYNC,S_AXIS_FIFO_77_IS_ASYNC,S_AXIS_FIFO_76_IS_ASYNC,S_AXIS_FIFO_75_IS_ASYNC,S_AXIS_FIFO_74_IS_ASYNC,S_AXIS_FIFO_73_IS_ASYNC,S_AXIS_FIFO_72_IS_ASYNC,S_AXIS_FIFO_71_IS_ASYNC,S_AXIS_FIFO_70_IS_ASYNC,S_AXIS_FIFO_69_IS_ASYNC,S_AXIS_FIFO_68_IS_ASYNC,S_AXIS_FIFO_67_IS_ASYNC,S_AXIS_FIFO_66_IS_ASYNC,S_AXIS_FIFO_65_IS_ASYNC,S_AXIS_FIFO_64_IS_ASYNC,S_AXIS_FIFO_63_IS_ASYNC,S_AXIS_FIFO_62_IS_ASYNC,S_AXIS_FIFO_61_IS_ASYNC,S_AXIS_FIFO_60_IS_ASYNC,S_AXIS_FIFO_59_IS_ASYNC,S_AXIS_FIFO_58_IS_ASYNC,S_AXIS_FIFO_57_IS_ASYNC,S_AXIS_FIFO_56_IS_ASYNC,S_AXIS_FIFO_55_IS_ASYNC,S_AXIS_FIFO_54_IS_ASYNC,S_AXIS_FIFO_53_IS_ASYNC,S_AXIS_FIFO_52_IS_ASYNC,S_AXIS_FIFO_51_IS_ASYNC,S_AXIS_FIFO_50_IS_ASYNC,S_AXIS_FIFO_49_IS_ASYNC,S_AXIS_FIFO_48_IS_ASYNC,S_AXIS_FIFO_47_IS_ASYNC,S_AXIS_FIFO_46_IS_ASYNC,S_AXIS_FIFO_45_IS_ASYNC,S_AXIS_FIFO_44_IS_ASYNC,S_AXIS_FIFO_43_IS_ASYNC,S_AXIS_FIFO_42_IS_ASYNC,S_AXIS_FIFO_41_IS_ASYNC,S_AXIS_FIFO_40_IS_ASYNC,S_AXIS_FIFO_39_IS_ASYNC,S_AXIS_FIFO_38_IS_ASYNC,S_AXIS_FIFO_37_IS_ASYNC,S_AXIS_FIFO_36_IS_ASYNC,S_AXIS_FIFO_35_IS_ASYNC,S_AXIS_FIFO_34_IS_ASYNC,S_AXIS_FIFO_33_IS_ASYNC,S_AXIS_FIFO_32_IS_ASYNC,S_AXIS_FIFO_31_IS_ASYNC,S_AXIS_FIFO_30_IS_ASYNC,S_AXIS_FIFO_29_IS_ASYNC,S_AXIS_FIFO_28_IS_ASYNC,S_AXIS_FIFO_27_IS_ASYNC,S_AXIS_FIFO_26_IS_ASYNC,S_AXIS_FIFO_25_IS_ASYNC,S_AXIS_FIFO_24_IS_ASYNC,S_AXIS_FIFO_23_IS_ASYNC,S_AXIS_FIFO_22_IS_ASYNC,S_AXIS_FIFO_21_IS_ASYNC,S_AXIS_FIFO_20_IS_ASYNC,S_AXIS_FIFO_19_IS_ASYNC,S_AXIS_FIFO_18_IS_ASYNC,S_AXIS_FIFO_17_IS_ASYNC,S_AXIS_FIFO_16_IS_ASYNC,S_AXIS_FIFO_15_IS_ASYNC,S_AXIS_FIFO_14_IS_ASYNC,S_AXIS_FIFO_13_IS_ASYNC,S_AXIS_FIFO_12_IS_ASYNC,S_AXIS_FIFO_11_IS_ASYNC,S_AXIS_FIFO_10_IS_ASYNC,S_AXIS_FIFO_9_IS_ASYNC,S_AXIS_FIFO_8_IS_ASYNC,S_AXIS_FIFO_7_IS_ASYNC,S_AXIS_FIFO_6_IS_ASYNC,S_AXIS_FIFO_5_IS_ASYNC,S_AXIS_FIFO_4_IS_ASYNC,S_AXIS_FIFO_3_IS_ASYNC,S_AXIS_FIFO_2_IS_ASYNC,S_AXIS_FIFO_1_IS_ASYNC,S_AXIS_FIFO_0_IS_ASYNC};
    
    wire [C_NUM_INPUT_FIFOs-1:0] axis_clk;
    wire [C_NUM_INPUT_FIFOs-1:0] axis_rst;
    
    wire [C_NUM_INPUT_FIFOs-1:0] tlast;
    wire [C_NUM_INPUT_FIFOs-1:0] tvalid;
    wire [C_MAX_BIT_WIDTH/8-1:0] tkeep [C_NUM_INPUT_FIFOs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] tstrb [C_NUM_INPUT_FIFOs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0]   tdata [C_NUM_INPUT_FIFOs-1:0];
    wire [C_NUM_INPUT_FIFOs-1:0] tready;
    
    wire [C_NUM_INPUT_FIFOs-1:0] dwconv_tlast;
    wire [C_NUM_INPUT_FIFOs-1:0] dwconv_tvalid;
    wire [C_MAX_BIT_WIDTH-1:0] dwconv_tdata [C_NUM_INPUT_FIFOs-1:0];
    wire [C_NUM_INPUT_FIFOs-1:0] dwconv_tready;
    
    wire [C_NUM_INPUT_FIFOs-1:0] trunc_tlast;
    wire [C_NUM_INPUT_FIFOs-1:0] trunc_tvalid;
    wire [C_MAX_BIT_WIDTH-1:0] trunc_tdata [C_NUM_INPUT_FIFOs-1:0];
    wire [C_NUM_INPUT_FIFOs-1:0] trunc_tready;
    
    wire [C_NUM_INPUT_FIFOs-1:0] buf_tlast;
    wire [C_NUM_INPUT_FIFOs-1:0] buf_tvalid;
    wire [C_MAX_BIT_WIDTH-1:0] buf_tdata [C_NUM_INPUT_FIFOs-1:0];
    wire [C_NUM_INPUT_FIFOs-1:0] buf_tready;
    
    wire [C_NUM_INPUT_FIFOs-1:0] read;
    wire [C_NUM_INPUT_FIFOs-1:0] empty;
    wire [C_MAX_BIT_WIDTH-1:0] dout [C_NUM_INPUT_FIFOs-1:0];
    
    //assign inputs to buses, and buses to outputs
    generate
        if(C_NUM_INPUT_FIFOs > 0) begin
            assign axis_clk[0] = s_axis_fifo_0_aclk;
            assign axis_rst[0] = s_axis_fifo_0_aresetn;
            assign tlast[0] = s_axis_fifo_0_tlast;
            assign tvalid[0] = s_axis_fifo_0_tvalid;
            assign read[0] = ap_fifo_iarg_0_read;
            assign tkeep[0][S_AXIS_FIFO_0_DMWIDTH/8-1:0] = s_axis_fifo_0_tkeep;
            assign tstrb[0][S_AXIS_FIFO_0_DMWIDTH/8-1:0] = s_axis_fifo_0_tstrb;
            assign tdata[0][S_AXIS_FIFO_0_DMWIDTH-1:0] = s_axis_fifo_0_tdata;
            assign s_axis_fifo_0_tready = tready[0];
            assign ap_fifo_iarg_0_empty_n = empty[0];
            assign ap_fifo_iarg_0_dout = dout[0][S_AXIS_FIFO_0_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 1) begin
            assign axis_clk[1] = s_axis_fifo_1_aclk;
            assign axis_rst[1] = s_axis_fifo_1_aresetn;
            assign tlast[1] = s_axis_fifo_1_tlast;
            assign tvalid[1] = s_axis_fifo_1_tvalid;
            assign read[1] = ap_fifo_iarg_1_read;
            assign tkeep[1][S_AXIS_FIFO_1_DMWIDTH/8-1:0] = s_axis_fifo_1_tkeep;
            assign tstrb[1][S_AXIS_FIFO_1_DMWIDTH/8-1:0] = s_axis_fifo_1_tstrb;
            assign tdata[1][S_AXIS_FIFO_1_DMWIDTH-1:0] = s_axis_fifo_1_tdata;
            assign s_axis_fifo_1_tready = tready[1];
            assign ap_fifo_iarg_1_empty_n = empty[1];
            assign ap_fifo_iarg_1_dout = dout[1][S_AXIS_FIFO_1_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 2) begin
            assign axis_clk[2] = s_axis_fifo_2_aclk;
            assign axis_rst[2] = s_axis_fifo_2_aresetn;
            assign tlast[2] = s_axis_fifo_2_tlast;
            assign tvalid[2] = s_axis_fifo_2_tvalid;
            assign read[2] = ap_fifo_iarg_2_read;
            assign tkeep[2][S_AXIS_FIFO_2_DMWIDTH/8-1:0] = s_axis_fifo_2_tkeep;
            assign tstrb[2][S_AXIS_FIFO_2_DMWIDTH/8-1:0] = s_axis_fifo_2_tstrb;
            assign tdata[2][S_AXIS_FIFO_2_DMWIDTH-1:0] = s_axis_fifo_2_tdata;
            assign s_axis_fifo_2_tready = tready[2];
            assign ap_fifo_iarg_2_empty_n = empty[2];
            assign ap_fifo_iarg_2_dout = dout[2][S_AXIS_FIFO_2_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 3) begin
            assign axis_clk[3] = s_axis_fifo_3_aclk;
            assign axis_rst[3] = s_axis_fifo_3_aresetn;
            assign tlast[3] = s_axis_fifo_3_tlast;
            assign tvalid[3] = s_axis_fifo_3_tvalid;
            assign read[3] = ap_fifo_iarg_3_read;
            assign tkeep[3][S_AXIS_FIFO_3_DMWIDTH/8-1:0] = s_axis_fifo_3_tkeep;
            assign tstrb[3][S_AXIS_FIFO_3_DMWIDTH/8-1:0] = s_axis_fifo_3_tstrb;
            assign tdata[3][S_AXIS_FIFO_3_DMWIDTH-1:0] = s_axis_fifo_3_tdata;
            assign s_axis_fifo_3_tready = tready[3];
            assign ap_fifo_iarg_3_empty_n = empty[3];
            assign ap_fifo_iarg_3_dout = dout[3][S_AXIS_FIFO_3_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 4) begin
            assign axis_clk[4] = s_axis_fifo_4_aclk;
            assign axis_rst[4] = s_axis_fifo_4_aresetn;
            assign tlast[4] = s_axis_fifo_4_tlast;
            assign tvalid[4] = s_axis_fifo_4_tvalid;
            assign read[4] = ap_fifo_iarg_4_read;
            assign tkeep[4][S_AXIS_FIFO_4_DMWIDTH/8-1:0] = s_axis_fifo_4_tkeep;
            assign tstrb[4][S_AXIS_FIFO_4_DMWIDTH/8-1:0] = s_axis_fifo_4_tstrb;
            assign tdata[4][S_AXIS_FIFO_4_DMWIDTH-1:0] = s_axis_fifo_4_tdata;
            assign s_axis_fifo_4_tready = tready[4];
            assign ap_fifo_iarg_4_empty_n = empty[4];
            assign ap_fifo_iarg_4_dout = dout[4][S_AXIS_FIFO_4_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 5) begin
            assign axis_clk[5] = s_axis_fifo_5_aclk;
            assign axis_rst[5] = s_axis_fifo_5_aresetn;
            assign tlast[5] = s_axis_fifo_5_tlast;
            assign tvalid[5] = s_axis_fifo_5_tvalid;
            assign read[5] = ap_fifo_iarg_5_read;
            assign tkeep[5][S_AXIS_FIFO_5_DMWIDTH/8-1:0] = s_axis_fifo_5_tkeep;
            assign tstrb[5][S_AXIS_FIFO_5_DMWIDTH/8-1:0] = s_axis_fifo_5_tstrb;
            assign tdata[5][S_AXIS_FIFO_5_DMWIDTH-1:0] = s_axis_fifo_5_tdata;
            assign s_axis_fifo_5_tready = tready[5];
            assign ap_fifo_iarg_5_empty_n = empty[5];
            assign ap_fifo_iarg_5_dout = dout[5][S_AXIS_FIFO_5_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 6) begin
            assign axis_clk[6] = s_axis_fifo_6_aclk;
            assign axis_rst[6] = s_axis_fifo_6_aresetn;
            assign tlast[6] = s_axis_fifo_6_tlast;
            assign tvalid[6] = s_axis_fifo_6_tvalid;
            assign read[6] = ap_fifo_iarg_6_read;
            assign tkeep[6][S_AXIS_FIFO_6_DMWIDTH/8-1:0] = s_axis_fifo_6_tkeep;
            assign tstrb[6][S_AXIS_FIFO_6_DMWIDTH/8-1:0] = s_axis_fifo_6_tstrb;
            assign tdata[6][S_AXIS_FIFO_6_DMWIDTH-1:0] = s_axis_fifo_6_tdata;
            assign s_axis_fifo_6_tready = tready[6];
            assign ap_fifo_iarg_6_empty_n = empty[6];
            assign ap_fifo_iarg_6_dout = dout[6][S_AXIS_FIFO_6_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 7) begin
            assign axis_clk[7] = s_axis_fifo_7_aclk;
            assign axis_rst[7] = s_axis_fifo_7_aresetn;
            assign tlast[7] = s_axis_fifo_7_tlast;
            assign tvalid[7] = s_axis_fifo_7_tvalid;
            assign read[7] = ap_fifo_iarg_7_read;
            assign tkeep[7][S_AXIS_FIFO_7_DMWIDTH/8-1:0] = s_axis_fifo_7_tkeep;
            assign tstrb[7][S_AXIS_FIFO_7_DMWIDTH/8-1:0] = s_axis_fifo_7_tstrb;
            assign tdata[7][S_AXIS_FIFO_7_DMWIDTH-1:0] = s_axis_fifo_7_tdata;
            assign s_axis_fifo_7_tready = tready[7];
            assign ap_fifo_iarg_7_empty_n = empty[7];
            assign ap_fifo_iarg_7_dout = dout[7][S_AXIS_FIFO_7_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 8) begin
            assign axis_clk[8] = s_axis_fifo_8_aclk;
            assign axis_rst[8] = s_axis_fifo_8_aresetn;
            assign tlast[8] = s_axis_fifo_8_tlast;
            assign tvalid[8] = s_axis_fifo_8_tvalid;
            assign read[8] = ap_fifo_iarg_8_read;
            assign tkeep[8][S_AXIS_FIFO_8_DMWIDTH/8-1:0] = s_axis_fifo_8_tkeep;
            assign tstrb[8][S_AXIS_FIFO_8_DMWIDTH/8-1:0] = s_axis_fifo_8_tstrb;
            assign tdata[8][S_AXIS_FIFO_8_DMWIDTH-1:0] = s_axis_fifo_8_tdata;
            assign s_axis_fifo_8_tready = tready[8];
            assign ap_fifo_iarg_8_empty_n = empty[8];
            assign ap_fifo_iarg_8_dout = dout[8][S_AXIS_FIFO_8_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 9) begin
            assign axis_clk[9] = s_axis_fifo_9_aclk;
            assign axis_rst[9] = s_axis_fifo_9_aresetn;
            assign tlast[9] = s_axis_fifo_9_tlast;
            assign tvalid[9] = s_axis_fifo_9_tvalid;
            assign read[9] = ap_fifo_iarg_9_read;
            assign tkeep[9][S_AXIS_FIFO_9_DMWIDTH/8-1:0] = s_axis_fifo_9_tkeep;
            assign tstrb[9][S_AXIS_FIFO_9_DMWIDTH/8-1:0] = s_axis_fifo_9_tstrb;
            assign tdata[9][S_AXIS_FIFO_9_DMWIDTH-1:0] = s_axis_fifo_9_tdata;
            assign s_axis_fifo_9_tready = tready[9];
            assign ap_fifo_iarg_9_empty_n = empty[9];
            assign ap_fifo_iarg_9_dout = dout[9][S_AXIS_FIFO_9_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 10) begin
            assign axis_clk[10] = s_axis_fifo_10_aclk;
            assign axis_rst[10] = s_axis_fifo_10_aresetn;
            assign tlast[10] = s_axis_fifo_10_tlast;
            assign tvalid[10] = s_axis_fifo_10_tvalid;
            assign read[10] = ap_fifo_iarg_10_read;
            assign tkeep[10][S_AXIS_FIFO_10_DMWIDTH/8-1:0] = s_axis_fifo_10_tkeep;
            assign tstrb[10][S_AXIS_FIFO_10_DMWIDTH/8-1:0] = s_axis_fifo_10_tstrb;
            assign tdata[10][S_AXIS_FIFO_10_DMWIDTH-1:0] = s_axis_fifo_10_tdata;
            assign s_axis_fifo_10_tready = tready[10];
            assign ap_fifo_iarg_10_empty_n = empty[10];
            assign ap_fifo_iarg_10_dout = dout[10][S_AXIS_FIFO_10_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 11) begin
            assign axis_clk[11] = s_axis_fifo_11_aclk;
            assign axis_rst[11] = s_axis_fifo_11_aresetn;
            assign tlast[11] = s_axis_fifo_11_tlast;
            assign tvalid[11] = s_axis_fifo_11_tvalid;
            assign read[11] = ap_fifo_iarg_11_read;
            assign tkeep[11][S_AXIS_FIFO_11_DMWIDTH/8-1:0] = s_axis_fifo_11_tkeep;
            assign tstrb[11][S_AXIS_FIFO_11_DMWIDTH/8-1:0] = s_axis_fifo_11_tstrb;
            assign tdata[11][S_AXIS_FIFO_11_DMWIDTH-1:0] = s_axis_fifo_11_tdata;
            assign s_axis_fifo_11_tready = tready[11];
            assign ap_fifo_iarg_11_empty_n = empty[11];
            assign ap_fifo_iarg_11_dout = dout[11][S_AXIS_FIFO_11_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 12) begin
            assign axis_clk[12] = s_axis_fifo_12_aclk;
            assign axis_rst[12] = s_axis_fifo_12_aresetn;
            assign tlast[12] = s_axis_fifo_12_tlast;
            assign tvalid[12] = s_axis_fifo_12_tvalid;
            assign read[12] = ap_fifo_iarg_12_read;
            assign tkeep[12][S_AXIS_FIFO_12_DMWIDTH/8-1:0] = s_axis_fifo_12_tkeep;
            assign tstrb[12][S_AXIS_FIFO_12_DMWIDTH/8-1:0] = s_axis_fifo_12_tstrb;
            assign tdata[12][S_AXIS_FIFO_12_DMWIDTH-1:0] = s_axis_fifo_12_tdata;
            assign s_axis_fifo_12_tready = tready[12];
            assign ap_fifo_iarg_12_empty_n = empty[12];
            assign ap_fifo_iarg_12_dout = dout[12][S_AXIS_FIFO_12_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 13) begin
            assign axis_clk[13] = s_axis_fifo_13_aclk;
            assign axis_rst[13] = s_axis_fifo_13_aresetn;
            assign tlast[13] = s_axis_fifo_13_tlast;
            assign tvalid[13] = s_axis_fifo_13_tvalid;
            assign read[13] = ap_fifo_iarg_13_read;
            assign tkeep[13][S_AXIS_FIFO_13_DMWIDTH/8-1:0] = s_axis_fifo_13_tkeep;
            assign tstrb[13][S_AXIS_FIFO_13_DMWIDTH/8-1:0] = s_axis_fifo_13_tstrb;
            assign tdata[13][S_AXIS_FIFO_13_DMWIDTH-1:0] = s_axis_fifo_13_tdata;
            assign s_axis_fifo_13_tready = tready[13];
            assign ap_fifo_iarg_13_empty_n = empty[13];
            assign ap_fifo_iarg_13_dout = dout[13][S_AXIS_FIFO_13_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 14) begin
            assign axis_clk[14] = s_axis_fifo_14_aclk;
            assign axis_rst[14] = s_axis_fifo_14_aresetn;
            assign tlast[14] = s_axis_fifo_14_tlast;
            assign tvalid[14] = s_axis_fifo_14_tvalid;
            assign read[14] = ap_fifo_iarg_14_read;
            assign tkeep[14][S_AXIS_FIFO_14_DMWIDTH/8-1:0] = s_axis_fifo_14_tkeep;
            assign tstrb[14][S_AXIS_FIFO_14_DMWIDTH/8-1:0] = s_axis_fifo_14_tstrb;
            assign tdata[14][S_AXIS_FIFO_14_DMWIDTH-1:0] = s_axis_fifo_14_tdata;
            assign s_axis_fifo_14_tready = tready[14];
            assign ap_fifo_iarg_14_empty_n = empty[14];
            assign ap_fifo_iarg_14_dout = dout[14][S_AXIS_FIFO_14_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 15) begin
            assign axis_clk[15] = s_axis_fifo_15_aclk;
            assign axis_rst[15] = s_axis_fifo_15_aresetn;
            assign tlast[15] = s_axis_fifo_15_tlast;
            assign tvalid[15] = s_axis_fifo_15_tvalid;
            assign read[15] = ap_fifo_iarg_15_read;
            assign tkeep[15][S_AXIS_FIFO_15_DMWIDTH/8-1:0] = s_axis_fifo_15_tkeep;
            assign tstrb[15][S_AXIS_FIFO_15_DMWIDTH/8-1:0] = s_axis_fifo_15_tstrb;
            assign tdata[15][S_AXIS_FIFO_15_DMWIDTH-1:0] = s_axis_fifo_15_tdata;
            assign s_axis_fifo_15_tready = tready[15];
            assign ap_fifo_iarg_15_empty_n = empty[15];
            assign ap_fifo_iarg_15_dout = dout[15][S_AXIS_FIFO_15_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 16) begin
            assign axis_clk[16] = s_axis_fifo_16_aclk;
            assign axis_rst[16] = s_axis_fifo_16_aresetn;
            assign tlast[16] = s_axis_fifo_16_tlast;
            assign tvalid[16] = s_axis_fifo_16_tvalid;
            assign read[16] = ap_fifo_iarg_16_read;
            assign tkeep[16][S_AXIS_FIFO_16_DMWIDTH/8-1:0] = s_axis_fifo_16_tkeep;
            assign tstrb[16][S_AXIS_FIFO_16_DMWIDTH/8-1:0] = s_axis_fifo_16_tstrb;
            assign tdata[16][S_AXIS_FIFO_16_DMWIDTH-1:0] = s_axis_fifo_16_tdata;
            assign s_axis_fifo_16_tready = tready[16];
            assign ap_fifo_iarg_16_empty_n = empty[16];
            assign ap_fifo_iarg_16_dout = dout[16][S_AXIS_FIFO_16_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 17) begin
            assign axis_clk[17] = s_axis_fifo_17_aclk;
            assign axis_rst[17] = s_axis_fifo_17_aresetn;
            assign tlast[17] = s_axis_fifo_17_tlast;
            assign tvalid[17] = s_axis_fifo_17_tvalid;
            assign read[17] = ap_fifo_iarg_17_read;
            assign tkeep[17][S_AXIS_FIFO_17_DMWIDTH/8-1:0] = s_axis_fifo_17_tkeep;
            assign tstrb[17][S_AXIS_FIFO_17_DMWIDTH/8-1:0] = s_axis_fifo_17_tstrb;
            assign tdata[17][S_AXIS_FIFO_17_DMWIDTH-1:0] = s_axis_fifo_17_tdata;
            assign s_axis_fifo_17_tready = tready[17];
            assign ap_fifo_iarg_17_empty_n = empty[17];
            assign ap_fifo_iarg_17_dout = dout[17][S_AXIS_FIFO_17_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 18) begin
            assign axis_clk[18] = s_axis_fifo_18_aclk;
            assign axis_rst[18] = s_axis_fifo_18_aresetn;
            assign tlast[18] = s_axis_fifo_18_tlast;
            assign tvalid[18] = s_axis_fifo_18_tvalid;
            assign read[18] = ap_fifo_iarg_18_read;
            assign tkeep[18][S_AXIS_FIFO_18_DMWIDTH/8-1:0] = s_axis_fifo_18_tkeep;
            assign tstrb[18][S_AXIS_FIFO_18_DMWIDTH/8-1:0] = s_axis_fifo_18_tstrb;
            assign tdata[18][S_AXIS_FIFO_18_DMWIDTH-1:0] = s_axis_fifo_18_tdata;
            assign s_axis_fifo_18_tready = tready[18];
            assign ap_fifo_iarg_18_empty_n = empty[18];
            assign ap_fifo_iarg_18_dout = dout[18][S_AXIS_FIFO_18_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 19) begin
            assign axis_clk[19] = s_axis_fifo_19_aclk;
            assign axis_rst[19] = s_axis_fifo_19_aresetn;
            assign tlast[19] = s_axis_fifo_19_tlast;
            assign tvalid[19] = s_axis_fifo_19_tvalid;
            assign read[19] = ap_fifo_iarg_19_read;
            assign tkeep[19][S_AXIS_FIFO_19_DMWIDTH/8-1:0] = s_axis_fifo_19_tkeep;
            assign tstrb[19][S_AXIS_FIFO_19_DMWIDTH/8-1:0] = s_axis_fifo_19_tstrb;
            assign tdata[19][S_AXIS_FIFO_19_DMWIDTH-1:0] = s_axis_fifo_19_tdata;
            assign s_axis_fifo_19_tready = tready[19];
            assign ap_fifo_iarg_19_empty_n = empty[19];
            assign ap_fifo_iarg_19_dout = dout[19][S_AXIS_FIFO_19_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 20) begin
            assign axis_clk[20] = s_axis_fifo_20_aclk;
            assign axis_rst[20] = s_axis_fifo_20_aresetn;
            assign tlast[20] = s_axis_fifo_20_tlast;
            assign tvalid[20] = s_axis_fifo_20_tvalid;
            assign read[20] = ap_fifo_iarg_20_read;
            assign tkeep[20][S_AXIS_FIFO_20_DMWIDTH/8-1:0] = s_axis_fifo_20_tkeep;
            assign tstrb[20][S_AXIS_FIFO_20_DMWIDTH/8-1:0] = s_axis_fifo_20_tstrb;
            assign tdata[20][S_AXIS_FIFO_20_DMWIDTH-1:0] = s_axis_fifo_20_tdata;
            assign s_axis_fifo_20_tready = tready[20];
            assign ap_fifo_iarg_20_empty_n = empty[20];
            assign ap_fifo_iarg_20_dout = dout[20][S_AXIS_FIFO_20_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 21) begin
            assign axis_clk[21] = s_axis_fifo_21_aclk;
            assign axis_rst[21] = s_axis_fifo_21_aresetn;
            assign tlast[21] = s_axis_fifo_21_tlast;
            assign tvalid[21] = s_axis_fifo_21_tvalid;
            assign read[21] = ap_fifo_iarg_21_read;
            assign tkeep[21][S_AXIS_FIFO_21_DMWIDTH/8-1:0] = s_axis_fifo_21_tkeep;
            assign tstrb[21][S_AXIS_FIFO_21_DMWIDTH/8-1:0] = s_axis_fifo_21_tstrb;
            assign tdata[21][S_AXIS_FIFO_21_DMWIDTH-1:0] = s_axis_fifo_21_tdata;
            assign s_axis_fifo_21_tready = tready[21];
            assign ap_fifo_iarg_21_empty_n = empty[21];
            assign ap_fifo_iarg_21_dout = dout[21][S_AXIS_FIFO_21_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 22) begin
            assign axis_clk[22] = s_axis_fifo_22_aclk;
            assign axis_rst[22] = s_axis_fifo_22_aresetn;
            assign tlast[22] = s_axis_fifo_22_tlast;
            assign tvalid[22] = s_axis_fifo_22_tvalid;
            assign read[22] = ap_fifo_iarg_22_read;
            assign tkeep[22][S_AXIS_FIFO_22_DMWIDTH/8-1:0] = s_axis_fifo_22_tkeep;
            assign tstrb[22][S_AXIS_FIFO_22_DMWIDTH/8-1:0] = s_axis_fifo_22_tstrb;
            assign tdata[22][S_AXIS_FIFO_22_DMWIDTH-1:0] = s_axis_fifo_22_tdata;
            assign s_axis_fifo_22_tready = tready[22];
            assign ap_fifo_iarg_22_empty_n = empty[22];
            assign ap_fifo_iarg_22_dout = dout[22][S_AXIS_FIFO_22_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 23) begin
            assign axis_clk[23] = s_axis_fifo_23_aclk;
            assign axis_rst[23] = s_axis_fifo_23_aresetn;
            assign tlast[23] = s_axis_fifo_23_tlast;
            assign tvalid[23] = s_axis_fifo_23_tvalid;
            assign read[23] = ap_fifo_iarg_23_read;
            assign tkeep[23][S_AXIS_FIFO_23_DMWIDTH/8-1:0] = s_axis_fifo_23_tkeep;
            assign tstrb[23][S_AXIS_FIFO_23_DMWIDTH/8-1:0] = s_axis_fifo_23_tstrb;
            assign tdata[23][S_AXIS_FIFO_23_DMWIDTH-1:0] = s_axis_fifo_23_tdata;
            assign s_axis_fifo_23_tready = tready[23];
            assign ap_fifo_iarg_23_empty_n = empty[23];
            assign ap_fifo_iarg_23_dout = dout[23][S_AXIS_FIFO_23_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 24) begin
            assign axis_clk[24] = s_axis_fifo_24_aclk;
            assign axis_rst[24] = s_axis_fifo_24_aresetn;
            assign tlast[24] = s_axis_fifo_24_tlast;
            assign tvalid[24] = s_axis_fifo_24_tvalid;
            assign read[24] = ap_fifo_iarg_24_read;
            assign tkeep[24][S_AXIS_FIFO_24_DMWIDTH/8-1:0] = s_axis_fifo_24_tkeep;
            assign tstrb[24][S_AXIS_FIFO_24_DMWIDTH/8-1:0] = s_axis_fifo_24_tstrb;
            assign tdata[24][S_AXIS_FIFO_24_DMWIDTH-1:0] = s_axis_fifo_24_tdata;
            assign s_axis_fifo_24_tready = tready[24];
            assign ap_fifo_iarg_24_empty_n = empty[24];
            assign ap_fifo_iarg_24_dout = dout[24][S_AXIS_FIFO_24_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 25) begin
            assign axis_clk[25] = s_axis_fifo_25_aclk;
            assign axis_rst[25] = s_axis_fifo_25_aresetn;
            assign tlast[25] = s_axis_fifo_25_tlast;
            assign tvalid[25] = s_axis_fifo_25_tvalid;
            assign read[25] = ap_fifo_iarg_25_read;
            assign tkeep[25][S_AXIS_FIFO_25_DMWIDTH/8-1:0] = s_axis_fifo_25_tkeep;
            assign tstrb[25][S_AXIS_FIFO_25_DMWIDTH/8-1:0] = s_axis_fifo_25_tstrb;
            assign tdata[25][S_AXIS_FIFO_25_DMWIDTH-1:0] = s_axis_fifo_25_tdata;
            assign s_axis_fifo_25_tready = tready[25];
            assign ap_fifo_iarg_25_empty_n = empty[25];
            assign ap_fifo_iarg_25_dout = dout[25][S_AXIS_FIFO_25_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 26) begin
            assign axis_clk[26] = s_axis_fifo_26_aclk;
            assign axis_rst[26] = s_axis_fifo_26_aresetn;
            assign tlast[26] = s_axis_fifo_26_tlast;
            assign tvalid[26] = s_axis_fifo_26_tvalid;
            assign read[26] = ap_fifo_iarg_26_read;
            assign tkeep[26][S_AXIS_FIFO_26_DMWIDTH/8-1:0] = s_axis_fifo_26_tkeep;
            assign tstrb[26][S_AXIS_FIFO_26_DMWIDTH/8-1:0] = s_axis_fifo_26_tstrb;
            assign tdata[26][S_AXIS_FIFO_26_DMWIDTH-1:0] = s_axis_fifo_26_tdata;
            assign s_axis_fifo_26_tready = tready[26];
            assign ap_fifo_iarg_26_empty_n = empty[26];
            assign ap_fifo_iarg_26_dout = dout[26][S_AXIS_FIFO_26_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 27) begin
            assign axis_clk[27] = s_axis_fifo_27_aclk;
            assign axis_rst[27] = s_axis_fifo_27_aresetn;
            assign tlast[27] = s_axis_fifo_27_tlast;
            assign tvalid[27] = s_axis_fifo_27_tvalid;
            assign read[27] = ap_fifo_iarg_27_read;
            assign tkeep[27][S_AXIS_FIFO_27_DMWIDTH/8-1:0] = s_axis_fifo_27_tkeep;
            assign tstrb[27][S_AXIS_FIFO_27_DMWIDTH/8-1:0] = s_axis_fifo_27_tstrb;
            assign tdata[27][S_AXIS_FIFO_27_DMWIDTH-1:0] = s_axis_fifo_27_tdata;
            assign s_axis_fifo_27_tready = tready[27];
            assign ap_fifo_iarg_27_empty_n = empty[27];
            assign ap_fifo_iarg_27_dout = dout[27][S_AXIS_FIFO_27_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 28) begin
            assign axis_clk[28] = s_axis_fifo_28_aclk;
            assign axis_rst[28] = s_axis_fifo_28_aresetn;
            assign tlast[28] = s_axis_fifo_28_tlast;
            assign tvalid[28] = s_axis_fifo_28_tvalid;
            assign read[28] = ap_fifo_iarg_28_read;
            assign tkeep[28][S_AXIS_FIFO_28_DMWIDTH/8-1:0] = s_axis_fifo_28_tkeep;
            assign tstrb[28][S_AXIS_FIFO_28_DMWIDTH/8-1:0] = s_axis_fifo_28_tstrb;
            assign tdata[28][S_AXIS_FIFO_28_DMWIDTH-1:0] = s_axis_fifo_28_tdata;
            assign s_axis_fifo_28_tready = tready[28];
            assign ap_fifo_iarg_28_empty_n = empty[28];
            assign ap_fifo_iarg_28_dout = dout[28][S_AXIS_FIFO_28_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 29) begin
            assign axis_clk[29] = s_axis_fifo_29_aclk;
            assign axis_rst[29] = s_axis_fifo_29_aresetn;
            assign tlast[29] = s_axis_fifo_29_tlast;
            assign tvalid[29] = s_axis_fifo_29_tvalid;
            assign read[29] = ap_fifo_iarg_29_read;
            assign tkeep[29][S_AXIS_FIFO_29_DMWIDTH/8-1:0] = s_axis_fifo_29_tkeep;
            assign tstrb[29][S_AXIS_FIFO_29_DMWIDTH/8-1:0] = s_axis_fifo_29_tstrb;
            assign tdata[29][S_AXIS_FIFO_29_DMWIDTH-1:0] = s_axis_fifo_29_tdata;
            assign s_axis_fifo_29_tready = tready[29];
            assign ap_fifo_iarg_29_empty_n = empty[29];
            assign ap_fifo_iarg_29_dout = dout[29][S_AXIS_FIFO_29_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 30) begin
            assign axis_clk[30] = s_axis_fifo_30_aclk;
            assign axis_rst[30] = s_axis_fifo_30_aresetn;
            assign tlast[30] = s_axis_fifo_30_tlast;
            assign tvalid[30] = s_axis_fifo_30_tvalid;
            assign read[30] = ap_fifo_iarg_30_read;
            assign tkeep[30][S_AXIS_FIFO_30_DMWIDTH/8-1:0] = s_axis_fifo_30_tkeep;
            assign tstrb[30][S_AXIS_FIFO_30_DMWIDTH/8-1:0] = s_axis_fifo_30_tstrb;
            assign tdata[30][S_AXIS_FIFO_30_DMWIDTH-1:0] = s_axis_fifo_30_tdata;
            assign s_axis_fifo_30_tready = tready[30];
            assign ap_fifo_iarg_30_empty_n = empty[30];
            assign ap_fifo_iarg_30_dout = dout[30][S_AXIS_FIFO_30_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 31) begin
            assign axis_clk[31] = s_axis_fifo_31_aclk;
            assign axis_rst[31] = s_axis_fifo_31_aresetn;
            assign tlast[31] = s_axis_fifo_31_tlast;
            assign tvalid[31] = s_axis_fifo_31_tvalid;
            assign read[31] = ap_fifo_iarg_31_read;
            assign tkeep[31][S_AXIS_FIFO_31_DMWIDTH/8-1:0] = s_axis_fifo_31_tkeep;
            assign tstrb[31][S_AXIS_FIFO_31_DMWIDTH/8-1:0] = s_axis_fifo_31_tstrb;
            assign tdata[31][S_AXIS_FIFO_31_DMWIDTH-1:0] = s_axis_fifo_31_tdata;
            assign s_axis_fifo_31_tready = tready[31];
            assign ap_fifo_iarg_31_empty_n = empty[31];
            assign ap_fifo_iarg_31_dout = dout[31][S_AXIS_FIFO_31_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 32) begin
            assign axis_clk[32] = s_axis_fifo_32_aclk;
            assign axis_rst[32] = s_axis_fifo_32_aresetn;
            assign tlast[32] = s_axis_fifo_32_tlast;
            assign tvalid[32] = s_axis_fifo_32_tvalid;
            assign read[32] = ap_fifo_iarg_32_read;
            assign tkeep[32][S_AXIS_FIFO_32_DMWIDTH/8-1:0] = s_axis_fifo_32_tkeep;
            assign tstrb[32][S_AXIS_FIFO_32_DMWIDTH/8-1:0] = s_axis_fifo_32_tstrb;
            assign tdata[32][S_AXIS_FIFO_32_DMWIDTH-1:0] = s_axis_fifo_32_tdata;
            assign s_axis_fifo_32_tready = tready[32];
            assign ap_fifo_iarg_32_empty_n = empty[32];
            assign ap_fifo_iarg_32_dout = dout[32][S_AXIS_FIFO_32_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 33) begin
            assign axis_clk[33] = s_axis_fifo_33_aclk;
            assign axis_rst[33] = s_axis_fifo_33_aresetn;
            assign tlast[33] = s_axis_fifo_33_tlast;
            assign tvalid[33] = s_axis_fifo_33_tvalid;
            assign read[33] = ap_fifo_iarg_33_read;
            assign tkeep[33][S_AXIS_FIFO_33_DMWIDTH/8-1:0] = s_axis_fifo_33_tkeep;
            assign tstrb[33][S_AXIS_FIFO_33_DMWIDTH/8-1:0] = s_axis_fifo_33_tstrb;
            assign tdata[33][S_AXIS_FIFO_33_DMWIDTH-1:0] = s_axis_fifo_33_tdata;
            assign s_axis_fifo_33_tready = tready[33];
            assign ap_fifo_iarg_33_empty_n = empty[33];
            assign ap_fifo_iarg_33_dout = dout[33][S_AXIS_FIFO_33_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 34) begin
            assign axis_clk[34] = s_axis_fifo_34_aclk;
            assign axis_rst[34] = s_axis_fifo_34_aresetn;
            assign tlast[34] = s_axis_fifo_34_tlast;
            assign tvalid[34] = s_axis_fifo_34_tvalid;
            assign read[34] = ap_fifo_iarg_34_read;
            assign tkeep[34][S_AXIS_FIFO_34_DMWIDTH/8-1:0] = s_axis_fifo_34_tkeep;
            assign tstrb[34][S_AXIS_FIFO_34_DMWIDTH/8-1:0] = s_axis_fifo_34_tstrb;
            assign tdata[34][S_AXIS_FIFO_34_DMWIDTH-1:0] = s_axis_fifo_34_tdata;
            assign s_axis_fifo_34_tready = tready[34];
            assign ap_fifo_iarg_34_empty_n = empty[34];
            assign ap_fifo_iarg_34_dout = dout[34][S_AXIS_FIFO_34_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 35) begin
            assign axis_clk[35] = s_axis_fifo_35_aclk;
            assign axis_rst[35] = s_axis_fifo_35_aresetn;
            assign tlast[35] = s_axis_fifo_35_tlast;
            assign tvalid[35] = s_axis_fifo_35_tvalid;
            assign read[35] = ap_fifo_iarg_35_read;
            assign tkeep[35][S_AXIS_FIFO_35_DMWIDTH/8-1:0] = s_axis_fifo_35_tkeep;
            assign tstrb[35][S_AXIS_FIFO_35_DMWIDTH/8-1:0] = s_axis_fifo_35_tstrb;
            assign tdata[35][S_AXIS_FIFO_35_DMWIDTH-1:0] = s_axis_fifo_35_tdata;
            assign s_axis_fifo_35_tready = tready[35];
            assign ap_fifo_iarg_35_empty_n = empty[35];
            assign ap_fifo_iarg_35_dout = dout[35][S_AXIS_FIFO_35_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 36) begin
            assign axis_clk[36] = s_axis_fifo_36_aclk;
            assign axis_rst[36] = s_axis_fifo_36_aresetn;
            assign tlast[36] = s_axis_fifo_36_tlast;
            assign tvalid[36] = s_axis_fifo_36_tvalid;
            assign read[36] = ap_fifo_iarg_36_read;
            assign tkeep[36][S_AXIS_FIFO_36_DMWIDTH/8-1:0] = s_axis_fifo_36_tkeep;
            assign tstrb[36][S_AXIS_FIFO_36_DMWIDTH/8-1:0] = s_axis_fifo_36_tstrb;
            assign tdata[36][S_AXIS_FIFO_36_DMWIDTH-1:0] = s_axis_fifo_36_tdata;
            assign s_axis_fifo_36_tready = tready[36];
            assign ap_fifo_iarg_36_empty_n = empty[36];
            assign ap_fifo_iarg_36_dout = dout[36][S_AXIS_FIFO_36_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 37) begin
            assign axis_clk[37] = s_axis_fifo_37_aclk;
            assign axis_rst[37] = s_axis_fifo_37_aresetn;
            assign tlast[37] = s_axis_fifo_37_tlast;
            assign tvalid[37] = s_axis_fifo_37_tvalid;
            assign read[37] = ap_fifo_iarg_37_read;
            assign tkeep[37][S_AXIS_FIFO_37_DMWIDTH/8-1:0] = s_axis_fifo_37_tkeep;
            assign tstrb[37][S_AXIS_FIFO_37_DMWIDTH/8-1:0] = s_axis_fifo_37_tstrb;
            assign tdata[37][S_AXIS_FIFO_37_DMWIDTH-1:0] = s_axis_fifo_37_tdata;
            assign s_axis_fifo_37_tready = tready[37];
            assign ap_fifo_iarg_37_empty_n = empty[37];
            assign ap_fifo_iarg_37_dout = dout[37][S_AXIS_FIFO_37_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 38) begin
            assign axis_clk[38] = s_axis_fifo_38_aclk;
            assign axis_rst[38] = s_axis_fifo_38_aresetn;
            assign tlast[38] = s_axis_fifo_38_tlast;
            assign tvalid[38] = s_axis_fifo_38_tvalid;
            assign read[38] = ap_fifo_iarg_38_read;
            assign tkeep[38][S_AXIS_FIFO_38_DMWIDTH/8-1:0] = s_axis_fifo_38_tkeep;
            assign tstrb[38][S_AXIS_FIFO_38_DMWIDTH/8-1:0] = s_axis_fifo_38_tstrb;
            assign tdata[38][S_AXIS_FIFO_38_DMWIDTH-1:0] = s_axis_fifo_38_tdata;
            assign s_axis_fifo_38_tready = tready[38];
            assign ap_fifo_iarg_38_empty_n = empty[38];
            assign ap_fifo_iarg_38_dout = dout[38][S_AXIS_FIFO_38_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 39) begin
            assign axis_clk[39] = s_axis_fifo_39_aclk;
            assign axis_rst[39] = s_axis_fifo_39_aresetn;
            assign tlast[39] = s_axis_fifo_39_tlast;
            assign tvalid[39] = s_axis_fifo_39_tvalid;
            assign read[39] = ap_fifo_iarg_39_read;
            assign tkeep[39][S_AXIS_FIFO_39_DMWIDTH/8-1:0] = s_axis_fifo_39_tkeep;
            assign tstrb[39][S_AXIS_FIFO_39_DMWIDTH/8-1:0] = s_axis_fifo_39_tstrb;
            assign tdata[39][S_AXIS_FIFO_39_DMWIDTH-1:0] = s_axis_fifo_39_tdata;
            assign s_axis_fifo_39_tready = tready[39];
            assign ap_fifo_iarg_39_empty_n = empty[39];
            assign ap_fifo_iarg_39_dout = dout[39][S_AXIS_FIFO_39_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 40) begin
            assign axis_clk[40] = s_axis_fifo_40_aclk;
            assign axis_rst[40] = s_axis_fifo_40_aresetn;
            assign tlast[40] = s_axis_fifo_40_tlast;
            assign tvalid[40] = s_axis_fifo_40_tvalid;
            assign read[40] = ap_fifo_iarg_40_read;
            assign tkeep[40][S_AXIS_FIFO_40_DMWIDTH/8-1:0] = s_axis_fifo_40_tkeep;
            assign tstrb[40][S_AXIS_FIFO_40_DMWIDTH/8-1:0] = s_axis_fifo_40_tstrb;
            assign tdata[40][S_AXIS_FIFO_40_DMWIDTH-1:0] = s_axis_fifo_40_tdata;
            assign s_axis_fifo_40_tready = tready[40];
            assign ap_fifo_iarg_40_empty_n = empty[40];
            assign ap_fifo_iarg_40_dout = dout[40][S_AXIS_FIFO_40_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 41) begin
            assign axis_clk[41] = s_axis_fifo_41_aclk;
            assign axis_rst[41] = s_axis_fifo_41_aresetn;
            assign tlast[41] = s_axis_fifo_41_tlast;
            assign tvalid[41] = s_axis_fifo_41_tvalid;
            assign read[41] = ap_fifo_iarg_41_read;
            assign tkeep[41][S_AXIS_FIFO_41_DMWIDTH/8-1:0] = s_axis_fifo_41_tkeep;
            assign tstrb[41][S_AXIS_FIFO_41_DMWIDTH/8-1:0] = s_axis_fifo_41_tstrb;
            assign tdata[41][S_AXIS_FIFO_41_DMWIDTH-1:0] = s_axis_fifo_41_tdata;
            assign s_axis_fifo_41_tready = tready[41];
            assign ap_fifo_iarg_41_empty_n = empty[41];
            assign ap_fifo_iarg_41_dout = dout[41][S_AXIS_FIFO_41_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 42) begin
            assign axis_clk[42] = s_axis_fifo_42_aclk;
            assign axis_rst[42] = s_axis_fifo_42_aresetn;
            assign tlast[42] = s_axis_fifo_42_tlast;
            assign tvalid[42] = s_axis_fifo_42_tvalid;
            assign read[42] = ap_fifo_iarg_42_read;
            assign tkeep[42][S_AXIS_FIFO_42_DMWIDTH/8-1:0] = s_axis_fifo_42_tkeep;
            assign tstrb[42][S_AXIS_FIFO_42_DMWIDTH/8-1:0] = s_axis_fifo_42_tstrb;
            assign tdata[42][S_AXIS_FIFO_42_DMWIDTH-1:0] = s_axis_fifo_42_tdata;
            assign s_axis_fifo_42_tready = tready[42];
            assign ap_fifo_iarg_42_empty_n = empty[42];
            assign ap_fifo_iarg_42_dout = dout[42][S_AXIS_FIFO_42_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 43) begin
            assign axis_clk[43] = s_axis_fifo_43_aclk;
            assign axis_rst[43] = s_axis_fifo_43_aresetn;
            assign tlast[43] = s_axis_fifo_43_tlast;
            assign tvalid[43] = s_axis_fifo_43_tvalid;
            assign read[43] = ap_fifo_iarg_43_read;
            assign tkeep[43][S_AXIS_FIFO_43_DMWIDTH/8-1:0] = s_axis_fifo_43_tkeep;
            assign tstrb[43][S_AXIS_FIFO_43_DMWIDTH/8-1:0] = s_axis_fifo_43_tstrb;
            assign tdata[43][S_AXIS_FIFO_43_DMWIDTH-1:0] = s_axis_fifo_43_tdata;
            assign s_axis_fifo_43_tready = tready[43];
            assign ap_fifo_iarg_43_empty_n = empty[43];
            assign ap_fifo_iarg_43_dout = dout[43][S_AXIS_FIFO_43_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 44) begin
            assign axis_clk[44] = s_axis_fifo_44_aclk;
            assign axis_rst[44] = s_axis_fifo_44_aresetn;
            assign tlast[44] = s_axis_fifo_44_tlast;
            assign tvalid[44] = s_axis_fifo_44_tvalid;
            assign read[44] = ap_fifo_iarg_44_read;
            assign tkeep[44][S_AXIS_FIFO_44_DMWIDTH/8-1:0] = s_axis_fifo_44_tkeep;
            assign tstrb[44][S_AXIS_FIFO_44_DMWIDTH/8-1:0] = s_axis_fifo_44_tstrb;
            assign tdata[44][S_AXIS_FIFO_44_DMWIDTH-1:0] = s_axis_fifo_44_tdata;
            assign s_axis_fifo_44_tready = tready[44];
            assign ap_fifo_iarg_44_empty_n = empty[44];
            assign ap_fifo_iarg_44_dout = dout[44][S_AXIS_FIFO_44_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 45) begin
            assign axis_clk[45] = s_axis_fifo_45_aclk;
            assign axis_rst[45] = s_axis_fifo_45_aresetn;
            assign tlast[45] = s_axis_fifo_45_tlast;
            assign tvalid[45] = s_axis_fifo_45_tvalid;
            assign read[45] = ap_fifo_iarg_45_read;
            assign tkeep[45][S_AXIS_FIFO_45_DMWIDTH/8-1:0] = s_axis_fifo_45_tkeep;
            assign tstrb[45][S_AXIS_FIFO_45_DMWIDTH/8-1:0] = s_axis_fifo_45_tstrb;
            assign tdata[45][S_AXIS_FIFO_45_DMWIDTH-1:0] = s_axis_fifo_45_tdata;
            assign s_axis_fifo_45_tready = tready[45];
            assign ap_fifo_iarg_45_empty_n = empty[45];
            assign ap_fifo_iarg_45_dout = dout[45][S_AXIS_FIFO_45_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 46) begin
            assign axis_clk[46] = s_axis_fifo_46_aclk;
            assign axis_rst[46] = s_axis_fifo_46_aresetn;
            assign tlast[46] = s_axis_fifo_46_tlast;
            assign tvalid[46] = s_axis_fifo_46_tvalid;
            assign read[46] = ap_fifo_iarg_46_read;
            assign tkeep[46][S_AXIS_FIFO_46_DMWIDTH/8-1:0] = s_axis_fifo_46_tkeep;
            assign tstrb[46][S_AXIS_FIFO_46_DMWIDTH/8-1:0] = s_axis_fifo_46_tstrb;
            assign tdata[46][S_AXIS_FIFO_46_DMWIDTH-1:0] = s_axis_fifo_46_tdata;
            assign s_axis_fifo_46_tready = tready[46];
            assign ap_fifo_iarg_46_empty_n = empty[46];
            assign ap_fifo_iarg_46_dout = dout[46][S_AXIS_FIFO_46_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 47) begin
            assign axis_clk[47] = s_axis_fifo_47_aclk;
            assign axis_rst[47] = s_axis_fifo_47_aresetn;
            assign tlast[47] = s_axis_fifo_47_tlast;
            assign tvalid[47] = s_axis_fifo_47_tvalid;
            assign read[47] = ap_fifo_iarg_47_read;
            assign tkeep[47][S_AXIS_FIFO_47_DMWIDTH/8-1:0] = s_axis_fifo_47_tkeep;
            assign tstrb[47][S_AXIS_FIFO_47_DMWIDTH/8-1:0] = s_axis_fifo_47_tstrb;
            assign tdata[47][S_AXIS_FIFO_47_DMWIDTH-1:0] = s_axis_fifo_47_tdata;
            assign s_axis_fifo_47_tready = tready[47];
            assign ap_fifo_iarg_47_empty_n = empty[47];
            assign ap_fifo_iarg_47_dout = dout[47][S_AXIS_FIFO_47_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 48) begin
            assign axis_clk[48] = s_axis_fifo_48_aclk;
            assign axis_rst[48] = s_axis_fifo_48_aresetn;
            assign tlast[48] = s_axis_fifo_48_tlast;
            assign tvalid[48] = s_axis_fifo_48_tvalid;
            assign read[48] = ap_fifo_iarg_48_read;
            assign tkeep[48][S_AXIS_FIFO_48_DMWIDTH/8-1:0] = s_axis_fifo_48_tkeep;
            assign tstrb[48][S_AXIS_FIFO_48_DMWIDTH/8-1:0] = s_axis_fifo_48_tstrb;
            assign tdata[48][S_AXIS_FIFO_48_DMWIDTH-1:0] = s_axis_fifo_48_tdata;
            assign s_axis_fifo_48_tready = tready[48];
            assign ap_fifo_iarg_48_empty_n = empty[48];
            assign ap_fifo_iarg_48_dout = dout[48][S_AXIS_FIFO_48_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 49) begin
            assign axis_clk[49] = s_axis_fifo_49_aclk;
            assign axis_rst[49] = s_axis_fifo_49_aresetn;
            assign tlast[49] = s_axis_fifo_49_tlast;
            assign tvalid[49] = s_axis_fifo_49_tvalid;
            assign read[49] = ap_fifo_iarg_49_read;
            assign tkeep[49][S_AXIS_FIFO_49_DMWIDTH/8-1:0] = s_axis_fifo_49_tkeep;
            assign tstrb[49][S_AXIS_FIFO_49_DMWIDTH/8-1:0] = s_axis_fifo_49_tstrb;
            assign tdata[49][S_AXIS_FIFO_49_DMWIDTH-1:0] = s_axis_fifo_49_tdata;
            assign s_axis_fifo_49_tready = tready[49];
            assign ap_fifo_iarg_49_empty_n = empty[49];
            assign ap_fifo_iarg_49_dout = dout[49][S_AXIS_FIFO_49_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 50) begin
            assign axis_clk[50] = s_axis_fifo_50_aclk;
            assign axis_rst[50] = s_axis_fifo_50_aresetn;
            assign tlast[50] = s_axis_fifo_50_tlast;
            assign tvalid[50] = s_axis_fifo_50_tvalid;
            assign read[50] = ap_fifo_iarg_50_read;
            assign tkeep[50][S_AXIS_FIFO_50_DMWIDTH/8-1:0] = s_axis_fifo_50_tkeep;
            assign tstrb[50][S_AXIS_FIFO_50_DMWIDTH/8-1:0] = s_axis_fifo_50_tstrb;
            assign tdata[50][S_AXIS_FIFO_50_DMWIDTH-1:0] = s_axis_fifo_50_tdata;
            assign s_axis_fifo_50_tready = tready[50];
            assign ap_fifo_iarg_50_empty_n = empty[50];
            assign ap_fifo_iarg_50_dout = dout[50][S_AXIS_FIFO_50_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 51) begin
            assign axis_clk[51] = s_axis_fifo_51_aclk;
            assign axis_rst[51] = s_axis_fifo_51_aresetn;
            assign tlast[51] = s_axis_fifo_51_tlast;
            assign tvalid[51] = s_axis_fifo_51_tvalid;
            assign read[51] = ap_fifo_iarg_51_read;
            assign tkeep[51][S_AXIS_FIFO_51_DMWIDTH/8-1:0] = s_axis_fifo_51_tkeep;
            assign tstrb[51][S_AXIS_FIFO_51_DMWIDTH/8-1:0] = s_axis_fifo_51_tstrb;
            assign tdata[51][S_AXIS_FIFO_51_DMWIDTH-1:0] = s_axis_fifo_51_tdata;
            assign s_axis_fifo_51_tready = tready[51];
            assign ap_fifo_iarg_51_empty_n = empty[51];
            assign ap_fifo_iarg_51_dout = dout[51][S_AXIS_FIFO_51_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 52) begin
            assign axis_clk[52] = s_axis_fifo_52_aclk;
            assign axis_rst[52] = s_axis_fifo_52_aresetn;
            assign tlast[52] = s_axis_fifo_52_tlast;
            assign tvalid[52] = s_axis_fifo_52_tvalid;
            assign read[52] = ap_fifo_iarg_52_read;
            assign tkeep[52][S_AXIS_FIFO_52_DMWIDTH/8-1:0] = s_axis_fifo_52_tkeep;
            assign tstrb[52][S_AXIS_FIFO_52_DMWIDTH/8-1:0] = s_axis_fifo_52_tstrb;
            assign tdata[52][S_AXIS_FIFO_52_DMWIDTH-1:0] = s_axis_fifo_52_tdata;
            assign s_axis_fifo_52_tready = tready[52];
            assign ap_fifo_iarg_52_empty_n = empty[52];
            assign ap_fifo_iarg_52_dout = dout[52][S_AXIS_FIFO_52_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 53) begin
            assign axis_clk[53] = s_axis_fifo_53_aclk;
            assign axis_rst[53] = s_axis_fifo_53_aresetn;
            assign tlast[53] = s_axis_fifo_53_tlast;
            assign tvalid[53] = s_axis_fifo_53_tvalid;
            assign read[53] = ap_fifo_iarg_53_read;
            assign tkeep[53][S_AXIS_FIFO_53_DMWIDTH/8-1:0] = s_axis_fifo_53_tkeep;
            assign tstrb[53][S_AXIS_FIFO_53_DMWIDTH/8-1:0] = s_axis_fifo_53_tstrb;
            assign tdata[53][S_AXIS_FIFO_53_DMWIDTH-1:0] = s_axis_fifo_53_tdata;
            assign s_axis_fifo_53_tready = tready[53];
            assign ap_fifo_iarg_53_empty_n = empty[53];
            assign ap_fifo_iarg_53_dout = dout[53][S_AXIS_FIFO_53_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 54) begin
            assign axis_clk[54] = s_axis_fifo_54_aclk;
            assign axis_rst[54] = s_axis_fifo_54_aresetn;
            assign tlast[54] = s_axis_fifo_54_tlast;
            assign tvalid[54] = s_axis_fifo_54_tvalid;
            assign read[54] = ap_fifo_iarg_54_read;
            assign tkeep[54][S_AXIS_FIFO_54_DMWIDTH/8-1:0] = s_axis_fifo_54_tkeep;
            assign tstrb[54][S_AXIS_FIFO_54_DMWIDTH/8-1:0] = s_axis_fifo_54_tstrb;
            assign tdata[54][S_AXIS_FIFO_54_DMWIDTH-1:0] = s_axis_fifo_54_tdata;
            assign s_axis_fifo_54_tready = tready[54];
            assign ap_fifo_iarg_54_empty_n = empty[54];
            assign ap_fifo_iarg_54_dout = dout[54][S_AXIS_FIFO_54_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 55) begin
            assign axis_clk[55] = s_axis_fifo_55_aclk;
            assign axis_rst[55] = s_axis_fifo_55_aresetn;
            assign tlast[55] = s_axis_fifo_55_tlast;
            assign tvalid[55] = s_axis_fifo_55_tvalid;
            assign read[55] = ap_fifo_iarg_55_read;
            assign tkeep[55][S_AXIS_FIFO_55_DMWIDTH/8-1:0] = s_axis_fifo_55_tkeep;
            assign tstrb[55][S_AXIS_FIFO_55_DMWIDTH/8-1:0] = s_axis_fifo_55_tstrb;
            assign tdata[55][S_AXIS_FIFO_55_DMWIDTH-1:0] = s_axis_fifo_55_tdata;
            assign s_axis_fifo_55_tready = tready[55];
            assign ap_fifo_iarg_55_empty_n = empty[55];
            assign ap_fifo_iarg_55_dout = dout[55][S_AXIS_FIFO_55_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 56) begin
            assign axis_clk[56] = s_axis_fifo_56_aclk;
            assign axis_rst[56] = s_axis_fifo_56_aresetn;
            assign tlast[56] = s_axis_fifo_56_tlast;
            assign tvalid[56] = s_axis_fifo_56_tvalid;
            assign read[56] = ap_fifo_iarg_56_read;
            assign tkeep[56][S_AXIS_FIFO_56_DMWIDTH/8-1:0] = s_axis_fifo_56_tkeep;
            assign tstrb[56][S_AXIS_FIFO_56_DMWIDTH/8-1:0] = s_axis_fifo_56_tstrb;
            assign tdata[56][S_AXIS_FIFO_56_DMWIDTH-1:0] = s_axis_fifo_56_tdata;
            assign s_axis_fifo_56_tready = tready[56];
            assign ap_fifo_iarg_56_empty_n = empty[56];
            assign ap_fifo_iarg_56_dout = dout[56][S_AXIS_FIFO_56_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 57) begin
            assign axis_clk[57] = s_axis_fifo_57_aclk;
            assign axis_rst[57] = s_axis_fifo_57_aresetn;
            assign tlast[57] = s_axis_fifo_57_tlast;
            assign tvalid[57] = s_axis_fifo_57_tvalid;
            assign read[57] = ap_fifo_iarg_57_read;
            assign tkeep[57][S_AXIS_FIFO_57_DMWIDTH/8-1:0] = s_axis_fifo_57_tkeep;
            assign tstrb[57][S_AXIS_FIFO_57_DMWIDTH/8-1:0] = s_axis_fifo_57_tstrb;
            assign tdata[57][S_AXIS_FIFO_57_DMWIDTH-1:0] = s_axis_fifo_57_tdata;
            assign s_axis_fifo_57_tready = tready[57];
            assign ap_fifo_iarg_57_empty_n = empty[57];
            assign ap_fifo_iarg_57_dout = dout[57][S_AXIS_FIFO_57_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 58) begin
            assign axis_clk[58] = s_axis_fifo_58_aclk;
            assign axis_rst[58] = s_axis_fifo_58_aresetn;
            assign tlast[58] = s_axis_fifo_58_tlast;
            assign tvalid[58] = s_axis_fifo_58_tvalid;
            assign read[58] = ap_fifo_iarg_58_read;
            assign tkeep[58][S_AXIS_FIFO_58_DMWIDTH/8-1:0] = s_axis_fifo_58_tkeep;
            assign tstrb[58][S_AXIS_FIFO_58_DMWIDTH/8-1:0] = s_axis_fifo_58_tstrb;
            assign tdata[58][S_AXIS_FIFO_58_DMWIDTH-1:0] = s_axis_fifo_58_tdata;
            assign s_axis_fifo_58_tready = tready[58];
            assign ap_fifo_iarg_58_empty_n = empty[58];
            assign ap_fifo_iarg_58_dout = dout[58][S_AXIS_FIFO_58_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 59) begin
            assign axis_clk[59] = s_axis_fifo_59_aclk;
            assign axis_rst[59] = s_axis_fifo_59_aresetn;
            assign tlast[59] = s_axis_fifo_59_tlast;
            assign tvalid[59] = s_axis_fifo_59_tvalid;
            assign read[59] = ap_fifo_iarg_59_read;
            assign tkeep[59][S_AXIS_FIFO_59_DMWIDTH/8-1:0] = s_axis_fifo_59_tkeep;
            assign tstrb[59][S_AXIS_FIFO_59_DMWIDTH/8-1:0] = s_axis_fifo_59_tstrb;
            assign tdata[59][S_AXIS_FIFO_59_DMWIDTH-1:0] = s_axis_fifo_59_tdata;
            assign s_axis_fifo_59_tready = tready[59];
            assign ap_fifo_iarg_59_empty_n = empty[59];
            assign ap_fifo_iarg_59_dout = dout[59][S_AXIS_FIFO_59_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 60) begin
            assign axis_clk[60] = s_axis_fifo_60_aclk;
            assign axis_rst[60] = s_axis_fifo_60_aresetn;
            assign tlast[60] = s_axis_fifo_60_tlast;
            assign tvalid[60] = s_axis_fifo_60_tvalid;
            assign read[60] = ap_fifo_iarg_60_read;
            assign tkeep[60][S_AXIS_FIFO_60_DMWIDTH/8-1:0] = s_axis_fifo_60_tkeep;
            assign tstrb[60][S_AXIS_FIFO_60_DMWIDTH/8-1:0] = s_axis_fifo_60_tstrb;
            assign tdata[60][S_AXIS_FIFO_60_DMWIDTH-1:0] = s_axis_fifo_60_tdata;
            assign s_axis_fifo_60_tready = tready[60];
            assign ap_fifo_iarg_60_empty_n = empty[60];
            assign ap_fifo_iarg_60_dout = dout[60][S_AXIS_FIFO_60_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 61) begin
            assign axis_clk[61] = s_axis_fifo_61_aclk;
            assign axis_rst[61] = s_axis_fifo_61_aresetn;
            assign tlast[61] = s_axis_fifo_61_tlast;
            assign tvalid[61] = s_axis_fifo_61_tvalid;
            assign read[61] = ap_fifo_iarg_61_read;
            assign tkeep[61][S_AXIS_FIFO_61_DMWIDTH/8-1:0] = s_axis_fifo_61_tkeep;
            assign tstrb[61][S_AXIS_FIFO_61_DMWIDTH/8-1:0] = s_axis_fifo_61_tstrb;
            assign tdata[61][S_AXIS_FIFO_61_DMWIDTH-1:0] = s_axis_fifo_61_tdata;
            assign s_axis_fifo_61_tready = tready[61];
            assign ap_fifo_iarg_61_empty_n = empty[61];
            assign ap_fifo_iarg_61_dout = dout[61][S_AXIS_FIFO_61_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 62) begin
            assign axis_clk[62] = s_axis_fifo_62_aclk;
            assign axis_rst[62] = s_axis_fifo_62_aresetn;
            assign tlast[62] = s_axis_fifo_62_tlast;
            assign tvalid[62] = s_axis_fifo_62_tvalid;
            assign read[62] = ap_fifo_iarg_62_read;
            assign tkeep[62][S_AXIS_FIFO_62_DMWIDTH/8-1:0] = s_axis_fifo_62_tkeep;
            assign tstrb[62][S_AXIS_FIFO_62_DMWIDTH/8-1:0] = s_axis_fifo_62_tstrb;
            assign tdata[62][S_AXIS_FIFO_62_DMWIDTH-1:0] = s_axis_fifo_62_tdata;
            assign s_axis_fifo_62_tready = tready[62];
            assign ap_fifo_iarg_62_empty_n = empty[62];
            assign ap_fifo_iarg_62_dout = dout[62][S_AXIS_FIFO_62_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 63) begin
            assign axis_clk[63] = s_axis_fifo_63_aclk;
            assign axis_rst[63] = s_axis_fifo_63_aresetn;
            assign tlast[63] = s_axis_fifo_63_tlast;
            assign tvalid[63] = s_axis_fifo_63_tvalid;
            assign read[63] = ap_fifo_iarg_63_read;
            assign tkeep[63][S_AXIS_FIFO_63_DMWIDTH/8-1:0] = s_axis_fifo_63_tkeep;
            assign tstrb[63][S_AXIS_FIFO_63_DMWIDTH/8-1:0] = s_axis_fifo_63_tstrb;
            assign tdata[63][S_AXIS_FIFO_63_DMWIDTH-1:0] = s_axis_fifo_63_tdata;
            assign s_axis_fifo_63_tready = tready[63];
            assign ap_fifo_iarg_63_empty_n = empty[63];
            assign ap_fifo_iarg_63_dout = dout[63][S_AXIS_FIFO_63_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 64) begin
            assign axis_clk[64] = s_axis_fifo_64_aclk;
            assign axis_rst[64] = s_axis_fifo_64_aresetn;
            assign tlast[64] = s_axis_fifo_64_tlast;
            assign tvalid[64] = s_axis_fifo_64_tvalid;
            assign read[64] = ap_fifo_iarg_64_read;
            assign tkeep[64][S_AXIS_FIFO_64_DMWIDTH/8-1:0] = s_axis_fifo_64_tkeep;
            assign tstrb[64][S_AXIS_FIFO_64_DMWIDTH/8-1:0] = s_axis_fifo_64_tstrb;
            assign tdata[64][S_AXIS_FIFO_64_DMWIDTH-1:0] = s_axis_fifo_64_tdata;
            assign s_axis_fifo_64_tready = tready[64];
            assign ap_fifo_iarg_64_empty_n = empty[64];
            assign ap_fifo_iarg_64_dout = dout[64][S_AXIS_FIFO_64_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 65) begin
            assign axis_clk[65] = s_axis_fifo_65_aclk;
            assign axis_rst[65] = s_axis_fifo_65_aresetn;
            assign tlast[65] = s_axis_fifo_65_tlast;
            assign tvalid[65] = s_axis_fifo_65_tvalid;
            assign read[65] = ap_fifo_iarg_65_read;
            assign tkeep[65][S_AXIS_FIFO_65_DMWIDTH/8-1:0] = s_axis_fifo_65_tkeep;
            assign tstrb[65][S_AXIS_FIFO_65_DMWIDTH/8-1:0] = s_axis_fifo_65_tstrb;
            assign tdata[65][S_AXIS_FIFO_65_DMWIDTH-1:0] = s_axis_fifo_65_tdata;
            assign s_axis_fifo_65_tready = tready[65];
            assign ap_fifo_iarg_65_empty_n = empty[65];
            assign ap_fifo_iarg_65_dout = dout[65][S_AXIS_FIFO_65_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 66) begin
            assign axis_clk[66] = s_axis_fifo_66_aclk;
            assign axis_rst[66] = s_axis_fifo_66_aresetn;
            assign tlast[66] = s_axis_fifo_66_tlast;
            assign tvalid[66] = s_axis_fifo_66_tvalid;
            assign read[66] = ap_fifo_iarg_66_read;
            assign tkeep[66][S_AXIS_FIFO_66_DMWIDTH/8-1:0] = s_axis_fifo_66_tkeep;
            assign tstrb[66][S_AXIS_FIFO_66_DMWIDTH/8-1:0] = s_axis_fifo_66_tstrb;
            assign tdata[66][S_AXIS_FIFO_66_DMWIDTH-1:0] = s_axis_fifo_66_tdata;
            assign s_axis_fifo_66_tready = tready[66];
            assign ap_fifo_iarg_66_empty_n = empty[66];
            assign ap_fifo_iarg_66_dout = dout[66][S_AXIS_FIFO_66_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 67) begin
            assign axis_clk[67] = s_axis_fifo_67_aclk;
            assign axis_rst[67] = s_axis_fifo_67_aresetn;
            assign tlast[67] = s_axis_fifo_67_tlast;
            assign tvalid[67] = s_axis_fifo_67_tvalid;
            assign read[67] = ap_fifo_iarg_67_read;
            assign tkeep[67][S_AXIS_FIFO_67_DMWIDTH/8-1:0] = s_axis_fifo_67_tkeep;
            assign tstrb[67][S_AXIS_FIFO_67_DMWIDTH/8-1:0] = s_axis_fifo_67_tstrb;
            assign tdata[67][S_AXIS_FIFO_67_DMWIDTH-1:0] = s_axis_fifo_67_tdata;
            assign s_axis_fifo_67_tready = tready[67];
            assign ap_fifo_iarg_67_empty_n = empty[67];
            assign ap_fifo_iarg_67_dout = dout[67][S_AXIS_FIFO_67_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 68) begin
            assign axis_clk[68] = s_axis_fifo_68_aclk;
            assign axis_rst[68] = s_axis_fifo_68_aresetn;
            assign tlast[68] = s_axis_fifo_68_tlast;
            assign tvalid[68] = s_axis_fifo_68_tvalid;
            assign read[68] = ap_fifo_iarg_68_read;
            assign tkeep[68][S_AXIS_FIFO_68_DMWIDTH/8-1:0] = s_axis_fifo_68_tkeep;
            assign tstrb[68][S_AXIS_FIFO_68_DMWIDTH/8-1:0] = s_axis_fifo_68_tstrb;
            assign tdata[68][S_AXIS_FIFO_68_DMWIDTH-1:0] = s_axis_fifo_68_tdata;
            assign s_axis_fifo_68_tready = tready[68];
            assign ap_fifo_iarg_68_empty_n = empty[68];
            assign ap_fifo_iarg_68_dout = dout[68][S_AXIS_FIFO_68_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 69) begin
            assign axis_clk[69] = s_axis_fifo_69_aclk;
            assign axis_rst[69] = s_axis_fifo_69_aresetn;
            assign tlast[69] = s_axis_fifo_69_tlast;
            assign tvalid[69] = s_axis_fifo_69_tvalid;
            assign read[69] = ap_fifo_iarg_69_read;
            assign tkeep[69][S_AXIS_FIFO_69_DMWIDTH/8-1:0] = s_axis_fifo_69_tkeep;
            assign tstrb[69][S_AXIS_FIFO_69_DMWIDTH/8-1:0] = s_axis_fifo_69_tstrb;
            assign tdata[69][S_AXIS_FIFO_69_DMWIDTH-1:0] = s_axis_fifo_69_tdata;
            assign s_axis_fifo_69_tready = tready[69];
            assign ap_fifo_iarg_69_empty_n = empty[69];
            assign ap_fifo_iarg_69_dout = dout[69][S_AXIS_FIFO_69_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 70) begin
            assign axis_clk[70] = s_axis_fifo_70_aclk;
            assign axis_rst[70] = s_axis_fifo_70_aresetn;
            assign tlast[70] = s_axis_fifo_70_tlast;
            assign tvalid[70] = s_axis_fifo_70_tvalid;
            assign read[70] = ap_fifo_iarg_70_read;
            assign tkeep[70][S_AXIS_FIFO_70_DMWIDTH/8-1:0] = s_axis_fifo_70_tkeep;
            assign tstrb[70][S_AXIS_FIFO_70_DMWIDTH/8-1:0] = s_axis_fifo_70_tstrb;
            assign tdata[70][S_AXIS_FIFO_70_DMWIDTH-1:0] = s_axis_fifo_70_tdata;
            assign s_axis_fifo_70_tready = tready[70];
            assign ap_fifo_iarg_70_empty_n = empty[70];
            assign ap_fifo_iarg_70_dout = dout[70][S_AXIS_FIFO_70_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 71) begin
            assign axis_clk[71] = s_axis_fifo_71_aclk;
            assign axis_rst[71] = s_axis_fifo_71_aresetn;
            assign tlast[71] = s_axis_fifo_71_tlast;
            assign tvalid[71] = s_axis_fifo_71_tvalid;
            assign read[71] = ap_fifo_iarg_71_read;
            assign tkeep[71][S_AXIS_FIFO_71_DMWIDTH/8-1:0] = s_axis_fifo_71_tkeep;
            assign tstrb[71][S_AXIS_FIFO_71_DMWIDTH/8-1:0] = s_axis_fifo_71_tstrb;
            assign tdata[71][S_AXIS_FIFO_71_DMWIDTH-1:0] = s_axis_fifo_71_tdata;
            assign s_axis_fifo_71_tready = tready[71];
            assign ap_fifo_iarg_71_empty_n = empty[71];
            assign ap_fifo_iarg_71_dout = dout[71][S_AXIS_FIFO_71_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 72) begin
            assign axis_clk[72] = s_axis_fifo_72_aclk;
            assign axis_rst[72] = s_axis_fifo_72_aresetn;
            assign tlast[72] = s_axis_fifo_72_tlast;
            assign tvalid[72] = s_axis_fifo_72_tvalid;
            assign read[72] = ap_fifo_iarg_72_read;
            assign tkeep[72][S_AXIS_FIFO_72_DMWIDTH/8-1:0] = s_axis_fifo_72_tkeep;
            assign tstrb[72][S_AXIS_FIFO_72_DMWIDTH/8-1:0] = s_axis_fifo_72_tstrb;
            assign tdata[72][S_AXIS_FIFO_72_DMWIDTH-1:0] = s_axis_fifo_72_tdata;
            assign s_axis_fifo_72_tready = tready[72];
            assign ap_fifo_iarg_72_empty_n = empty[72];
            assign ap_fifo_iarg_72_dout = dout[72][S_AXIS_FIFO_72_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 73) begin
            assign axis_clk[73] = s_axis_fifo_73_aclk;
            assign axis_rst[73] = s_axis_fifo_73_aresetn;
            assign tlast[73] = s_axis_fifo_73_tlast;
            assign tvalid[73] = s_axis_fifo_73_tvalid;
            assign read[73] = ap_fifo_iarg_73_read;
            assign tkeep[73][S_AXIS_FIFO_73_DMWIDTH/8-1:0] = s_axis_fifo_73_tkeep;
            assign tstrb[73][S_AXIS_FIFO_73_DMWIDTH/8-1:0] = s_axis_fifo_73_tstrb;
            assign tdata[73][S_AXIS_FIFO_73_DMWIDTH-1:0] = s_axis_fifo_73_tdata;
            assign s_axis_fifo_73_tready = tready[73];
            assign ap_fifo_iarg_73_empty_n = empty[73];
            assign ap_fifo_iarg_73_dout = dout[73][S_AXIS_FIFO_73_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 74) begin
            assign axis_clk[74] = s_axis_fifo_74_aclk;
            assign axis_rst[74] = s_axis_fifo_74_aresetn;
            assign tlast[74] = s_axis_fifo_74_tlast;
            assign tvalid[74] = s_axis_fifo_74_tvalid;
            assign read[74] = ap_fifo_iarg_74_read;
            assign tkeep[74][S_AXIS_FIFO_74_DMWIDTH/8-1:0] = s_axis_fifo_74_tkeep;
            assign tstrb[74][S_AXIS_FIFO_74_DMWIDTH/8-1:0] = s_axis_fifo_74_tstrb;
            assign tdata[74][S_AXIS_FIFO_74_DMWIDTH-1:0] = s_axis_fifo_74_tdata;
            assign s_axis_fifo_74_tready = tready[74];
            assign ap_fifo_iarg_74_empty_n = empty[74];
            assign ap_fifo_iarg_74_dout = dout[74][S_AXIS_FIFO_74_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 75) begin
            assign axis_clk[75] = s_axis_fifo_75_aclk;
            assign axis_rst[75] = s_axis_fifo_75_aresetn;
            assign tlast[75] = s_axis_fifo_75_tlast;
            assign tvalid[75] = s_axis_fifo_75_tvalid;
            assign read[75] = ap_fifo_iarg_75_read;
            assign tkeep[75][S_AXIS_FIFO_75_DMWIDTH/8-1:0] = s_axis_fifo_75_tkeep;
            assign tstrb[75][S_AXIS_FIFO_75_DMWIDTH/8-1:0] = s_axis_fifo_75_tstrb;
            assign tdata[75][S_AXIS_FIFO_75_DMWIDTH-1:0] = s_axis_fifo_75_tdata;
            assign s_axis_fifo_75_tready = tready[75];
            assign ap_fifo_iarg_75_empty_n = empty[75];
            assign ap_fifo_iarg_75_dout = dout[75][S_AXIS_FIFO_75_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 76) begin
            assign axis_clk[76] = s_axis_fifo_76_aclk;
            assign axis_rst[76] = s_axis_fifo_76_aresetn;
            assign tlast[76] = s_axis_fifo_76_tlast;
            assign tvalid[76] = s_axis_fifo_76_tvalid;
            assign read[76] = ap_fifo_iarg_76_read;
            assign tkeep[76][S_AXIS_FIFO_76_DMWIDTH/8-1:0] = s_axis_fifo_76_tkeep;
            assign tstrb[76][S_AXIS_FIFO_76_DMWIDTH/8-1:0] = s_axis_fifo_76_tstrb;
            assign tdata[76][S_AXIS_FIFO_76_DMWIDTH-1:0] = s_axis_fifo_76_tdata;
            assign s_axis_fifo_76_tready = tready[76];
            assign ap_fifo_iarg_76_empty_n = empty[76];
            assign ap_fifo_iarg_76_dout = dout[76][S_AXIS_FIFO_76_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 77) begin
            assign axis_clk[77] = s_axis_fifo_77_aclk;
            assign axis_rst[77] = s_axis_fifo_77_aresetn;
            assign tlast[77] = s_axis_fifo_77_tlast;
            assign tvalid[77] = s_axis_fifo_77_tvalid;
            assign read[77] = ap_fifo_iarg_77_read;
            assign tkeep[77][S_AXIS_FIFO_77_DMWIDTH/8-1:0] = s_axis_fifo_77_tkeep;
            assign tstrb[77][S_AXIS_FIFO_77_DMWIDTH/8-1:0] = s_axis_fifo_77_tstrb;
            assign tdata[77][S_AXIS_FIFO_77_DMWIDTH-1:0] = s_axis_fifo_77_tdata;
            assign s_axis_fifo_77_tready = tready[77];
            assign ap_fifo_iarg_77_empty_n = empty[77];
            assign ap_fifo_iarg_77_dout = dout[77][S_AXIS_FIFO_77_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 78) begin
            assign axis_clk[78] = s_axis_fifo_78_aclk;
            assign axis_rst[78] = s_axis_fifo_78_aresetn;
            assign tlast[78] = s_axis_fifo_78_tlast;
            assign tvalid[78] = s_axis_fifo_78_tvalid;
            assign read[78] = ap_fifo_iarg_78_read;
            assign tkeep[78][S_AXIS_FIFO_78_DMWIDTH/8-1:0] = s_axis_fifo_78_tkeep;
            assign tstrb[78][S_AXIS_FIFO_78_DMWIDTH/8-1:0] = s_axis_fifo_78_tstrb;
            assign tdata[78][S_AXIS_FIFO_78_DMWIDTH-1:0] = s_axis_fifo_78_tdata;
            assign s_axis_fifo_78_tready = tready[78];
            assign ap_fifo_iarg_78_empty_n = empty[78];
            assign ap_fifo_iarg_78_dout = dout[78][S_AXIS_FIFO_78_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 79) begin
            assign axis_clk[79] = s_axis_fifo_79_aclk;
            assign axis_rst[79] = s_axis_fifo_79_aresetn;
            assign tlast[79] = s_axis_fifo_79_tlast;
            assign tvalid[79] = s_axis_fifo_79_tvalid;
            assign read[79] = ap_fifo_iarg_79_read;
            assign tkeep[79][S_AXIS_FIFO_79_DMWIDTH/8-1:0] = s_axis_fifo_79_tkeep;
            assign tstrb[79][S_AXIS_FIFO_79_DMWIDTH/8-1:0] = s_axis_fifo_79_tstrb;
            assign tdata[79][S_AXIS_FIFO_79_DMWIDTH-1:0] = s_axis_fifo_79_tdata;
            assign s_axis_fifo_79_tready = tready[79];
            assign ap_fifo_iarg_79_empty_n = empty[79];
            assign ap_fifo_iarg_79_dout = dout[79][S_AXIS_FIFO_79_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 80) begin
            assign axis_clk[80] = s_axis_fifo_80_aclk;
            assign axis_rst[80] = s_axis_fifo_80_aresetn;
            assign tlast[80] = s_axis_fifo_80_tlast;
            assign tvalid[80] = s_axis_fifo_80_tvalid;
            assign read[80] = ap_fifo_iarg_80_read;
            assign tkeep[80][S_AXIS_FIFO_80_DMWIDTH/8-1:0] = s_axis_fifo_80_tkeep;
            assign tstrb[80][S_AXIS_FIFO_80_DMWIDTH/8-1:0] = s_axis_fifo_80_tstrb;
            assign tdata[80][S_AXIS_FIFO_80_DMWIDTH-1:0] = s_axis_fifo_80_tdata;
            assign s_axis_fifo_80_tready = tready[80];
            assign ap_fifo_iarg_80_empty_n = empty[80];
            assign ap_fifo_iarg_80_dout = dout[80][S_AXIS_FIFO_80_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 81) begin
            assign axis_clk[81] = s_axis_fifo_81_aclk;
            assign axis_rst[81] = s_axis_fifo_81_aresetn;
            assign tlast[81] = s_axis_fifo_81_tlast;
            assign tvalid[81] = s_axis_fifo_81_tvalid;
            assign read[81] = ap_fifo_iarg_81_read;
            assign tkeep[81][S_AXIS_FIFO_81_DMWIDTH/8-1:0] = s_axis_fifo_81_tkeep;
            assign tstrb[81][S_AXIS_FIFO_81_DMWIDTH/8-1:0] = s_axis_fifo_81_tstrb;
            assign tdata[81][S_AXIS_FIFO_81_DMWIDTH-1:0] = s_axis_fifo_81_tdata;
            assign s_axis_fifo_81_tready = tready[81];
            assign ap_fifo_iarg_81_empty_n = empty[81];
            assign ap_fifo_iarg_81_dout = dout[81][S_AXIS_FIFO_81_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 82) begin
            assign axis_clk[82] = s_axis_fifo_82_aclk;
            assign axis_rst[82] = s_axis_fifo_82_aresetn;
            assign tlast[82] = s_axis_fifo_82_tlast;
            assign tvalid[82] = s_axis_fifo_82_tvalid;
            assign read[82] = ap_fifo_iarg_82_read;
            assign tkeep[82][S_AXIS_FIFO_82_DMWIDTH/8-1:0] = s_axis_fifo_82_tkeep;
            assign tstrb[82][S_AXIS_FIFO_82_DMWIDTH/8-1:0] = s_axis_fifo_82_tstrb;
            assign tdata[82][S_AXIS_FIFO_82_DMWIDTH-1:0] = s_axis_fifo_82_tdata;
            assign s_axis_fifo_82_tready = tready[82];
            assign ap_fifo_iarg_82_empty_n = empty[82];
            assign ap_fifo_iarg_82_dout = dout[82][S_AXIS_FIFO_82_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 83) begin
            assign axis_clk[83] = s_axis_fifo_83_aclk;
            assign axis_rst[83] = s_axis_fifo_83_aresetn;
            assign tlast[83] = s_axis_fifo_83_tlast;
            assign tvalid[83] = s_axis_fifo_83_tvalid;
            assign read[83] = ap_fifo_iarg_83_read;
            assign tkeep[83][S_AXIS_FIFO_83_DMWIDTH/8-1:0] = s_axis_fifo_83_tkeep;
            assign tstrb[83][S_AXIS_FIFO_83_DMWIDTH/8-1:0] = s_axis_fifo_83_tstrb;
            assign tdata[83][S_AXIS_FIFO_83_DMWIDTH-1:0] = s_axis_fifo_83_tdata;
            assign s_axis_fifo_83_tready = tready[83];
            assign ap_fifo_iarg_83_empty_n = empty[83];
            assign ap_fifo_iarg_83_dout = dout[83][S_AXIS_FIFO_83_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 84) begin
            assign axis_clk[84] = s_axis_fifo_84_aclk;
            assign axis_rst[84] = s_axis_fifo_84_aresetn;
            assign tlast[84] = s_axis_fifo_84_tlast;
            assign tvalid[84] = s_axis_fifo_84_tvalid;
            assign read[84] = ap_fifo_iarg_84_read;
            assign tkeep[84][S_AXIS_FIFO_84_DMWIDTH/8-1:0] = s_axis_fifo_84_tkeep;
            assign tstrb[84][S_AXIS_FIFO_84_DMWIDTH/8-1:0] = s_axis_fifo_84_tstrb;
            assign tdata[84][S_AXIS_FIFO_84_DMWIDTH-1:0] = s_axis_fifo_84_tdata;
            assign s_axis_fifo_84_tready = tready[84];
            assign ap_fifo_iarg_84_empty_n = empty[84];
            assign ap_fifo_iarg_84_dout = dout[84][S_AXIS_FIFO_84_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 85) begin
            assign axis_clk[85] = s_axis_fifo_85_aclk;
            assign axis_rst[85] = s_axis_fifo_85_aresetn;
            assign tlast[85] = s_axis_fifo_85_tlast;
            assign tvalid[85] = s_axis_fifo_85_tvalid;
            assign read[85] = ap_fifo_iarg_85_read;
            assign tkeep[85][S_AXIS_FIFO_85_DMWIDTH/8-1:0] = s_axis_fifo_85_tkeep;
            assign tstrb[85][S_AXIS_FIFO_85_DMWIDTH/8-1:0] = s_axis_fifo_85_tstrb;
            assign tdata[85][S_AXIS_FIFO_85_DMWIDTH-1:0] = s_axis_fifo_85_tdata;
            assign s_axis_fifo_85_tready = tready[85];
            assign ap_fifo_iarg_85_empty_n = empty[85];
            assign ap_fifo_iarg_85_dout = dout[85][S_AXIS_FIFO_85_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 86) begin
            assign axis_clk[86] = s_axis_fifo_86_aclk;
            assign axis_rst[86] = s_axis_fifo_86_aresetn;
            assign tlast[86] = s_axis_fifo_86_tlast;
            assign tvalid[86] = s_axis_fifo_86_tvalid;
            assign read[86] = ap_fifo_iarg_86_read;
            assign tkeep[86][S_AXIS_FIFO_86_DMWIDTH/8-1:0] = s_axis_fifo_86_tkeep;
            assign tstrb[86][S_AXIS_FIFO_86_DMWIDTH/8-1:0] = s_axis_fifo_86_tstrb;
            assign tdata[86][S_AXIS_FIFO_86_DMWIDTH-1:0] = s_axis_fifo_86_tdata;
            assign s_axis_fifo_86_tready = tready[86];
            assign ap_fifo_iarg_86_empty_n = empty[86];
            assign ap_fifo_iarg_86_dout = dout[86][S_AXIS_FIFO_86_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 87) begin
            assign axis_clk[87] = s_axis_fifo_87_aclk;
            assign axis_rst[87] = s_axis_fifo_87_aresetn;
            assign tlast[87] = s_axis_fifo_87_tlast;
            assign tvalid[87] = s_axis_fifo_87_tvalid;
            assign read[87] = ap_fifo_iarg_87_read;
            assign tkeep[87][S_AXIS_FIFO_87_DMWIDTH/8-1:0] = s_axis_fifo_87_tkeep;
            assign tstrb[87][S_AXIS_FIFO_87_DMWIDTH/8-1:0] = s_axis_fifo_87_tstrb;
            assign tdata[87][S_AXIS_FIFO_87_DMWIDTH-1:0] = s_axis_fifo_87_tdata;
            assign s_axis_fifo_87_tready = tready[87];
            assign ap_fifo_iarg_87_empty_n = empty[87];
            assign ap_fifo_iarg_87_dout = dout[87][S_AXIS_FIFO_87_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 88) begin
            assign axis_clk[88] = s_axis_fifo_88_aclk;
            assign axis_rst[88] = s_axis_fifo_88_aresetn;
            assign tlast[88] = s_axis_fifo_88_tlast;
            assign tvalid[88] = s_axis_fifo_88_tvalid;
            assign read[88] = ap_fifo_iarg_88_read;
            assign tkeep[88][S_AXIS_FIFO_88_DMWIDTH/8-1:0] = s_axis_fifo_88_tkeep;
            assign tstrb[88][S_AXIS_FIFO_88_DMWIDTH/8-1:0] = s_axis_fifo_88_tstrb;
            assign tdata[88][S_AXIS_FIFO_88_DMWIDTH-1:0] = s_axis_fifo_88_tdata;
            assign s_axis_fifo_88_tready = tready[88];
            assign ap_fifo_iarg_88_empty_n = empty[88];
            assign ap_fifo_iarg_88_dout = dout[88][S_AXIS_FIFO_88_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 89) begin
            assign axis_clk[89] = s_axis_fifo_89_aclk;
            assign axis_rst[89] = s_axis_fifo_89_aresetn;
            assign tlast[89] = s_axis_fifo_89_tlast;
            assign tvalid[89] = s_axis_fifo_89_tvalid;
            assign read[89] = ap_fifo_iarg_89_read;
            assign tkeep[89][S_AXIS_FIFO_89_DMWIDTH/8-1:0] = s_axis_fifo_89_tkeep;
            assign tstrb[89][S_AXIS_FIFO_89_DMWIDTH/8-1:0] = s_axis_fifo_89_tstrb;
            assign tdata[89][S_AXIS_FIFO_89_DMWIDTH-1:0] = s_axis_fifo_89_tdata;
            assign s_axis_fifo_89_tready = tready[89];
            assign ap_fifo_iarg_89_empty_n = empty[89];
            assign ap_fifo_iarg_89_dout = dout[89][S_AXIS_FIFO_89_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 90) begin
            assign axis_clk[90] = s_axis_fifo_90_aclk;
            assign axis_rst[90] = s_axis_fifo_90_aresetn;
            assign tlast[90] = s_axis_fifo_90_tlast;
            assign tvalid[90] = s_axis_fifo_90_tvalid;
            assign read[90] = ap_fifo_iarg_90_read;
            assign tkeep[90][S_AXIS_FIFO_90_DMWIDTH/8-1:0] = s_axis_fifo_90_tkeep;
            assign tstrb[90][S_AXIS_FIFO_90_DMWIDTH/8-1:0] = s_axis_fifo_90_tstrb;
            assign tdata[90][S_AXIS_FIFO_90_DMWIDTH-1:0] = s_axis_fifo_90_tdata;
            assign s_axis_fifo_90_tready = tready[90];
            assign ap_fifo_iarg_90_empty_n = empty[90];
            assign ap_fifo_iarg_90_dout = dout[90][S_AXIS_FIFO_90_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 91) begin
            assign axis_clk[91] = s_axis_fifo_91_aclk;
            assign axis_rst[91] = s_axis_fifo_91_aresetn;
            assign tlast[91] = s_axis_fifo_91_tlast;
            assign tvalid[91] = s_axis_fifo_91_tvalid;
            assign read[91] = ap_fifo_iarg_91_read;
            assign tkeep[91][S_AXIS_FIFO_91_DMWIDTH/8-1:0] = s_axis_fifo_91_tkeep;
            assign tstrb[91][S_AXIS_FIFO_91_DMWIDTH/8-1:0] = s_axis_fifo_91_tstrb;
            assign tdata[91][S_AXIS_FIFO_91_DMWIDTH-1:0] = s_axis_fifo_91_tdata;
            assign s_axis_fifo_91_tready = tready[91];
            assign ap_fifo_iarg_91_empty_n = empty[91];
            assign ap_fifo_iarg_91_dout = dout[91][S_AXIS_FIFO_91_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 92) begin
            assign axis_clk[92] = s_axis_fifo_92_aclk;
            assign axis_rst[92] = s_axis_fifo_92_aresetn;
            assign tlast[92] = s_axis_fifo_92_tlast;
            assign tvalid[92] = s_axis_fifo_92_tvalid;
            assign read[92] = ap_fifo_iarg_92_read;
            assign tkeep[92][S_AXIS_FIFO_92_DMWIDTH/8-1:0] = s_axis_fifo_92_tkeep;
            assign tstrb[92][S_AXIS_FIFO_92_DMWIDTH/8-1:0] = s_axis_fifo_92_tstrb;
            assign tdata[92][S_AXIS_FIFO_92_DMWIDTH-1:0] = s_axis_fifo_92_tdata;
            assign s_axis_fifo_92_tready = tready[92];
            assign ap_fifo_iarg_92_empty_n = empty[92];
            assign ap_fifo_iarg_92_dout = dout[92][S_AXIS_FIFO_92_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 93) begin
            assign axis_clk[93] = s_axis_fifo_93_aclk;
            assign axis_rst[93] = s_axis_fifo_93_aresetn;
            assign tlast[93] = s_axis_fifo_93_tlast;
            assign tvalid[93] = s_axis_fifo_93_tvalid;
            assign read[93] = ap_fifo_iarg_93_read;
            assign tkeep[93][S_AXIS_FIFO_93_DMWIDTH/8-1:0] = s_axis_fifo_93_tkeep;
            assign tstrb[93][S_AXIS_FIFO_93_DMWIDTH/8-1:0] = s_axis_fifo_93_tstrb;
            assign tdata[93][S_AXIS_FIFO_93_DMWIDTH-1:0] = s_axis_fifo_93_tdata;
            assign s_axis_fifo_93_tready = tready[93];
            assign ap_fifo_iarg_93_empty_n = empty[93];
            assign ap_fifo_iarg_93_dout = dout[93][S_AXIS_FIFO_93_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 94) begin
            assign axis_clk[94] = s_axis_fifo_94_aclk;
            assign axis_rst[94] = s_axis_fifo_94_aresetn;
            assign tlast[94] = s_axis_fifo_94_tlast;
            assign tvalid[94] = s_axis_fifo_94_tvalid;
            assign read[94] = ap_fifo_iarg_94_read;
            assign tkeep[94][S_AXIS_FIFO_94_DMWIDTH/8-1:0] = s_axis_fifo_94_tkeep;
            assign tstrb[94][S_AXIS_FIFO_94_DMWIDTH/8-1:0] = s_axis_fifo_94_tstrb;
            assign tdata[94][S_AXIS_FIFO_94_DMWIDTH-1:0] = s_axis_fifo_94_tdata;
            assign s_axis_fifo_94_tready = tready[94];
            assign ap_fifo_iarg_94_empty_n = empty[94];
            assign ap_fifo_iarg_94_dout = dout[94][S_AXIS_FIFO_94_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 95) begin
            assign axis_clk[95] = s_axis_fifo_95_aclk;
            assign axis_rst[95] = s_axis_fifo_95_aresetn;
            assign tlast[95] = s_axis_fifo_95_tlast;
            assign tvalid[95] = s_axis_fifo_95_tvalid;
            assign read[95] = ap_fifo_iarg_95_read;
            assign tkeep[95][S_AXIS_FIFO_95_DMWIDTH/8-1:0] = s_axis_fifo_95_tkeep;
            assign tstrb[95][S_AXIS_FIFO_95_DMWIDTH/8-1:0] = s_axis_fifo_95_tstrb;
            assign tdata[95][S_AXIS_FIFO_95_DMWIDTH-1:0] = s_axis_fifo_95_tdata;
            assign s_axis_fifo_95_tready = tready[95];
            assign ap_fifo_iarg_95_empty_n = empty[95];
            assign ap_fifo_iarg_95_dout = dout[95][S_AXIS_FIFO_95_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 96) begin
            assign axis_clk[96] = s_axis_fifo_96_aclk;
            assign axis_rst[96] = s_axis_fifo_96_aresetn;
            assign tlast[96] = s_axis_fifo_96_tlast;
            assign tvalid[96] = s_axis_fifo_96_tvalid;
            assign read[96] = ap_fifo_iarg_96_read;
            assign tkeep[96][S_AXIS_FIFO_96_DMWIDTH/8-1:0] = s_axis_fifo_96_tkeep;
            assign tstrb[96][S_AXIS_FIFO_96_DMWIDTH/8-1:0] = s_axis_fifo_96_tstrb;
            assign tdata[96][S_AXIS_FIFO_96_DMWIDTH-1:0] = s_axis_fifo_96_tdata;
            assign s_axis_fifo_96_tready = tready[96];
            assign ap_fifo_iarg_96_empty_n = empty[96];
            assign ap_fifo_iarg_96_dout = dout[96][S_AXIS_FIFO_96_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 97) begin
            assign axis_clk[97] = s_axis_fifo_97_aclk;
            assign axis_rst[97] = s_axis_fifo_97_aresetn;
            assign tlast[97] = s_axis_fifo_97_tlast;
            assign tvalid[97] = s_axis_fifo_97_tvalid;
            assign read[97] = ap_fifo_iarg_97_read;
            assign tkeep[97][S_AXIS_FIFO_97_DMWIDTH/8-1:0] = s_axis_fifo_97_tkeep;
            assign tstrb[97][S_AXIS_FIFO_97_DMWIDTH/8-1:0] = s_axis_fifo_97_tstrb;
            assign tdata[97][S_AXIS_FIFO_97_DMWIDTH-1:0] = s_axis_fifo_97_tdata;
            assign s_axis_fifo_97_tready = tready[97];
            assign ap_fifo_iarg_97_empty_n = empty[97];
            assign ap_fifo_iarg_97_dout = dout[97][S_AXIS_FIFO_97_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 98) begin
            assign axis_clk[98] = s_axis_fifo_98_aclk;
            assign axis_rst[98] = s_axis_fifo_98_aresetn;
            assign tlast[98] = s_axis_fifo_98_tlast;
            assign tvalid[98] = s_axis_fifo_98_tvalid;
            assign read[98] = ap_fifo_iarg_98_read;
            assign tkeep[98][S_AXIS_FIFO_98_DMWIDTH/8-1:0] = s_axis_fifo_98_tkeep;
            assign tstrb[98][S_AXIS_FIFO_98_DMWIDTH/8-1:0] = s_axis_fifo_98_tstrb;
            assign tdata[98][S_AXIS_FIFO_98_DMWIDTH-1:0] = s_axis_fifo_98_tdata;
            assign s_axis_fifo_98_tready = tready[98];
            assign ap_fifo_iarg_98_empty_n = empty[98];
            assign ap_fifo_iarg_98_dout = dout[98][S_AXIS_FIFO_98_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 99) begin
            assign axis_clk[99] = s_axis_fifo_99_aclk;
            assign axis_rst[99] = s_axis_fifo_99_aresetn;
            assign tlast[99] = s_axis_fifo_99_tlast;
            assign tvalid[99] = s_axis_fifo_99_tvalid;
            assign read[99] = ap_fifo_iarg_99_read;
            assign tkeep[99][S_AXIS_FIFO_99_DMWIDTH/8-1:0] = s_axis_fifo_99_tkeep;
            assign tstrb[99][S_AXIS_FIFO_99_DMWIDTH/8-1:0] = s_axis_fifo_99_tstrb;
            assign tdata[99][S_AXIS_FIFO_99_DMWIDTH-1:0] = s_axis_fifo_99_tdata;
            assign s_axis_fifo_99_tready = tready[99];
            assign ap_fifo_iarg_99_empty_n = empty[99];
            assign ap_fifo_iarg_99_dout = dout[99][S_AXIS_FIFO_99_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 100) begin
            assign axis_clk[100] = s_axis_fifo_100_aclk;
            assign axis_rst[100] = s_axis_fifo_100_aresetn;
            assign tlast[100] = s_axis_fifo_100_tlast;
            assign tvalid[100] = s_axis_fifo_100_tvalid;
            assign read[100] = ap_fifo_iarg_100_read;
            assign tkeep[100][S_AXIS_FIFO_100_DMWIDTH/8-1:0] = s_axis_fifo_100_tkeep;
            assign tstrb[100][S_AXIS_FIFO_100_DMWIDTH/8-1:0] = s_axis_fifo_100_tstrb;
            assign tdata[100][S_AXIS_FIFO_100_DMWIDTH-1:0] = s_axis_fifo_100_tdata;
            assign s_axis_fifo_100_tready = tready[100];
            assign ap_fifo_iarg_100_empty_n = empty[100];
            assign ap_fifo_iarg_100_dout = dout[100][S_AXIS_FIFO_100_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 101) begin
            assign axis_clk[101] = s_axis_fifo_101_aclk;
            assign axis_rst[101] = s_axis_fifo_101_aresetn;
            assign tlast[101] = s_axis_fifo_101_tlast;
            assign tvalid[101] = s_axis_fifo_101_tvalid;
            assign read[101] = ap_fifo_iarg_101_read;
            assign tkeep[101][S_AXIS_FIFO_101_DMWIDTH/8-1:0] = s_axis_fifo_101_tkeep;
            assign tstrb[101][S_AXIS_FIFO_101_DMWIDTH/8-1:0] = s_axis_fifo_101_tstrb;
            assign tdata[101][S_AXIS_FIFO_101_DMWIDTH-1:0] = s_axis_fifo_101_tdata;
            assign s_axis_fifo_101_tready = tready[101];
            assign ap_fifo_iarg_101_empty_n = empty[101];
            assign ap_fifo_iarg_101_dout = dout[101][S_AXIS_FIFO_101_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 102) begin
            assign axis_clk[102] = s_axis_fifo_102_aclk;
            assign axis_rst[102] = s_axis_fifo_102_aresetn;
            assign tlast[102] = s_axis_fifo_102_tlast;
            assign tvalid[102] = s_axis_fifo_102_tvalid;
            assign read[102] = ap_fifo_iarg_102_read;
            assign tkeep[102][S_AXIS_FIFO_102_DMWIDTH/8-1:0] = s_axis_fifo_102_tkeep;
            assign tstrb[102][S_AXIS_FIFO_102_DMWIDTH/8-1:0] = s_axis_fifo_102_tstrb;
            assign tdata[102][S_AXIS_FIFO_102_DMWIDTH-1:0] = s_axis_fifo_102_tdata;
            assign s_axis_fifo_102_tready = tready[102];
            assign ap_fifo_iarg_102_empty_n = empty[102];
            assign ap_fifo_iarg_102_dout = dout[102][S_AXIS_FIFO_102_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 103) begin
            assign axis_clk[103] = s_axis_fifo_103_aclk;
            assign axis_rst[103] = s_axis_fifo_103_aresetn;
            assign tlast[103] = s_axis_fifo_103_tlast;
            assign tvalid[103] = s_axis_fifo_103_tvalid;
            assign read[103] = ap_fifo_iarg_103_read;
            assign tkeep[103][S_AXIS_FIFO_103_DMWIDTH/8-1:0] = s_axis_fifo_103_tkeep;
            assign tstrb[103][S_AXIS_FIFO_103_DMWIDTH/8-1:0] = s_axis_fifo_103_tstrb;
            assign tdata[103][S_AXIS_FIFO_103_DMWIDTH-1:0] = s_axis_fifo_103_tdata;
            assign s_axis_fifo_103_tready = tready[103];
            assign ap_fifo_iarg_103_empty_n = empty[103];
            assign ap_fifo_iarg_103_dout = dout[103][S_AXIS_FIFO_103_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 104) begin
            assign axis_clk[104] = s_axis_fifo_104_aclk;
            assign axis_rst[104] = s_axis_fifo_104_aresetn;
            assign tlast[104] = s_axis_fifo_104_tlast;
            assign tvalid[104] = s_axis_fifo_104_tvalid;
            assign read[104] = ap_fifo_iarg_104_read;
            assign tkeep[104][S_AXIS_FIFO_104_DMWIDTH/8-1:0] = s_axis_fifo_104_tkeep;
            assign tstrb[104][S_AXIS_FIFO_104_DMWIDTH/8-1:0] = s_axis_fifo_104_tstrb;
            assign tdata[104][S_AXIS_FIFO_104_DMWIDTH-1:0] = s_axis_fifo_104_tdata;
            assign s_axis_fifo_104_tready = tready[104];
            assign ap_fifo_iarg_104_empty_n = empty[104];
            assign ap_fifo_iarg_104_dout = dout[104][S_AXIS_FIFO_104_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 105) begin
            assign axis_clk[105] = s_axis_fifo_105_aclk;
            assign axis_rst[105] = s_axis_fifo_105_aresetn;
            assign tlast[105] = s_axis_fifo_105_tlast;
            assign tvalid[105] = s_axis_fifo_105_tvalid;
            assign read[105] = ap_fifo_iarg_105_read;
            assign tkeep[105][S_AXIS_FIFO_105_DMWIDTH/8-1:0] = s_axis_fifo_105_tkeep;
            assign tstrb[105][S_AXIS_FIFO_105_DMWIDTH/8-1:0] = s_axis_fifo_105_tstrb;
            assign tdata[105][S_AXIS_FIFO_105_DMWIDTH-1:0] = s_axis_fifo_105_tdata;
            assign s_axis_fifo_105_tready = tready[105];
            assign ap_fifo_iarg_105_empty_n = empty[105];
            assign ap_fifo_iarg_105_dout = dout[105][S_AXIS_FIFO_105_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 106) begin
            assign axis_clk[106] = s_axis_fifo_106_aclk;
            assign axis_rst[106] = s_axis_fifo_106_aresetn;
            assign tlast[106] = s_axis_fifo_106_tlast;
            assign tvalid[106] = s_axis_fifo_106_tvalid;
            assign read[106] = ap_fifo_iarg_106_read;
            assign tkeep[106][S_AXIS_FIFO_106_DMWIDTH/8-1:0] = s_axis_fifo_106_tkeep;
            assign tstrb[106][S_AXIS_FIFO_106_DMWIDTH/8-1:0] = s_axis_fifo_106_tstrb;
            assign tdata[106][S_AXIS_FIFO_106_DMWIDTH-1:0] = s_axis_fifo_106_tdata;
            assign s_axis_fifo_106_tready = tready[106];
            assign ap_fifo_iarg_106_empty_n = empty[106];
            assign ap_fifo_iarg_106_dout = dout[106][S_AXIS_FIFO_106_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 107) begin
            assign axis_clk[107] = s_axis_fifo_107_aclk;
            assign axis_rst[107] = s_axis_fifo_107_aresetn;
            assign tlast[107] = s_axis_fifo_107_tlast;
            assign tvalid[107] = s_axis_fifo_107_tvalid;
            assign read[107] = ap_fifo_iarg_107_read;
            assign tkeep[107][S_AXIS_FIFO_107_DMWIDTH/8-1:0] = s_axis_fifo_107_tkeep;
            assign tstrb[107][S_AXIS_FIFO_107_DMWIDTH/8-1:0] = s_axis_fifo_107_tstrb;
            assign tdata[107][S_AXIS_FIFO_107_DMWIDTH-1:0] = s_axis_fifo_107_tdata;
            assign s_axis_fifo_107_tready = tready[107];
            assign ap_fifo_iarg_107_empty_n = empty[107];
            assign ap_fifo_iarg_107_dout = dout[107][S_AXIS_FIFO_107_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 108) begin
            assign axis_clk[108] = s_axis_fifo_108_aclk;
            assign axis_rst[108] = s_axis_fifo_108_aresetn;
            assign tlast[108] = s_axis_fifo_108_tlast;
            assign tvalid[108] = s_axis_fifo_108_tvalid;
            assign read[108] = ap_fifo_iarg_108_read;
            assign tkeep[108][S_AXIS_FIFO_108_DMWIDTH/8-1:0] = s_axis_fifo_108_tkeep;
            assign tstrb[108][S_AXIS_FIFO_108_DMWIDTH/8-1:0] = s_axis_fifo_108_tstrb;
            assign tdata[108][S_AXIS_FIFO_108_DMWIDTH-1:0] = s_axis_fifo_108_tdata;
            assign s_axis_fifo_108_tready = tready[108];
            assign ap_fifo_iarg_108_empty_n = empty[108];
            assign ap_fifo_iarg_108_dout = dout[108][S_AXIS_FIFO_108_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 109) begin
            assign axis_clk[109] = s_axis_fifo_109_aclk;
            assign axis_rst[109] = s_axis_fifo_109_aresetn;
            assign tlast[109] = s_axis_fifo_109_tlast;
            assign tvalid[109] = s_axis_fifo_109_tvalid;
            assign read[109] = ap_fifo_iarg_109_read;
            assign tkeep[109][S_AXIS_FIFO_109_DMWIDTH/8-1:0] = s_axis_fifo_109_tkeep;
            assign tstrb[109][S_AXIS_FIFO_109_DMWIDTH/8-1:0] = s_axis_fifo_109_tstrb;
            assign tdata[109][S_AXIS_FIFO_109_DMWIDTH-1:0] = s_axis_fifo_109_tdata;
            assign s_axis_fifo_109_tready = tready[109];
            assign ap_fifo_iarg_109_empty_n = empty[109];
            assign ap_fifo_iarg_109_dout = dout[109][S_AXIS_FIFO_109_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 110) begin
            assign axis_clk[110] = s_axis_fifo_110_aclk;
            assign axis_rst[110] = s_axis_fifo_110_aresetn;
            assign tlast[110] = s_axis_fifo_110_tlast;
            assign tvalid[110] = s_axis_fifo_110_tvalid;
            assign read[110] = ap_fifo_iarg_110_read;
            assign tkeep[110][S_AXIS_FIFO_110_DMWIDTH/8-1:0] = s_axis_fifo_110_tkeep;
            assign tstrb[110][S_AXIS_FIFO_110_DMWIDTH/8-1:0] = s_axis_fifo_110_tstrb;
            assign tdata[110][S_AXIS_FIFO_110_DMWIDTH-1:0] = s_axis_fifo_110_tdata;
            assign s_axis_fifo_110_tready = tready[110];
            assign ap_fifo_iarg_110_empty_n = empty[110];
            assign ap_fifo_iarg_110_dout = dout[110][S_AXIS_FIFO_110_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 111) begin
            assign axis_clk[111] = s_axis_fifo_111_aclk;
            assign axis_rst[111] = s_axis_fifo_111_aresetn;
            assign tlast[111] = s_axis_fifo_111_tlast;
            assign tvalid[111] = s_axis_fifo_111_tvalid;
            assign read[111] = ap_fifo_iarg_111_read;
            assign tkeep[111][S_AXIS_FIFO_111_DMWIDTH/8-1:0] = s_axis_fifo_111_tkeep;
            assign tstrb[111][S_AXIS_FIFO_111_DMWIDTH/8-1:0] = s_axis_fifo_111_tstrb;
            assign tdata[111][S_AXIS_FIFO_111_DMWIDTH-1:0] = s_axis_fifo_111_tdata;
            assign s_axis_fifo_111_tready = tready[111];
            assign ap_fifo_iarg_111_empty_n = empty[111];
            assign ap_fifo_iarg_111_dout = dout[111][S_AXIS_FIFO_111_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 112) begin
            assign axis_clk[112] = s_axis_fifo_112_aclk;
            assign axis_rst[112] = s_axis_fifo_112_aresetn;
            assign tlast[112] = s_axis_fifo_112_tlast;
            assign tvalid[112] = s_axis_fifo_112_tvalid;
            assign read[112] = ap_fifo_iarg_112_read;
            assign tkeep[112][S_AXIS_FIFO_112_DMWIDTH/8-1:0] = s_axis_fifo_112_tkeep;
            assign tstrb[112][S_AXIS_FIFO_112_DMWIDTH/8-1:0] = s_axis_fifo_112_tstrb;
            assign tdata[112][S_AXIS_FIFO_112_DMWIDTH-1:0] = s_axis_fifo_112_tdata;
            assign s_axis_fifo_112_tready = tready[112];
            assign ap_fifo_iarg_112_empty_n = empty[112];
            assign ap_fifo_iarg_112_dout = dout[112][S_AXIS_FIFO_112_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 113) begin
            assign axis_clk[113] = s_axis_fifo_113_aclk;
            assign axis_rst[113] = s_axis_fifo_113_aresetn;
            assign tlast[113] = s_axis_fifo_113_tlast;
            assign tvalid[113] = s_axis_fifo_113_tvalid;
            assign read[113] = ap_fifo_iarg_113_read;
            assign tkeep[113][S_AXIS_FIFO_113_DMWIDTH/8-1:0] = s_axis_fifo_113_tkeep;
            assign tstrb[113][S_AXIS_FIFO_113_DMWIDTH/8-1:0] = s_axis_fifo_113_tstrb;
            assign tdata[113][S_AXIS_FIFO_113_DMWIDTH-1:0] = s_axis_fifo_113_tdata;
            assign s_axis_fifo_113_tready = tready[113];
            assign ap_fifo_iarg_113_empty_n = empty[113];
            assign ap_fifo_iarg_113_dout = dout[113][S_AXIS_FIFO_113_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 114) begin
            assign axis_clk[114] = s_axis_fifo_114_aclk;
            assign axis_rst[114] = s_axis_fifo_114_aresetn;
            assign tlast[114] = s_axis_fifo_114_tlast;
            assign tvalid[114] = s_axis_fifo_114_tvalid;
            assign read[114] = ap_fifo_iarg_114_read;
            assign tkeep[114][S_AXIS_FIFO_114_DMWIDTH/8-1:0] = s_axis_fifo_114_tkeep;
            assign tstrb[114][S_AXIS_FIFO_114_DMWIDTH/8-1:0] = s_axis_fifo_114_tstrb;
            assign tdata[114][S_AXIS_FIFO_114_DMWIDTH-1:0] = s_axis_fifo_114_tdata;
            assign s_axis_fifo_114_tready = tready[114];
            assign ap_fifo_iarg_114_empty_n = empty[114];
            assign ap_fifo_iarg_114_dout = dout[114][S_AXIS_FIFO_114_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 115) begin
            assign axis_clk[115] = s_axis_fifo_115_aclk;
            assign axis_rst[115] = s_axis_fifo_115_aresetn;
            assign tlast[115] = s_axis_fifo_115_tlast;
            assign tvalid[115] = s_axis_fifo_115_tvalid;
            assign read[115] = ap_fifo_iarg_115_read;
            assign tkeep[115][S_AXIS_FIFO_115_DMWIDTH/8-1:0] = s_axis_fifo_115_tkeep;
            assign tstrb[115][S_AXIS_FIFO_115_DMWIDTH/8-1:0] = s_axis_fifo_115_tstrb;
            assign tdata[115][S_AXIS_FIFO_115_DMWIDTH-1:0] = s_axis_fifo_115_tdata;
            assign s_axis_fifo_115_tready = tready[115];
            assign ap_fifo_iarg_115_empty_n = empty[115];
            assign ap_fifo_iarg_115_dout = dout[115][S_AXIS_FIFO_115_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 116) begin
            assign axis_clk[116] = s_axis_fifo_116_aclk;
            assign axis_rst[116] = s_axis_fifo_116_aresetn;
            assign tlast[116] = s_axis_fifo_116_tlast;
            assign tvalid[116] = s_axis_fifo_116_tvalid;
            assign read[116] = ap_fifo_iarg_116_read;
            assign tkeep[116][S_AXIS_FIFO_116_DMWIDTH/8-1:0] = s_axis_fifo_116_tkeep;
            assign tstrb[116][S_AXIS_FIFO_116_DMWIDTH/8-1:0] = s_axis_fifo_116_tstrb;
            assign tdata[116][S_AXIS_FIFO_116_DMWIDTH-1:0] = s_axis_fifo_116_tdata;
            assign s_axis_fifo_116_tready = tready[116];
            assign ap_fifo_iarg_116_empty_n = empty[116];
            assign ap_fifo_iarg_116_dout = dout[116][S_AXIS_FIFO_116_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 117) begin
            assign axis_clk[117] = s_axis_fifo_117_aclk;
            assign axis_rst[117] = s_axis_fifo_117_aresetn;
            assign tlast[117] = s_axis_fifo_117_tlast;
            assign tvalid[117] = s_axis_fifo_117_tvalid;
            assign read[117] = ap_fifo_iarg_117_read;
            assign tkeep[117][S_AXIS_FIFO_117_DMWIDTH/8-1:0] = s_axis_fifo_117_tkeep;
            assign tstrb[117][S_AXIS_FIFO_117_DMWIDTH/8-1:0] = s_axis_fifo_117_tstrb;
            assign tdata[117][S_AXIS_FIFO_117_DMWIDTH-1:0] = s_axis_fifo_117_tdata;
            assign s_axis_fifo_117_tready = tready[117];
            assign ap_fifo_iarg_117_empty_n = empty[117];
            assign ap_fifo_iarg_117_dout = dout[117][S_AXIS_FIFO_117_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 118) begin
            assign axis_clk[118] = s_axis_fifo_118_aclk;
            assign axis_rst[118] = s_axis_fifo_118_aresetn;
            assign tlast[118] = s_axis_fifo_118_tlast;
            assign tvalid[118] = s_axis_fifo_118_tvalid;
            assign read[118] = ap_fifo_iarg_118_read;
            assign tkeep[118][S_AXIS_FIFO_118_DMWIDTH/8-1:0] = s_axis_fifo_118_tkeep;
            assign tstrb[118][S_AXIS_FIFO_118_DMWIDTH/8-1:0] = s_axis_fifo_118_tstrb;
            assign tdata[118][S_AXIS_FIFO_118_DMWIDTH-1:0] = s_axis_fifo_118_tdata;
            assign s_axis_fifo_118_tready = tready[118];
            assign ap_fifo_iarg_118_empty_n = empty[118];
            assign ap_fifo_iarg_118_dout = dout[118][S_AXIS_FIFO_118_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 119) begin
            assign axis_clk[119] = s_axis_fifo_119_aclk;
            assign axis_rst[119] = s_axis_fifo_119_aresetn;
            assign tlast[119] = s_axis_fifo_119_tlast;
            assign tvalid[119] = s_axis_fifo_119_tvalid;
            assign read[119] = ap_fifo_iarg_119_read;
            assign tkeep[119][S_AXIS_FIFO_119_DMWIDTH/8-1:0] = s_axis_fifo_119_tkeep;
            assign tstrb[119][S_AXIS_FIFO_119_DMWIDTH/8-1:0] = s_axis_fifo_119_tstrb;
            assign tdata[119][S_AXIS_FIFO_119_DMWIDTH-1:0] = s_axis_fifo_119_tdata;
            assign s_axis_fifo_119_tready = tready[119];
            assign ap_fifo_iarg_119_empty_n = empty[119];
            assign ap_fifo_iarg_119_dout = dout[119][S_AXIS_FIFO_119_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 120) begin
            assign axis_clk[120] = s_axis_fifo_120_aclk;
            assign axis_rst[120] = s_axis_fifo_120_aresetn;
            assign tlast[120] = s_axis_fifo_120_tlast;
            assign tvalid[120] = s_axis_fifo_120_tvalid;
            assign read[120] = ap_fifo_iarg_120_read;
            assign tkeep[120][S_AXIS_FIFO_120_DMWIDTH/8-1:0] = s_axis_fifo_120_tkeep;
            assign tstrb[120][S_AXIS_FIFO_120_DMWIDTH/8-1:0] = s_axis_fifo_120_tstrb;
            assign tdata[120][S_AXIS_FIFO_120_DMWIDTH-1:0] = s_axis_fifo_120_tdata;
            assign s_axis_fifo_120_tready = tready[120];
            assign ap_fifo_iarg_120_empty_n = empty[120];
            assign ap_fifo_iarg_120_dout = dout[120][S_AXIS_FIFO_120_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 121) begin
            assign axis_clk[121] = s_axis_fifo_121_aclk;
            assign axis_rst[121] = s_axis_fifo_121_aresetn;
            assign tlast[121] = s_axis_fifo_121_tlast;
            assign tvalid[121] = s_axis_fifo_121_tvalid;
            assign read[121] = ap_fifo_iarg_121_read;
            assign tkeep[121][S_AXIS_FIFO_121_DMWIDTH/8-1:0] = s_axis_fifo_121_tkeep;
            assign tstrb[121][S_AXIS_FIFO_121_DMWIDTH/8-1:0] = s_axis_fifo_121_tstrb;
            assign tdata[121][S_AXIS_FIFO_121_DMWIDTH-1:0] = s_axis_fifo_121_tdata;
            assign s_axis_fifo_121_tready = tready[121];
            assign ap_fifo_iarg_121_empty_n = empty[121];
            assign ap_fifo_iarg_121_dout = dout[121][S_AXIS_FIFO_121_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 122) begin
            assign axis_clk[122] = s_axis_fifo_122_aclk;
            assign axis_rst[122] = s_axis_fifo_122_aresetn;
            assign tlast[122] = s_axis_fifo_122_tlast;
            assign tvalid[122] = s_axis_fifo_122_tvalid;
            assign read[122] = ap_fifo_iarg_122_read;
            assign tkeep[122][S_AXIS_FIFO_122_DMWIDTH/8-1:0] = s_axis_fifo_122_tkeep;
            assign tstrb[122][S_AXIS_FIFO_122_DMWIDTH/8-1:0] = s_axis_fifo_122_tstrb;
            assign tdata[122][S_AXIS_FIFO_122_DMWIDTH-1:0] = s_axis_fifo_122_tdata;
            assign s_axis_fifo_122_tready = tready[122];
            assign ap_fifo_iarg_122_empty_n = empty[122];
            assign ap_fifo_iarg_122_dout = dout[122][S_AXIS_FIFO_122_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 123) begin
            assign axis_clk[123] = s_axis_fifo_123_aclk;
            assign axis_rst[123] = s_axis_fifo_123_aresetn;
            assign tlast[123] = s_axis_fifo_123_tlast;
            assign tvalid[123] = s_axis_fifo_123_tvalid;
            assign read[123] = ap_fifo_iarg_123_read;
            assign tkeep[123][S_AXIS_FIFO_123_DMWIDTH/8-1:0] = s_axis_fifo_123_tkeep;
            assign tstrb[123][S_AXIS_FIFO_123_DMWIDTH/8-1:0] = s_axis_fifo_123_tstrb;
            assign tdata[123][S_AXIS_FIFO_123_DMWIDTH-1:0] = s_axis_fifo_123_tdata;
            assign s_axis_fifo_123_tready = tready[123];
            assign ap_fifo_iarg_123_empty_n = empty[123];
            assign ap_fifo_iarg_123_dout = dout[123][S_AXIS_FIFO_123_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 124) begin
            assign axis_clk[124] = s_axis_fifo_124_aclk;
            assign axis_rst[124] = s_axis_fifo_124_aresetn;
            assign tlast[124] = s_axis_fifo_124_tlast;
            assign tvalid[124] = s_axis_fifo_124_tvalid;
            assign read[124] = ap_fifo_iarg_124_read;
            assign tkeep[124][S_AXIS_FIFO_124_DMWIDTH/8-1:0] = s_axis_fifo_124_tkeep;
            assign tstrb[124][S_AXIS_FIFO_124_DMWIDTH/8-1:0] = s_axis_fifo_124_tstrb;
            assign tdata[124][S_AXIS_FIFO_124_DMWIDTH-1:0] = s_axis_fifo_124_tdata;
            assign s_axis_fifo_124_tready = tready[124];
            assign ap_fifo_iarg_124_empty_n = empty[124];
            assign ap_fifo_iarg_124_dout = dout[124][S_AXIS_FIFO_124_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 125) begin
            assign axis_clk[125] = s_axis_fifo_125_aclk;
            assign axis_rst[125] = s_axis_fifo_125_aresetn;
            assign tlast[125] = s_axis_fifo_125_tlast;
            assign tvalid[125] = s_axis_fifo_125_tvalid;
            assign read[125] = ap_fifo_iarg_125_read;
            assign tkeep[125][S_AXIS_FIFO_125_DMWIDTH/8-1:0] = s_axis_fifo_125_tkeep;
            assign tstrb[125][S_AXIS_FIFO_125_DMWIDTH/8-1:0] = s_axis_fifo_125_tstrb;
            assign tdata[125][S_AXIS_FIFO_125_DMWIDTH-1:0] = s_axis_fifo_125_tdata;
            assign s_axis_fifo_125_tready = tready[125];
            assign ap_fifo_iarg_125_empty_n = empty[125];
            assign ap_fifo_iarg_125_dout = dout[125][S_AXIS_FIFO_125_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 126) begin
            assign axis_clk[126] = s_axis_fifo_126_aclk;
            assign axis_rst[126] = s_axis_fifo_126_aresetn;
            assign tlast[126] = s_axis_fifo_126_tlast;
            assign tvalid[126] = s_axis_fifo_126_tvalid;
            assign read[126] = ap_fifo_iarg_126_read;
            assign tkeep[126][S_AXIS_FIFO_126_DMWIDTH/8-1:0] = s_axis_fifo_126_tkeep;
            assign tstrb[126][S_AXIS_FIFO_126_DMWIDTH/8-1:0] = s_axis_fifo_126_tstrb;
            assign tdata[126][S_AXIS_FIFO_126_DMWIDTH-1:0] = s_axis_fifo_126_tdata;
            assign s_axis_fifo_126_tready = tready[126];
            assign ap_fifo_iarg_126_empty_n = empty[126];
            assign ap_fifo_iarg_126_dout = dout[126][S_AXIS_FIFO_126_BYTE_WIDTH-1:0];
        end
        if(C_NUM_INPUT_FIFOs > 127) begin
            assign axis_clk[127] = s_axis_fifo_127_aclk;
            assign axis_rst[127] = s_axis_fifo_127_aresetn;
            assign tlast[127] = s_axis_fifo_127_tlast;
            assign tvalid[127] = s_axis_fifo_127_tvalid;
            assign read[127] = ap_fifo_iarg_127_read;
            assign tkeep[127][S_AXIS_FIFO_127_DMWIDTH/8-1:0] = s_axis_fifo_127_tkeep;
            assign tstrb[127][S_AXIS_FIFO_127_DMWIDTH/8-1:0] = s_axis_fifo_127_tstrb;
            assign tdata[127][S_AXIS_FIFO_127_DMWIDTH-1:0] = s_axis_fifo_127_tdata;
            assign s_axis_fifo_127_tready = tready[127];
            assign ap_fifo_iarg_127_empty_n = empty[127];
            assign ap_fifo_iarg_127_dout = dout[127][S_AXIS_FIFO_127_BYTE_WIDTH-1:0];
        end
    endgenerate
    
    //instantiate the axis2fifo modules
    genvar idx;
    generate
        for(idx=0; idx<C_NUM_INPUT_FIFOs; idx=idx+1) begin: IN_FIFO_GEN
            //check if data width converter is needed
            if(C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx] != C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]) begin
                 axis_dwidth_converter_v1_1_9_axis_dwidth_converter #(
                    .C_S_AXIS_TDATA_WIDTH(C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_M_AXIS_TDATA_WIDTH(C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_AXIS_TID_WIDTH(1),
                    .C_AXIS_TDEST_WIDTH(1),
                    .C_S_AXIS_TUSER_WIDTH(1),
                    .C_M_AXIS_TUSER_WIDTH(1),
                    .C_AXIS_SIGNAL_SET(32'h1F)  //Enabled: TLAST, TKEEP, TSTRB, TDATA, TREADY
                ) data_width_conv_i (
                    .aclk(axis_clk[idx]),
                    .aresetn(axis_rst[idx]),
                    .aclken(1'b1),
                    .s_axis_tvalid(tvalid[idx]),
                    .s_axis_tready(tready[idx]),
                    .s_axis_tdata(tdata[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .s_axis_tstrb(tstrb[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tkeep(tkeep[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tlast(tlast[idx]),
//                    .s_axis_tid(),
//                    .s_axis_tdest(),
//                    .s_axis_tuser(),
                    .m_axis_tvalid(dwconv_tvalid[idx]),
                    .m_axis_tready(dwconv_tready[idx]),
                    .m_axis_tdata(dwconv_tdata[idx][C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
//                    .m_axis_tstrb(),
//                    .m_axis_tkeep(),
                    .m_axis_tlast(dwconv_tlast[idx])
//                    .m_axis_tid(),
//                    .m_axis_tdest(),
//                    .m_axis_tuser()
                );
            end
            else begin
                //if no data width conversion, wire the input signals straight through
                assign dwconv_tlast[idx] = tlast[idx];
                assign dwconv_tvalid[idx] = tvalid[idx];
                assign tready[idx] = dwconv_tready[idx];   //output
                assign dwconv_tdata[idx][C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = tdata[idx][C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            end
            
            if(C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx] != C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]) begin
                //use truncator
                axisTrunc #(
                    .IN_WIDTH(C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .OUT_WIDTH(C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx])
                ) axis_trunc_i (
                    .IN_TLAST(dwconv_tlast[idx]),
                    .IN_TVALID(dwconv_tvalid[idx]),
                    .IN_TDATA(dwconv_tdata[idx][C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .IN_TREADY(dwconv_tready[idx]),
                    .OUT_TLAST(trunc_tlast[idx]),
                    .OUT_TVALID(trunc_tvalid[idx]),
                    .OUT_TDATA(trunc_tdata[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .OUT_TREADY(trunc_tready[idx])
                );
            end
            else begin
                //if not, wire the input signals straight through
                assign trunc_tlast[idx] = dwconv_tlast[idx];
                assign trunc_tvalid[idx] = dwconv_tvalid[idx];
                assign dwconv_tready[idx] = trunc_tready[idx];   //output
                assign trunc_tdata[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0] = dwconv_tdata[idx][C_INFIFO_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            end
            
            if(C_DEPTH_BIT_ARRAY[32*(idx+1)-1:32*idx] > 0) begin
                //use fifo
                axis_fifo #(
                    .C_DATA_WIDTH(C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_DATA_DEPTH(C_DEPTH_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_IS_ASYNC(C_IS_ASYNC_BIT_ARRAY[32*(idx+1)-1:32*idx])
                ) axis_fifo_i (
                    .aresetn(axis_rst[idx]),
                    .inclk(axis_clk[idx]),
                    .in_tdata(trunc_tdata[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .in_tlast(trunc_tlast[idx]),  
                    .in_tvalid(trunc_tvalid[idx]),
                    .in_tready(trunc_tready[idx]),
                    .outclk(acc_clk), 
                    .out_tdata(buf_tdata[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .out_tready(buf_tready[idx]),
                    .out_tvalid(buf_tvalid[idx]),
                    .out_tlast(buf_tlast[idx])
                );
            end
            else begin
                //if not, wire the input signals straight through
                assign buf_tlast[idx] = trunc_tlast[idx];
                assign buf_tvalid[idx] = trunc_tvalid[idx];
                assign trunc_tready[idx] = buf_tready[idx];   //output
                assign buf_tdata[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0] = trunc_tdata[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            end
            
            axis2fifo #( 
                .DATA_WIDTH(C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx])
            ) axis2fifo_i (
                .ACC_CLK(acc_clk),
                .ARESETN(acc_aresetn),
                .CTRL_ALLOW(in_fifo_allow),
                .CTRL_READY(in_fifo_ready[idx]),
                .CTRL_FINISHED(in_fifo_finished[idx]),
                .AXIS_TLAST(buf_tlast[idx]),
                .AXIS_TVALID(buf_tvalid[idx]),
                .AXIS_TDATA(buf_tdata[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .AXIS_TREADY(buf_tready[idx]),
                .FIFO_EMPTY(empty[idx]),
                .FIFO_DOUT(dout[idx][C_INFIFO_REAL_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .FIFO_READ(read[idx])
            );
        end
    endgenerate
endmodule
