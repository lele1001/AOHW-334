// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689
`timescale 1ns / 1ps

module in_axis_args #(
    parameter C_NUM_INPUT_AXISs = 0,
    parameter [31:0] S_AXIS_IARG_0_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_1_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_2_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_3_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_4_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_5_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_6_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_7_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_8_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_9_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_10_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_11_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_12_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_13_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_14_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_15_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_16_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_17_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_18_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_19_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_20_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_21_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_22_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_23_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_24_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_25_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_26_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_27_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_28_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_29_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_30_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_31_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_32_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_33_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_34_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_35_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_36_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_37_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_38_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_39_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_40_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_41_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_42_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_43_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_44_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_45_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_46_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_47_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_48_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_49_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_50_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_51_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_52_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_53_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_54_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_55_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_56_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_57_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_58_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_59_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_60_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_61_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_62_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_63_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_64_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_65_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_66_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_67_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_68_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_69_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_70_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_71_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_72_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_73_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_74_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_75_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_76_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_77_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_78_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_79_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_80_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_81_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_82_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_83_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_84_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_85_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_86_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_87_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_88_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_89_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_90_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_91_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_92_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_93_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_94_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_95_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_96_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_97_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_98_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_99_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_100_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_101_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_102_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_103_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_104_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_105_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_106_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_107_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_108_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_109_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_110_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_111_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_112_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_113_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_114_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_115_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_116_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_117_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_118_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_119_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_120_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_121_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_122_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_123_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_124_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_125_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_126_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_127_WIDTH = 8,     //width of input axis interface on the accelerator
    parameter [31:0] S_AXIS_IARG_0_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_1_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_2_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_3_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_4_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_5_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_6_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_7_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_8_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_9_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_10_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_11_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_12_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_13_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_14_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_15_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_16_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_17_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_18_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_19_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_20_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_21_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_22_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_23_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_24_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_25_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_26_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_27_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_28_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_29_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_30_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_31_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_32_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_33_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_34_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_35_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_36_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_37_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_38_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_39_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_40_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_41_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_42_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_43_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_44_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_45_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_46_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_47_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_48_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_49_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_50_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_51_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_52_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_53_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_54_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_55_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_56_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_57_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_58_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_59_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_60_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_61_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_62_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_63_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_64_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_65_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_66_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_67_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_68_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_69_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_70_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_71_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_72_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_73_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_74_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_75_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_76_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_77_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_78_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_79_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_80_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_81_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_82_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_83_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_84_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_85_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_86_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_87_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_88_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_89_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_90_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_91_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_92_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_93_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_94_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_95_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_96_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_97_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_98_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_99_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_100_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_101_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_102_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_103_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_104_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_105_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_106_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_107_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_108_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_109_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_110_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_111_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_112_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_113_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_114_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_115_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_116_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_117_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_118_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_119_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_120_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_121_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_122_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_123_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_124_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_125_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_126_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_127_DEPTH = 16,      //depth of AXIS in adapter for input axis interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_0_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_1_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_2_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_3_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_4_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_5_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_6_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_7_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_8_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_9_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_10_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_11_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_12_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_13_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_14_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_15_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_16_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_17_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_18_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_19_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_20_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_21_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_22_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_23_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_24_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_25_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_26_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_27_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_28_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_29_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_30_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_31_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_32_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_33_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_34_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_35_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_36_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_37_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_38_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_39_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_40_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_41_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_42_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_43_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_44_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_45_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_46_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_47_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_48_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_49_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_50_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_51_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_52_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_53_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_54_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_55_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_56_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_57_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_58_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_59_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_60_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_61_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_62_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_63_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_64_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_65_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_66_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_67_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_68_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_69_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_70_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_71_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_72_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_73_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_74_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_75_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_76_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_77_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_78_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_79_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_80_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_81_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_82_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_83_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_84_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_85_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_86_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_87_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_88_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_89_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_90_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_91_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_92_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_93_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_94_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_95_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_96_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_97_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_98_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_99_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_100_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_101_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_102_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_103_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_104_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_105_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_106_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_107_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_108_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_109_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_110_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_111_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_112_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_113_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_114_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_115_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_116_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_117_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_118_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_119_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_120_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_121_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_122_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_123_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_124_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_125_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_126_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_127_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input axis interface
    parameter [31:0] S_AXIS_IARG_0_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_1_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_2_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_3_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_4_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_5_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_6_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_7_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_8_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_9_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_10_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_11_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_12_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_13_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_14_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_15_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_16_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_17_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_18_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_19_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_20_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_21_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_22_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_23_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_24_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_25_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_26_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_27_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_28_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_29_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_30_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_31_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_32_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_33_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_34_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_35_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_36_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_37_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_38_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_39_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_40_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_41_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_42_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_43_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_44_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_45_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_46_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_47_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_48_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_49_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_50_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_51_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_52_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_53_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_54_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_55_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_56_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_57_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_58_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_59_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_60_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_61_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_62_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_63_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_64_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_65_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_66_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_67_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_68_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_69_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_70_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_71_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_72_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_73_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_74_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_75_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_76_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_77_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_78_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_79_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_80_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_81_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_82_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_83_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_84_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_85_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_86_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_87_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_88_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_89_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_90_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_91_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_92_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_93_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_94_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_95_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_96_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_97_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_98_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_99_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_100_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_101_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_102_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_103_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_104_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_105_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_106_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_107_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_108_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_109_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_110_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_111_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_112_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_113_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_114_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_115_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_116_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_117_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_118_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_119_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_120_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_121_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_122_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_123_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_124_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_125_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_126_IS_ASYNC = 0,   //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_127_IS_ASYNC = 0   //should fifo buffer be asynchronous (0) or synchronours (1)
 ) (
    input acc_clk,
    input acc_aresetn,
    //control interface
    input in_axis_allow,
    output [C_NUM_INPUT_AXISs-1:0] in_axis_ready,
    output [C_NUM_INPUT_AXISs-1:0] in_axis_finished,
    //input AXI-Stream pass-through interface 0
    input s_axis_iarg_0_aclk,
    input s_axis_iarg_0_aresetn,
    input s_axis_iarg_0_tlast,
    input s_axis_iarg_0_tvalid,
    input [S_AXIS_IARG_0_DMWIDTH/8-1:0] s_axis_iarg_0_tkeep,
    input [S_AXIS_IARG_0_DMWIDTH/8-1:0] s_axis_iarg_0_tstrb,
    input [S_AXIS_IARG_0_DMWIDTH-1:0] s_axis_iarg_0_tdata,
    output s_axis_iarg_0_tready,
    output ap_axis_iarg_0_tlast,
    output ap_axis_iarg_0_tvalid,
    output [S_AXIS_IARG_0_WIDTH/8-1:0] ap_axis_iarg_0_tkeep,
    output [S_AXIS_IARG_0_WIDTH/8-1:0] ap_axis_iarg_0_tstrb,
    output [S_AXIS_IARG_0_WIDTH-1:0] ap_axis_iarg_0_tdata,
    input ap_axis_iarg_0_tready,
    //input AXI-Stream pass-through interface 1
    input s_axis_iarg_1_aclk,
    input s_axis_iarg_1_aresetn,
    input s_axis_iarg_1_tlast,
    input s_axis_iarg_1_tvalid,
    input [S_AXIS_IARG_1_DMWIDTH/8-1:0] s_axis_iarg_1_tkeep,
    input [S_AXIS_IARG_1_DMWIDTH/8-1:0] s_axis_iarg_1_tstrb,
    input [S_AXIS_IARG_1_DMWIDTH-1:0] s_axis_iarg_1_tdata,
    output s_axis_iarg_1_tready,
    output ap_axis_iarg_1_tlast,
    output ap_axis_iarg_1_tvalid,
    output [S_AXIS_IARG_1_WIDTH/8-1:0] ap_axis_iarg_1_tkeep,
    output [S_AXIS_IARG_1_WIDTH/8-1:0] ap_axis_iarg_1_tstrb,
    output [S_AXIS_IARG_1_WIDTH-1:0] ap_axis_iarg_1_tdata,
    input ap_axis_iarg_1_tready,
    //input AXI-Stream pass-through interface 2
    input s_axis_iarg_2_aclk,
    input s_axis_iarg_2_aresetn,
    input s_axis_iarg_2_tlast,
    input s_axis_iarg_2_tvalid,
    input [S_AXIS_IARG_2_DMWIDTH/8-1:0] s_axis_iarg_2_tkeep,
    input [S_AXIS_IARG_2_DMWIDTH/8-1:0] s_axis_iarg_2_tstrb,
    input [S_AXIS_IARG_2_DMWIDTH-1:0] s_axis_iarg_2_tdata,
    output s_axis_iarg_2_tready,
    output ap_axis_iarg_2_tlast,
    output ap_axis_iarg_2_tvalid,
    output [S_AXIS_IARG_2_WIDTH/8-1:0] ap_axis_iarg_2_tkeep,
    output [S_AXIS_IARG_2_WIDTH/8-1:0] ap_axis_iarg_2_tstrb,
    output [S_AXIS_IARG_2_WIDTH-1:0] ap_axis_iarg_2_tdata,
    input ap_axis_iarg_2_tready,
    //input AXI-Stream pass-through interface 3
    input s_axis_iarg_3_aclk,
    input s_axis_iarg_3_aresetn,
    input s_axis_iarg_3_tlast,
    input s_axis_iarg_3_tvalid,
    input [S_AXIS_IARG_3_DMWIDTH/8-1:0] s_axis_iarg_3_tkeep,
    input [S_AXIS_IARG_3_DMWIDTH/8-1:0] s_axis_iarg_3_tstrb,
    input [S_AXIS_IARG_3_DMWIDTH-1:0] s_axis_iarg_3_tdata,
    output s_axis_iarg_3_tready,
    output ap_axis_iarg_3_tlast,
    output ap_axis_iarg_3_tvalid,
    output [S_AXIS_IARG_3_WIDTH/8-1:0] ap_axis_iarg_3_tkeep,
    output [S_AXIS_IARG_3_WIDTH/8-1:0] ap_axis_iarg_3_tstrb,
    output [S_AXIS_IARG_3_WIDTH-1:0] ap_axis_iarg_3_tdata,
    input ap_axis_iarg_3_tready,
    //input AXI-Stream pass-through interface 4
    input s_axis_iarg_4_aclk,
    input s_axis_iarg_4_aresetn,
    input s_axis_iarg_4_tlast,
    input s_axis_iarg_4_tvalid,
    input [S_AXIS_IARG_4_DMWIDTH/8-1:0] s_axis_iarg_4_tkeep,
    input [S_AXIS_IARG_4_DMWIDTH/8-1:0] s_axis_iarg_4_tstrb,
    input [S_AXIS_IARG_4_DMWIDTH-1:0] s_axis_iarg_4_tdata,
    output s_axis_iarg_4_tready,
    output ap_axis_iarg_4_tlast,
    output ap_axis_iarg_4_tvalid,
    output [S_AXIS_IARG_4_WIDTH/8-1:0] ap_axis_iarg_4_tkeep,
    output [S_AXIS_IARG_4_WIDTH/8-1:0] ap_axis_iarg_4_tstrb,
    output [S_AXIS_IARG_4_WIDTH-1:0] ap_axis_iarg_4_tdata,
    input ap_axis_iarg_4_tready,
    //input AXI-Stream pass-through interface 5
    input s_axis_iarg_5_aclk,
    input s_axis_iarg_5_aresetn,
    input s_axis_iarg_5_tlast,
    input s_axis_iarg_5_tvalid,
    input [S_AXIS_IARG_5_DMWIDTH/8-1:0] s_axis_iarg_5_tkeep,
    input [S_AXIS_IARG_5_DMWIDTH/8-1:0] s_axis_iarg_5_tstrb,
    input [S_AXIS_IARG_5_DMWIDTH-1:0] s_axis_iarg_5_tdata,
    output s_axis_iarg_5_tready,
    output ap_axis_iarg_5_tlast,
    output ap_axis_iarg_5_tvalid,
    output [S_AXIS_IARG_5_WIDTH/8-1:0] ap_axis_iarg_5_tkeep,
    output [S_AXIS_IARG_5_WIDTH/8-1:0] ap_axis_iarg_5_tstrb,
    output [S_AXIS_IARG_5_WIDTH-1:0] ap_axis_iarg_5_tdata,
    input ap_axis_iarg_5_tready,
    //input AXI-Stream pass-through interface 6
    input s_axis_iarg_6_aclk,
    input s_axis_iarg_6_aresetn,
    input s_axis_iarg_6_tlast,
    input s_axis_iarg_6_tvalid,
    input [S_AXIS_IARG_6_DMWIDTH/8-1:0] s_axis_iarg_6_tkeep,
    input [S_AXIS_IARG_6_DMWIDTH/8-1:0] s_axis_iarg_6_tstrb,
    input [S_AXIS_IARG_6_DMWIDTH-1:0] s_axis_iarg_6_tdata,
    output s_axis_iarg_6_tready,
    output ap_axis_iarg_6_tlast,
    output ap_axis_iarg_6_tvalid,
    output [S_AXIS_IARG_6_WIDTH/8-1:0] ap_axis_iarg_6_tkeep,
    output [S_AXIS_IARG_6_WIDTH/8-1:0] ap_axis_iarg_6_tstrb,
    output [S_AXIS_IARG_6_WIDTH-1:0] ap_axis_iarg_6_tdata,
    input ap_axis_iarg_6_tready,
    //input AXI-Stream pass-through interface 7
    input s_axis_iarg_7_aclk,
    input s_axis_iarg_7_aresetn,
    input s_axis_iarg_7_tlast,
    input s_axis_iarg_7_tvalid,
    input [S_AXIS_IARG_7_DMWIDTH/8-1:0] s_axis_iarg_7_tkeep,
    input [S_AXIS_IARG_7_DMWIDTH/8-1:0] s_axis_iarg_7_tstrb,
    input [S_AXIS_IARG_7_DMWIDTH-1:0] s_axis_iarg_7_tdata,
    output s_axis_iarg_7_tready,
    output ap_axis_iarg_7_tlast,
    output ap_axis_iarg_7_tvalid,
    output [S_AXIS_IARG_7_WIDTH/8-1:0] ap_axis_iarg_7_tkeep,
    output [S_AXIS_IARG_7_WIDTH/8-1:0] ap_axis_iarg_7_tstrb,
    output [S_AXIS_IARG_7_WIDTH-1:0] ap_axis_iarg_7_tdata,
    input ap_axis_iarg_7_tready,
    //input AXI-Stream pass-through interface 8
    input s_axis_iarg_8_aclk,
    input s_axis_iarg_8_aresetn,
    input s_axis_iarg_8_tlast,
    input s_axis_iarg_8_tvalid,
    input [S_AXIS_IARG_8_DMWIDTH/8-1:0] s_axis_iarg_8_tkeep,
    input [S_AXIS_IARG_8_DMWIDTH/8-1:0] s_axis_iarg_8_tstrb,
    input [S_AXIS_IARG_8_DMWIDTH-1:0] s_axis_iarg_8_tdata,
    output s_axis_iarg_8_tready,
    output ap_axis_iarg_8_tlast,
    output ap_axis_iarg_8_tvalid,
    output [S_AXIS_IARG_8_WIDTH/8-1:0] ap_axis_iarg_8_tkeep,
    output [S_AXIS_IARG_8_WIDTH/8-1:0] ap_axis_iarg_8_tstrb,
    output [S_AXIS_IARG_8_WIDTH-1:0] ap_axis_iarg_8_tdata,
    input ap_axis_iarg_8_tready,
    //input AXI-Stream pass-through interface 9
    input s_axis_iarg_9_aclk,
    input s_axis_iarg_9_aresetn,
    input s_axis_iarg_9_tlast,
    input s_axis_iarg_9_tvalid,
    input [S_AXIS_IARG_9_DMWIDTH/8-1:0] s_axis_iarg_9_tkeep,
    input [S_AXIS_IARG_9_DMWIDTH/8-1:0] s_axis_iarg_9_tstrb,
    input [S_AXIS_IARG_9_DMWIDTH-1:0] s_axis_iarg_9_tdata,
    output s_axis_iarg_9_tready,
    output ap_axis_iarg_9_tlast,
    output ap_axis_iarg_9_tvalid,
    output [S_AXIS_IARG_9_WIDTH/8-1:0] ap_axis_iarg_9_tkeep,
    output [S_AXIS_IARG_9_WIDTH/8-1:0] ap_axis_iarg_9_tstrb,
    output [S_AXIS_IARG_9_WIDTH-1:0] ap_axis_iarg_9_tdata,
    input ap_axis_iarg_9_tready,
    //input AXI-Stream pass-through interface 10
    input s_axis_iarg_10_aclk,
    input s_axis_iarg_10_aresetn,
    input s_axis_iarg_10_tlast,
    input s_axis_iarg_10_tvalid,
    input [S_AXIS_IARG_10_DMWIDTH/8-1:0] s_axis_iarg_10_tkeep,
    input [S_AXIS_IARG_10_DMWIDTH/8-1:0] s_axis_iarg_10_tstrb,
    input [S_AXIS_IARG_10_DMWIDTH-1:0] s_axis_iarg_10_tdata,
    output s_axis_iarg_10_tready,
    output ap_axis_iarg_10_tlast,
    output ap_axis_iarg_10_tvalid,
    output [S_AXIS_IARG_10_WIDTH/8-1:0] ap_axis_iarg_10_tkeep,
    output [S_AXIS_IARG_10_WIDTH/8-1:0] ap_axis_iarg_10_tstrb,
    output [S_AXIS_IARG_10_WIDTH-1:0] ap_axis_iarg_10_tdata,
    input ap_axis_iarg_10_tready,
    //input AXI-Stream pass-through interface 11
    input s_axis_iarg_11_aclk,
    input s_axis_iarg_11_aresetn,
    input s_axis_iarg_11_tlast,
    input s_axis_iarg_11_tvalid,
    input [S_AXIS_IARG_11_DMWIDTH/8-1:0] s_axis_iarg_11_tkeep,
    input [S_AXIS_IARG_11_DMWIDTH/8-1:0] s_axis_iarg_11_tstrb,
    input [S_AXIS_IARG_11_DMWIDTH-1:0] s_axis_iarg_11_tdata,
    output s_axis_iarg_11_tready,
    output ap_axis_iarg_11_tlast,
    output ap_axis_iarg_11_tvalid,
    output [S_AXIS_IARG_11_WIDTH/8-1:0] ap_axis_iarg_11_tkeep,
    output [S_AXIS_IARG_11_WIDTH/8-1:0] ap_axis_iarg_11_tstrb,
    output [S_AXIS_IARG_11_WIDTH-1:0] ap_axis_iarg_11_tdata,
    input ap_axis_iarg_11_tready,
    //input AXI-Stream pass-through interface 12
    input s_axis_iarg_12_aclk,
    input s_axis_iarg_12_aresetn,
    input s_axis_iarg_12_tlast,
    input s_axis_iarg_12_tvalid,
    input [S_AXIS_IARG_12_DMWIDTH/8-1:0] s_axis_iarg_12_tkeep,
    input [S_AXIS_IARG_12_DMWIDTH/8-1:0] s_axis_iarg_12_tstrb,
    input [S_AXIS_IARG_12_DMWIDTH-1:0] s_axis_iarg_12_tdata,
    output s_axis_iarg_12_tready,
    output ap_axis_iarg_12_tlast,
    output ap_axis_iarg_12_tvalid,
    output [S_AXIS_IARG_12_WIDTH/8-1:0] ap_axis_iarg_12_tkeep,
    output [S_AXIS_IARG_12_WIDTH/8-1:0] ap_axis_iarg_12_tstrb,
    output [S_AXIS_IARG_12_WIDTH-1:0] ap_axis_iarg_12_tdata,
    input ap_axis_iarg_12_tready,
    //input AXI-Stream pass-through interface 13
    input s_axis_iarg_13_aclk,
    input s_axis_iarg_13_aresetn,
    input s_axis_iarg_13_tlast,
    input s_axis_iarg_13_tvalid,
    input [S_AXIS_IARG_13_DMWIDTH/8-1:0] s_axis_iarg_13_tkeep,
    input [S_AXIS_IARG_13_DMWIDTH/8-1:0] s_axis_iarg_13_tstrb,
    input [S_AXIS_IARG_13_DMWIDTH-1:0] s_axis_iarg_13_tdata,
    output s_axis_iarg_13_tready,
    output ap_axis_iarg_13_tlast,
    output ap_axis_iarg_13_tvalid,
    output [S_AXIS_IARG_13_WIDTH/8-1:0] ap_axis_iarg_13_tkeep,
    output [S_AXIS_IARG_13_WIDTH/8-1:0] ap_axis_iarg_13_tstrb,
    output [S_AXIS_IARG_13_WIDTH-1:0] ap_axis_iarg_13_tdata,
    input ap_axis_iarg_13_tready,
    //input AXI-Stream pass-through interface 14
    input s_axis_iarg_14_aclk,
    input s_axis_iarg_14_aresetn,
    input s_axis_iarg_14_tlast,
    input s_axis_iarg_14_tvalid,
    input [S_AXIS_IARG_14_DMWIDTH/8-1:0] s_axis_iarg_14_tkeep,
    input [S_AXIS_IARG_14_DMWIDTH/8-1:0] s_axis_iarg_14_tstrb,
    input [S_AXIS_IARG_14_DMWIDTH-1:0] s_axis_iarg_14_tdata,
    output s_axis_iarg_14_tready,
    output ap_axis_iarg_14_tlast,
    output ap_axis_iarg_14_tvalid,
    output [S_AXIS_IARG_14_WIDTH/8-1:0] ap_axis_iarg_14_tkeep,
    output [S_AXIS_IARG_14_WIDTH/8-1:0] ap_axis_iarg_14_tstrb,
    output [S_AXIS_IARG_14_WIDTH-1:0] ap_axis_iarg_14_tdata,
    input ap_axis_iarg_14_tready,
    //input AXI-Stream pass-through interface 15
    input s_axis_iarg_15_aclk,
    input s_axis_iarg_15_aresetn,
    input s_axis_iarg_15_tlast,
    input s_axis_iarg_15_tvalid,
    input [S_AXIS_IARG_15_DMWIDTH/8-1:0] s_axis_iarg_15_tkeep,
    input [S_AXIS_IARG_15_DMWIDTH/8-1:0] s_axis_iarg_15_tstrb,
    input [S_AXIS_IARG_15_DMWIDTH-1:0] s_axis_iarg_15_tdata,
    output s_axis_iarg_15_tready,
    output ap_axis_iarg_15_tlast,
    output ap_axis_iarg_15_tvalid,
    output [S_AXIS_IARG_15_WIDTH/8-1:0] ap_axis_iarg_15_tkeep,
    output [S_AXIS_IARG_15_WIDTH/8-1:0] ap_axis_iarg_15_tstrb,
    output [S_AXIS_IARG_15_WIDTH-1:0] ap_axis_iarg_15_tdata,
    input ap_axis_iarg_15_tready,
    //input AXI-Stream pass-through interface 16
    input s_axis_iarg_16_aclk,
    input s_axis_iarg_16_aresetn,
    input s_axis_iarg_16_tlast,
    input s_axis_iarg_16_tvalid,
    input [S_AXIS_IARG_16_DMWIDTH/8-1:0] s_axis_iarg_16_tkeep,
    input [S_AXIS_IARG_16_DMWIDTH/8-1:0] s_axis_iarg_16_tstrb,
    input [S_AXIS_IARG_16_DMWIDTH-1:0] s_axis_iarg_16_tdata,
    output s_axis_iarg_16_tready,
    output ap_axis_iarg_16_tlast,
    output ap_axis_iarg_16_tvalid,
    output [S_AXIS_IARG_16_WIDTH/8-1:0] ap_axis_iarg_16_tkeep,
    output [S_AXIS_IARG_16_WIDTH/8-1:0] ap_axis_iarg_16_tstrb,
    output [S_AXIS_IARG_16_WIDTH-1:0] ap_axis_iarg_16_tdata,
    input ap_axis_iarg_16_tready,
    //input AXI-Stream pass-through interface 17
    input s_axis_iarg_17_aclk,
    input s_axis_iarg_17_aresetn,
    input s_axis_iarg_17_tlast,
    input s_axis_iarg_17_tvalid,
    input [S_AXIS_IARG_17_DMWIDTH/8-1:0] s_axis_iarg_17_tkeep,
    input [S_AXIS_IARG_17_DMWIDTH/8-1:0] s_axis_iarg_17_tstrb,
    input [S_AXIS_IARG_17_DMWIDTH-1:0] s_axis_iarg_17_tdata,
    output s_axis_iarg_17_tready,
    output ap_axis_iarg_17_tlast,
    output ap_axis_iarg_17_tvalid,
    output [S_AXIS_IARG_17_WIDTH/8-1:0] ap_axis_iarg_17_tkeep,
    output [S_AXIS_IARG_17_WIDTH/8-1:0] ap_axis_iarg_17_tstrb,
    output [S_AXIS_IARG_17_WIDTH-1:0] ap_axis_iarg_17_tdata,
    input ap_axis_iarg_17_tready,
    //input AXI-Stream pass-through interface 18
    input s_axis_iarg_18_aclk,
    input s_axis_iarg_18_aresetn,
    input s_axis_iarg_18_tlast,
    input s_axis_iarg_18_tvalid,
    input [S_AXIS_IARG_18_DMWIDTH/8-1:0] s_axis_iarg_18_tkeep,
    input [S_AXIS_IARG_18_DMWIDTH/8-1:0] s_axis_iarg_18_tstrb,
    input [S_AXIS_IARG_18_DMWIDTH-1:0] s_axis_iarg_18_tdata,
    output s_axis_iarg_18_tready,
    output ap_axis_iarg_18_tlast,
    output ap_axis_iarg_18_tvalid,
    output [S_AXIS_IARG_18_WIDTH/8-1:0] ap_axis_iarg_18_tkeep,
    output [S_AXIS_IARG_18_WIDTH/8-1:0] ap_axis_iarg_18_tstrb,
    output [S_AXIS_IARG_18_WIDTH-1:0] ap_axis_iarg_18_tdata,
    input ap_axis_iarg_18_tready,
    //input AXI-Stream pass-through interface 19
    input s_axis_iarg_19_aclk,
    input s_axis_iarg_19_aresetn,
    input s_axis_iarg_19_tlast,
    input s_axis_iarg_19_tvalid,
    input [S_AXIS_IARG_19_DMWIDTH/8-1:0] s_axis_iarg_19_tkeep,
    input [S_AXIS_IARG_19_DMWIDTH/8-1:0] s_axis_iarg_19_tstrb,
    input [S_AXIS_IARG_19_DMWIDTH-1:0] s_axis_iarg_19_tdata,
    output s_axis_iarg_19_tready,
    output ap_axis_iarg_19_tlast,
    output ap_axis_iarg_19_tvalid,
    output [S_AXIS_IARG_19_WIDTH/8-1:0] ap_axis_iarg_19_tkeep,
    output [S_AXIS_IARG_19_WIDTH/8-1:0] ap_axis_iarg_19_tstrb,
    output [S_AXIS_IARG_19_WIDTH-1:0] ap_axis_iarg_19_tdata,
    input ap_axis_iarg_19_tready,
    //input AXI-Stream pass-through interface 20
    input s_axis_iarg_20_aclk,
    input s_axis_iarg_20_aresetn,
    input s_axis_iarg_20_tlast,
    input s_axis_iarg_20_tvalid,
    input [S_AXIS_IARG_20_DMWIDTH/8-1:0] s_axis_iarg_20_tkeep,
    input [S_AXIS_IARG_20_DMWIDTH/8-1:0] s_axis_iarg_20_tstrb,
    input [S_AXIS_IARG_20_DMWIDTH-1:0] s_axis_iarg_20_tdata,
    output s_axis_iarg_20_tready,
    output ap_axis_iarg_20_tlast,
    output ap_axis_iarg_20_tvalid,
    output [S_AXIS_IARG_20_WIDTH/8-1:0] ap_axis_iarg_20_tkeep,
    output [S_AXIS_IARG_20_WIDTH/8-1:0] ap_axis_iarg_20_tstrb,
    output [S_AXIS_IARG_20_WIDTH-1:0] ap_axis_iarg_20_tdata,
    input ap_axis_iarg_20_tready,
    //input AXI-Stream pass-through interface 21
    input s_axis_iarg_21_aclk,
    input s_axis_iarg_21_aresetn,
    input s_axis_iarg_21_tlast,
    input s_axis_iarg_21_tvalid,
    input [S_AXIS_IARG_21_DMWIDTH/8-1:0] s_axis_iarg_21_tkeep,
    input [S_AXIS_IARG_21_DMWIDTH/8-1:0] s_axis_iarg_21_tstrb,
    input [S_AXIS_IARG_21_DMWIDTH-1:0] s_axis_iarg_21_tdata,
    output s_axis_iarg_21_tready,
    output ap_axis_iarg_21_tlast,
    output ap_axis_iarg_21_tvalid,
    output [S_AXIS_IARG_21_WIDTH/8-1:0] ap_axis_iarg_21_tkeep,
    output [S_AXIS_IARG_21_WIDTH/8-1:0] ap_axis_iarg_21_tstrb,
    output [S_AXIS_IARG_21_WIDTH-1:0] ap_axis_iarg_21_tdata,
    input ap_axis_iarg_21_tready,
    //input AXI-Stream pass-through interface 22
    input s_axis_iarg_22_aclk,
    input s_axis_iarg_22_aresetn,
    input s_axis_iarg_22_tlast,
    input s_axis_iarg_22_tvalid,
    input [S_AXIS_IARG_22_DMWIDTH/8-1:0] s_axis_iarg_22_tkeep,
    input [S_AXIS_IARG_22_DMWIDTH/8-1:0] s_axis_iarg_22_tstrb,
    input [S_AXIS_IARG_22_DMWIDTH-1:0] s_axis_iarg_22_tdata,
    output s_axis_iarg_22_tready,
    output ap_axis_iarg_22_tlast,
    output ap_axis_iarg_22_tvalid,
    output [S_AXIS_IARG_22_WIDTH/8-1:0] ap_axis_iarg_22_tkeep,
    output [S_AXIS_IARG_22_WIDTH/8-1:0] ap_axis_iarg_22_tstrb,
    output [S_AXIS_IARG_22_WIDTH-1:0] ap_axis_iarg_22_tdata,
    input ap_axis_iarg_22_tready,
    //input AXI-Stream pass-through interface 23
    input s_axis_iarg_23_aclk,
    input s_axis_iarg_23_aresetn,
    input s_axis_iarg_23_tlast,
    input s_axis_iarg_23_tvalid,
    input [S_AXIS_IARG_23_DMWIDTH/8-1:0] s_axis_iarg_23_tkeep,
    input [S_AXIS_IARG_23_DMWIDTH/8-1:0] s_axis_iarg_23_tstrb,
    input [S_AXIS_IARG_23_DMWIDTH-1:0] s_axis_iarg_23_tdata,
    output s_axis_iarg_23_tready,
    output ap_axis_iarg_23_tlast,
    output ap_axis_iarg_23_tvalid,
    output [S_AXIS_IARG_23_WIDTH/8-1:0] ap_axis_iarg_23_tkeep,
    output [S_AXIS_IARG_23_WIDTH/8-1:0] ap_axis_iarg_23_tstrb,
    output [S_AXIS_IARG_23_WIDTH-1:0] ap_axis_iarg_23_tdata,
    input ap_axis_iarg_23_tready,
    //input AXI-Stream pass-through interface 24
    input s_axis_iarg_24_aclk,
    input s_axis_iarg_24_aresetn,
    input s_axis_iarg_24_tlast,
    input s_axis_iarg_24_tvalid,
    input [S_AXIS_IARG_24_DMWIDTH/8-1:0] s_axis_iarg_24_tkeep,
    input [S_AXIS_IARG_24_DMWIDTH/8-1:0] s_axis_iarg_24_tstrb,
    input [S_AXIS_IARG_24_DMWIDTH-1:0] s_axis_iarg_24_tdata,
    output s_axis_iarg_24_tready,
    output ap_axis_iarg_24_tlast,
    output ap_axis_iarg_24_tvalid,
    output [S_AXIS_IARG_24_WIDTH/8-1:0] ap_axis_iarg_24_tkeep,
    output [S_AXIS_IARG_24_WIDTH/8-1:0] ap_axis_iarg_24_tstrb,
    output [S_AXIS_IARG_24_WIDTH-1:0] ap_axis_iarg_24_tdata,
    input ap_axis_iarg_24_tready,
    //input AXI-Stream pass-through interface 25
    input s_axis_iarg_25_aclk,
    input s_axis_iarg_25_aresetn,
    input s_axis_iarg_25_tlast,
    input s_axis_iarg_25_tvalid,
    input [S_AXIS_IARG_25_DMWIDTH/8-1:0] s_axis_iarg_25_tkeep,
    input [S_AXIS_IARG_25_DMWIDTH/8-1:0] s_axis_iarg_25_tstrb,
    input [S_AXIS_IARG_25_DMWIDTH-1:0] s_axis_iarg_25_tdata,
    output s_axis_iarg_25_tready,
    output ap_axis_iarg_25_tlast,
    output ap_axis_iarg_25_tvalid,
    output [S_AXIS_IARG_25_WIDTH/8-1:0] ap_axis_iarg_25_tkeep,
    output [S_AXIS_IARG_25_WIDTH/8-1:0] ap_axis_iarg_25_tstrb,
    output [S_AXIS_IARG_25_WIDTH-1:0] ap_axis_iarg_25_tdata,
    input ap_axis_iarg_25_tready,
    //input AXI-Stream pass-through interface 26
    input s_axis_iarg_26_aclk,
    input s_axis_iarg_26_aresetn,
    input s_axis_iarg_26_tlast,
    input s_axis_iarg_26_tvalid,
    input [S_AXIS_IARG_26_DMWIDTH/8-1:0] s_axis_iarg_26_tkeep,
    input [S_AXIS_IARG_26_DMWIDTH/8-1:0] s_axis_iarg_26_tstrb,
    input [S_AXIS_IARG_26_DMWIDTH-1:0] s_axis_iarg_26_tdata,
    output s_axis_iarg_26_tready,
    output ap_axis_iarg_26_tlast,
    output ap_axis_iarg_26_tvalid,
    output [S_AXIS_IARG_26_WIDTH/8-1:0] ap_axis_iarg_26_tkeep,
    output [S_AXIS_IARG_26_WIDTH/8-1:0] ap_axis_iarg_26_tstrb,
    output [S_AXIS_IARG_26_WIDTH-1:0] ap_axis_iarg_26_tdata,
    input ap_axis_iarg_26_tready,
    //input AXI-Stream pass-through interface 27
    input s_axis_iarg_27_aclk,
    input s_axis_iarg_27_aresetn,
    input s_axis_iarg_27_tlast,
    input s_axis_iarg_27_tvalid,
    input [S_AXIS_IARG_27_DMWIDTH/8-1:0] s_axis_iarg_27_tkeep,
    input [S_AXIS_IARG_27_DMWIDTH/8-1:0] s_axis_iarg_27_tstrb,
    input [S_AXIS_IARG_27_DMWIDTH-1:0] s_axis_iarg_27_tdata,
    output s_axis_iarg_27_tready,
    output ap_axis_iarg_27_tlast,
    output ap_axis_iarg_27_tvalid,
    output [S_AXIS_IARG_27_WIDTH/8-1:0] ap_axis_iarg_27_tkeep,
    output [S_AXIS_IARG_27_WIDTH/8-1:0] ap_axis_iarg_27_tstrb,
    output [S_AXIS_IARG_27_WIDTH-1:0] ap_axis_iarg_27_tdata,
    input ap_axis_iarg_27_tready,
    //input AXI-Stream pass-through interface 28
    input s_axis_iarg_28_aclk,
    input s_axis_iarg_28_aresetn,
    input s_axis_iarg_28_tlast,
    input s_axis_iarg_28_tvalid,
    input [S_AXIS_IARG_28_DMWIDTH/8-1:0] s_axis_iarg_28_tkeep,
    input [S_AXIS_IARG_28_DMWIDTH/8-1:0] s_axis_iarg_28_tstrb,
    input [S_AXIS_IARG_28_DMWIDTH-1:0] s_axis_iarg_28_tdata,
    output s_axis_iarg_28_tready,
    output ap_axis_iarg_28_tlast,
    output ap_axis_iarg_28_tvalid,
    output [S_AXIS_IARG_28_WIDTH/8-1:0] ap_axis_iarg_28_tkeep,
    output [S_AXIS_IARG_28_WIDTH/8-1:0] ap_axis_iarg_28_tstrb,
    output [S_AXIS_IARG_28_WIDTH-1:0] ap_axis_iarg_28_tdata,
    input ap_axis_iarg_28_tready,
    //input AXI-Stream pass-through interface 29
    input s_axis_iarg_29_aclk,
    input s_axis_iarg_29_aresetn,
    input s_axis_iarg_29_tlast,
    input s_axis_iarg_29_tvalid,
    input [S_AXIS_IARG_29_DMWIDTH/8-1:0] s_axis_iarg_29_tkeep,
    input [S_AXIS_IARG_29_DMWIDTH/8-1:0] s_axis_iarg_29_tstrb,
    input [S_AXIS_IARG_29_DMWIDTH-1:0] s_axis_iarg_29_tdata,
    output s_axis_iarg_29_tready,
    output ap_axis_iarg_29_tlast,
    output ap_axis_iarg_29_tvalid,
    output [S_AXIS_IARG_29_WIDTH/8-1:0] ap_axis_iarg_29_tkeep,
    output [S_AXIS_IARG_29_WIDTH/8-1:0] ap_axis_iarg_29_tstrb,
    output [S_AXIS_IARG_29_WIDTH-1:0] ap_axis_iarg_29_tdata,
    input ap_axis_iarg_29_tready,
    //input AXI-Stream pass-through interface 30
    input s_axis_iarg_30_aclk,
    input s_axis_iarg_30_aresetn,
    input s_axis_iarg_30_tlast,
    input s_axis_iarg_30_tvalid,
    input [S_AXIS_IARG_30_DMWIDTH/8-1:0] s_axis_iarg_30_tkeep,
    input [S_AXIS_IARG_30_DMWIDTH/8-1:0] s_axis_iarg_30_tstrb,
    input [S_AXIS_IARG_30_DMWIDTH-1:0] s_axis_iarg_30_tdata,
    output s_axis_iarg_30_tready,
    output ap_axis_iarg_30_tlast,
    output ap_axis_iarg_30_tvalid,
    output [S_AXIS_IARG_30_WIDTH/8-1:0] ap_axis_iarg_30_tkeep,
    output [S_AXIS_IARG_30_WIDTH/8-1:0] ap_axis_iarg_30_tstrb,
    output [S_AXIS_IARG_30_WIDTH-1:0] ap_axis_iarg_30_tdata,
    input ap_axis_iarg_30_tready,
    //input AXI-Stream pass-through interface 31
    input s_axis_iarg_31_aclk,
    input s_axis_iarg_31_aresetn,
    input s_axis_iarg_31_tlast,
    input s_axis_iarg_31_tvalid,
    input [S_AXIS_IARG_31_DMWIDTH/8-1:0] s_axis_iarg_31_tkeep,
    input [S_AXIS_IARG_31_DMWIDTH/8-1:0] s_axis_iarg_31_tstrb,
    input [S_AXIS_IARG_31_DMWIDTH-1:0] s_axis_iarg_31_tdata,
    output s_axis_iarg_31_tready,
    output ap_axis_iarg_31_tlast,
    output ap_axis_iarg_31_tvalid,
    output [S_AXIS_IARG_31_WIDTH/8-1:0] ap_axis_iarg_31_tkeep,
    output [S_AXIS_IARG_31_WIDTH/8-1:0] ap_axis_iarg_31_tstrb,
    output [S_AXIS_IARG_31_WIDTH-1:0] ap_axis_iarg_31_tdata,
    input ap_axis_iarg_31_tready,
    //input AXI-Stream pass-through interface 32
    input s_axis_iarg_32_aclk,
    input s_axis_iarg_32_aresetn,
    input s_axis_iarg_32_tlast,
    input s_axis_iarg_32_tvalid,
    input [S_AXIS_IARG_32_DMWIDTH/8-1:0] s_axis_iarg_32_tkeep,
    input [S_AXIS_IARG_32_DMWIDTH/8-1:0] s_axis_iarg_32_tstrb,
    input [S_AXIS_IARG_32_DMWIDTH-1:0] s_axis_iarg_32_tdata,
    output s_axis_iarg_32_tready,
    output ap_axis_iarg_32_tlast,
    output ap_axis_iarg_32_tvalid,
    output [S_AXIS_IARG_32_WIDTH/8-1:0] ap_axis_iarg_32_tkeep,
    output [S_AXIS_IARG_32_WIDTH/8-1:0] ap_axis_iarg_32_tstrb,
    output [S_AXIS_IARG_32_WIDTH-1:0] ap_axis_iarg_32_tdata,
    input ap_axis_iarg_32_tready,
    //input AXI-Stream pass-through interface 33
    input s_axis_iarg_33_aclk,
    input s_axis_iarg_33_aresetn,
    input s_axis_iarg_33_tlast,
    input s_axis_iarg_33_tvalid,
    input [S_AXIS_IARG_33_DMWIDTH/8-1:0] s_axis_iarg_33_tkeep,
    input [S_AXIS_IARG_33_DMWIDTH/8-1:0] s_axis_iarg_33_tstrb,
    input [S_AXIS_IARG_33_DMWIDTH-1:0] s_axis_iarg_33_tdata,
    output s_axis_iarg_33_tready,
    output ap_axis_iarg_33_tlast,
    output ap_axis_iarg_33_tvalid,
    output [S_AXIS_IARG_33_WIDTH/8-1:0] ap_axis_iarg_33_tkeep,
    output [S_AXIS_IARG_33_WIDTH/8-1:0] ap_axis_iarg_33_tstrb,
    output [S_AXIS_IARG_33_WIDTH-1:0] ap_axis_iarg_33_tdata,
    input ap_axis_iarg_33_tready,
    //input AXI-Stream pass-through interface 34
    input s_axis_iarg_34_aclk,
    input s_axis_iarg_34_aresetn,
    input s_axis_iarg_34_tlast,
    input s_axis_iarg_34_tvalid,
    input [S_AXIS_IARG_34_DMWIDTH/8-1:0] s_axis_iarg_34_tkeep,
    input [S_AXIS_IARG_34_DMWIDTH/8-1:0] s_axis_iarg_34_tstrb,
    input [S_AXIS_IARG_34_DMWIDTH-1:0] s_axis_iarg_34_tdata,
    output s_axis_iarg_34_tready,
    output ap_axis_iarg_34_tlast,
    output ap_axis_iarg_34_tvalid,
    output [S_AXIS_IARG_34_WIDTH/8-1:0] ap_axis_iarg_34_tkeep,
    output [S_AXIS_IARG_34_WIDTH/8-1:0] ap_axis_iarg_34_tstrb,
    output [S_AXIS_IARG_34_WIDTH-1:0] ap_axis_iarg_34_tdata,
    input ap_axis_iarg_34_tready,
    //input AXI-Stream pass-through interface 35
    input s_axis_iarg_35_aclk,
    input s_axis_iarg_35_aresetn,
    input s_axis_iarg_35_tlast,
    input s_axis_iarg_35_tvalid,
    input [S_AXIS_IARG_35_DMWIDTH/8-1:0] s_axis_iarg_35_tkeep,
    input [S_AXIS_IARG_35_DMWIDTH/8-1:0] s_axis_iarg_35_tstrb,
    input [S_AXIS_IARG_35_DMWIDTH-1:0] s_axis_iarg_35_tdata,
    output s_axis_iarg_35_tready,
    output ap_axis_iarg_35_tlast,
    output ap_axis_iarg_35_tvalid,
    output [S_AXIS_IARG_35_WIDTH/8-1:0] ap_axis_iarg_35_tkeep,
    output [S_AXIS_IARG_35_WIDTH/8-1:0] ap_axis_iarg_35_tstrb,
    output [S_AXIS_IARG_35_WIDTH-1:0] ap_axis_iarg_35_tdata,
    input ap_axis_iarg_35_tready,
    //input AXI-Stream pass-through interface 36
    input s_axis_iarg_36_aclk,
    input s_axis_iarg_36_aresetn,
    input s_axis_iarg_36_tlast,
    input s_axis_iarg_36_tvalid,
    input [S_AXIS_IARG_36_DMWIDTH/8-1:0] s_axis_iarg_36_tkeep,
    input [S_AXIS_IARG_36_DMWIDTH/8-1:0] s_axis_iarg_36_tstrb,
    input [S_AXIS_IARG_36_DMWIDTH-1:0] s_axis_iarg_36_tdata,
    output s_axis_iarg_36_tready,
    output ap_axis_iarg_36_tlast,
    output ap_axis_iarg_36_tvalid,
    output [S_AXIS_IARG_36_WIDTH/8-1:0] ap_axis_iarg_36_tkeep,
    output [S_AXIS_IARG_36_WIDTH/8-1:0] ap_axis_iarg_36_tstrb,
    output [S_AXIS_IARG_36_WIDTH-1:0] ap_axis_iarg_36_tdata,
    input ap_axis_iarg_36_tready,
    //input AXI-Stream pass-through interface 37
    input s_axis_iarg_37_aclk,
    input s_axis_iarg_37_aresetn,
    input s_axis_iarg_37_tlast,
    input s_axis_iarg_37_tvalid,
    input [S_AXIS_IARG_37_DMWIDTH/8-1:0] s_axis_iarg_37_tkeep,
    input [S_AXIS_IARG_37_DMWIDTH/8-1:0] s_axis_iarg_37_tstrb,
    input [S_AXIS_IARG_37_DMWIDTH-1:0] s_axis_iarg_37_tdata,
    output s_axis_iarg_37_tready,
    output ap_axis_iarg_37_tlast,
    output ap_axis_iarg_37_tvalid,
    output [S_AXIS_IARG_37_WIDTH/8-1:0] ap_axis_iarg_37_tkeep,
    output [S_AXIS_IARG_37_WIDTH/8-1:0] ap_axis_iarg_37_tstrb,
    output [S_AXIS_IARG_37_WIDTH-1:0] ap_axis_iarg_37_tdata,
    input ap_axis_iarg_37_tready,
    //input AXI-Stream pass-through interface 38
    input s_axis_iarg_38_aclk,
    input s_axis_iarg_38_aresetn,
    input s_axis_iarg_38_tlast,
    input s_axis_iarg_38_tvalid,
    input [S_AXIS_IARG_38_DMWIDTH/8-1:0] s_axis_iarg_38_tkeep,
    input [S_AXIS_IARG_38_DMWIDTH/8-1:0] s_axis_iarg_38_tstrb,
    input [S_AXIS_IARG_38_DMWIDTH-1:0] s_axis_iarg_38_tdata,
    output s_axis_iarg_38_tready,
    output ap_axis_iarg_38_tlast,
    output ap_axis_iarg_38_tvalid,
    output [S_AXIS_IARG_38_WIDTH/8-1:0] ap_axis_iarg_38_tkeep,
    output [S_AXIS_IARG_38_WIDTH/8-1:0] ap_axis_iarg_38_tstrb,
    output [S_AXIS_IARG_38_WIDTH-1:0] ap_axis_iarg_38_tdata,
    input ap_axis_iarg_38_tready,
    //input AXI-Stream pass-through interface 39
    input s_axis_iarg_39_aclk,
    input s_axis_iarg_39_aresetn,
    input s_axis_iarg_39_tlast,
    input s_axis_iarg_39_tvalid,
    input [S_AXIS_IARG_39_DMWIDTH/8-1:0] s_axis_iarg_39_tkeep,
    input [S_AXIS_IARG_39_DMWIDTH/8-1:0] s_axis_iarg_39_tstrb,
    input [S_AXIS_IARG_39_DMWIDTH-1:0] s_axis_iarg_39_tdata,
    output s_axis_iarg_39_tready,
    output ap_axis_iarg_39_tlast,
    output ap_axis_iarg_39_tvalid,
    output [S_AXIS_IARG_39_WIDTH/8-1:0] ap_axis_iarg_39_tkeep,
    output [S_AXIS_IARG_39_WIDTH/8-1:0] ap_axis_iarg_39_tstrb,
    output [S_AXIS_IARG_39_WIDTH-1:0] ap_axis_iarg_39_tdata,
    input ap_axis_iarg_39_tready,
    //input AXI-Stream pass-through interface 40
    input s_axis_iarg_40_aclk,
    input s_axis_iarg_40_aresetn,
    input s_axis_iarg_40_tlast,
    input s_axis_iarg_40_tvalid,
    input [S_AXIS_IARG_40_DMWIDTH/8-1:0] s_axis_iarg_40_tkeep,
    input [S_AXIS_IARG_40_DMWIDTH/8-1:0] s_axis_iarg_40_tstrb,
    input [S_AXIS_IARG_40_DMWIDTH-1:0] s_axis_iarg_40_tdata,
    output s_axis_iarg_40_tready,
    output ap_axis_iarg_40_tlast,
    output ap_axis_iarg_40_tvalid,
    output [S_AXIS_IARG_40_WIDTH/8-1:0] ap_axis_iarg_40_tkeep,
    output [S_AXIS_IARG_40_WIDTH/8-1:0] ap_axis_iarg_40_tstrb,
    output [S_AXIS_IARG_40_WIDTH-1:0] ap_axis_iarg_40_tdata,
    input ap_axis_iarg_40_tready,
    //input AXI-Stream pass-through interface 41
    input s_axis_iarg_41_aclk,
    input s_axis_iarg_41_aresetn,
    input s_axis_iarg_41_tlast,
    input s_axis_iarg_41_tvalid,
    input [S_AXIS_IARG_41_DMWIDTH/8-1:0] s_axis_iarg_41_tkeep,
    input [S_AXIS_IARG_41_DMWIDTH/8-1:0] s_axis_iarg_41_tstrb,
    input [S_AXIS_IARG_41_DMWIDTH-1:0] s_axis_iarg_41_tdata,
    output s_axis_iarg_41_tready,
    output ap_axis_iarg_41_tlast,
    output ap_axis_iarg_41_tvalid,
    output [S_AXIS_IARG_41_WIDTH/8-1:0] ap_axis_iarg_41_tkeep,
    output [S_AXIS_IARG_41_WIDTH/8-1:0] ap_axis_iarg_41_tstrb,
    output [S_AXIS_IARG_41_WIDTH-1:0] ap_axis_iarg_41_tdata,
    input ap_axis_iarg_41_tready,
    //input AXI-Stream pass-through interface 42
    input s_axis_iarg_42_aclk,
    input s_axis_iarg_42_aresetn,
    input s_axis_iarg_42_tlast,
    input s_axis_iarg_42_tvalid,
    input [S_AXIS_IARG_42_DMWIDTH/8-1:0] s_axis_iarg_42_tkeep,
    input [S_AXIS_IARG_42_DMWIDTH/8-1:0] s_axis_iarg_42_tstrb,
    input [S_AXIS_IARG_42_DMWIDTH-1:0] s_axis_iarg_42_tdata,
    output s_axis_iarg_42_tready,
    output ap_axis_iarg_42_tlast,
    output ap_axis_iarg_42_tvalid,
    output [S_AXIS_IARG_42_WIDTH/8-1:0] ap_axis_iarg_42_tkeep,
    output [S_AXIS_IARG_42_WIDTH/8-1:0] ap_axis_iarg_42_tstrb,
    output [S_AXIS_IARG_42_WIDTH-1:0] ap_axis_iarg_42_tdata,
    input ap_axis_iarg_42_tready,
    //input AXI-Stream pass-through interface 43
    input s_axis_iarg_43_aclk,
    input s_axis_iarg_43_aresetn,
    input s_axis_iarg_43_tlast,
    input s_axis_iarg_43_tvalid,
    input [S_AXIS_IARG_43_DMWIDTH/8-1:0] s_axis_iarg_43_tkeep,
    input [S_AXIS_IARG_43_DMWIDTH/8-1:0] s_axis_iarg_43_tstrb,
    input [S_AXIS_IARG_43_DMWIDTH-1:0] s_axis_iarg_43_tdata,
    output s_axis_iarg_43_tready,
    output ap_axis_iarg_43_tlast,
    output ap_axis_iarg_43_tvalid,
    output [S_AXIS_IARG_43_WIDTH/8-1:0] ap_axis_iarg_43_tkeep,
    output [S_AXIS_IARG_43_WIDTH/8-1:0] ap_axis_iarg_43_tstrb,
    output [S_AXIS_IARG_43_WIDTH-1:0] ap_axis_iarg_43_tdata,
    input ap_axis_iarg_43_tready,
    //input AXI-Stream pass-through interface 44
    input s_axis_iarg_44_aclk,
    input s_axis_iarg_44_aresetn,
    input s_axis_iarg_44_tlast,
    input s_axis_iarg_44_tvalid,
    input [S_AXIS_IARG_44_DMWIDTH/8-1:0] s_axis_iarg_44_tkeep,
    input [S_AXIS_IARG_44_DMWIDTH/8-1:0] s_axis_iarg_44_tstrb,
    input [S_AXIS_IARG_44_DMWIDTH-1:0] s_axis_iarg_44_tdata,
    output s_axis_iarg_44_tready,
    output ap_axis_iarg_44_tlast,
    output ap_axis_iarg_44_tvalid,
    output [S_AXIS_IARG_44_WIDTH/8-1:0] ap_axis_iarg_44_tkeep,
    output [S_AXIS_IARG_44_WIDTH/8-1:0] ap_axis_iarg_44_tstrb,
    output [S_AXIS_IARG_44_WIDTH-1:0] ap_axis_iarg_44_tdata,
    input ap_axis_iarg_44_tready,
    //input AXI-Stream pass-through interface 45
    input s_axis_iarg_45_aclk,
    input s_axis_iarg_45_aresetn,
    input s_axis_iarg_45_tlast,
    input s_axis_iarg_45_tvalid,
    input [S_AXIS_IARG_45_DMWIDTH/8-1:0] s_axis_iarg_45_tkeep,
    input [S_AXIS_IARG_45_DMWIDTH/8-1:0] s_axis_iarg_45_tstrb,
    input [S_AXIS_IARG_45_DMWIDTH-1:0] s_axis_iarg_45_tdata,
    output s_axis_iarg_45_tready,
    output ap_axis_iarg_45_tlast,
    output ap_axis_iarg_45_tvalid,
    output [S_AXIS_IARG_45_WIDTH/8-1:0] ap_axis_iarg_45_tkeep,
    output [S_AXIS_IARG_45_WIDTH/8-1:0] ap_axis_iarg_45_tstrb,
    output [S_AXIS_IARG_45_WIDTH-1:0] ap_axis_iarg_45_tdata,
    input ap_axis_iarg_45_tready,
    //input AXI-Stream pass-through interface 46
    input s_axis_iarg_46_aclk,
    input s_axis_iarg_46_aresetn,
    input s_axis_iarg_46_tlast,
    input s_axis_iarg_46_tvalid,
    input [S_AXIS_IARG_46_DMWIDTH/8-1:0] s_axis_iarg_46_tkeep,
    input [S_AXIS_IARG_46_DMWIDTH/8-1:0] s_axis_iarg_46_tstrb,
    input [S_AXIS_IARG_46_DMWIDTH-1:0] s_axis_iarg_46_tdata,
    output s_axis_iarg_46_tready,
    output ap_axis_iarg_46_tlast,
    output ap_axis_iarg_46_tvalid,
    output [S_AXIS_IARG_46_WIDTH/8-1:0] ap_axis_iarg_46_tkeep,
    output [S_AXIS_IARG_46_WIDTH/8-1:0] ap_axis_iarg_46_tstrb,
    output [S_AXIS_IARG_46_WIDTH-1:0] ap_axis_iarg_46_tdata,
    input ap_axis_iarg_46_tready,
    //input AXI-Stream pass-through interface 47
    input s_axis_iarg_47_aclk,
    input s_axis_iarg_47_aresetn,
    input s_axis_iarg_47_tlast,
    input s_axis_iarg_47_tvalid,
    input [S_AXIS_IARG_47_DMWIDTH/8-1:0] s_axis_iarg_47_tkeep,
    input [S_AXIS_IARG_47_DMWIDTH/8-1:0] s_axis_iarg_47_tstrb,
    input [S_AXIS_IARG_47_DMWIDTH-1:0] s_axis_iarg_47_tdata,
    output s_axis_iarg_47_tready,
    output ap_axis_iarg_47_tlast,
    output ap_axis_iarg_47_tvalid,
    output [S_AXIS_IARG_47_WIDTH/8-1:0] ap_axis_iarg_47_tkeep,
    output [S_AXIS_IARG_47_WIDTH/8-1:0] ap_axis_iarg_47_tstrb,
    output [S_AXIS_IARG_47_WIDTH-1:0] ap_axis_iarg_47_tdata,
    input ap_axis_iarg_47_tready,
    //input AXI-Stream pass-through interface 48
    input s_axis_iarg_48_aclk,
    input s_axis_iarg_48_aresetn,
    input s_axis_iarg_48_tlast,
    input s_axis_iarg_48_tvalid,
    input [S_AXIS_IARG_48_DMWIDTH/8-1:0] s_axis_iarg_48_tkeep,
    input [S_AXIS_IARG_48_DMWIDTH/8-1:0] s_axis_iarg_48_tstrb,
    input [S_AXIS_IARG_48_DMWIDTH-1:0] s_axis_iarg_48_tdata,
    output s_axis_iarg_48_tready,
    output ap_axis_iarg_48_tlast,
    output ap_axis_iarg_48_tvalid,
    output [S_AXIS_IARG_48_WIDTH/8-1:0] ap_axis_iarg_48_tkeep,
    output [S_AXIS_IARG_48_WIDTH/8-1:0] ap_axis_iarg_48_tstrb,
    output [S_AXIS_IARG_48_WIDTH-1:0] ap_axis_iarg_48_tdata,
    input ap_axis_iarg_48_tready,
    //input AXI-Stream pass-through interface 49
    input s_axis_iarg_49_aclk,
    input s_axis_iarg_49_aresetn,
    input s_axis_iarg_49_tlast,
    input s_axis_iarg_49_tvalid,
    input [S_AXIS_IARG_49_DMWIDTH/8-1:0] s_axis_iarg_49_tkeep,
    input [S_AXIS_IARG_49_DMWIDTH/8-1:0] s_axis_iarg_49_tstrb,
    input [S_AXIS_IARG_49_DMWIDTH-1:0] s_axis_iarg_49_tdata,
    output s_axis_iarg_49_tready,
    output ap_axis_iarg_49_tlast,
    output ap_axis_iarg_49_tvalid,
    output [S_AXIS_IARG_49_WIDTH/8-1:0] ap_axis_iarg_49_tkeep,
    output [S_AXIS_IARG_49_WIDTH/8-1:0] ap_axis_iarg_49_tstrb,
    output [S_AXIS_IARG_49_WIDTH-1:0] ap_axis_iarg_49_tdata,
    input ap_axis_iarg_49_tready,
    //input AXI-Stream pass-through interface 50
    input s_axis_iarg_50_aclk,
    input s_axis_iarg_50_aresetn,
    input s_axis_iarg_50_tlast,
    input s_axis_iarg_50_tvalid,
    input [S_AXIS_IARG_50_DMWIDTH/8-1:0] s_axis_iarg_50_tkeep,
    input [S_AXIS_IARG_50_DMWIDTH/8-1:0] s_axis_iarg_50_tstrb,
    input [S_AXIS_IARG_50_DMWIDTH-1:0] s_axis_iarg_50_tdata,
    output s_axis_iarg_50_tready,
    output ap_axis_iarg_50_tlast,
    output ap_axis_iarg_50_tvalid,
    output [S_AXIS_IARG_50_WIDTH/8-1:0] ap_axis_iarg_50_tkeep,
    output [S_AXIS_IARG_50_WIDTH/8-1:0] ap_axis_iarg_50_tstrb,
    output [S_AXIS_IARG_50_WIDTH-1:0] ap_axis_iarg_50_tdata,
    input ap_axis_iarg_50_tready,
    //input AXI-Stream pass-through interface 51
    input s_axis_iarg_51_aclk,
    input s_axis_iarg_51_aresetn,
    input s_axis_iarg_51_tlast,
    input s_axis_iarg_51_tvalid,
    input [S_AXIS_IARG_51_DMWIDTH/8-1:0] s_axis_iarg_51_tkeep,
    input [S_AXIS_IARG_51_DMWIDTH/8-1:0] s_axis_iarg_51_tstrb,
    input [S_AXIS_IARG_51_DMWIDTH-1:0] s_axis_iarg_51_tdata,
    output s_axis_iarg_51_tready,
    output ap_axis_iarg_51_tlast,
    output ap_axis_iarg_51_tvalid,
    output [S_AXIS_IARG_51_WIDTH/8-1:0] ap_axis_iarg_51_tkeep,
    output [S_AXIS_IARG_51_WIDTH/8-1:0] ap_axis_iarg_51_tstrb,
    output [S_AXIS_IARG_51_WIDTH-1:0] ap_axis_iarg_51_tdata,
    input ap_axis_iarg_51_tready,
    //input AXI-Stream pass-through interface 52
    input s_axis_iarg_52_aclk,
    input s_axis_iarg_52_aresetn,
    input s_axis_iarg_52_tlast,
    input s_axis_iarg_52_tvalid,
    input [S_AXIS_IARG_52_DMWIDTH/8-1:0] s_axis_iarg_52_tkeep,
    input [S_AXIS_IARG_52_DMWIDTH/8-1:0] s_axis_iarg_52_tstrb,
    input [S_AXIS_IARG_52_DMWIDTH-1:0] s_axis_iarg_52_tdata,
    output s_axis_iarg_52_tready,
    output ap_axis_iarg_52_tlast,
    output ap_axis_iarg_52_tvalid,
    output [S_AXIS_IARG_52_WIDTH/8-1:0] ap_axis_iarg_52_tkeep,
    output [S_AXIS_IARG_52_WIDTH/8-1:0] ap_axis_iarg_52_tstrb,
    output [S_AXIS_IARG_52_WIDTH-1:0] ap_axis_iarg_52_tdata,
    input ap_axis_iarg_52_tready,
    //input AXI-Stream pass-through interface 53
    input s_axis_iarg_53_aclk,
    input s_axis_iarg_53_aresetn,
    input s_axis_iarg_53_tlast,
    input s_axis_iarg_53_tvalid,
    input [S_AXIS_IARG_53_DMWIDTH/8-1:0] s_axis_iarg_53_tkeep,
    input [S_AXIS_IARG_53_DMWIDTH/8-1:0] s_axis_iarg_53_tstrb,
    input [S_AXIS_IARG_53_DMWIDTH-1:0] s_axis_iarg_53_tdata,
    output s_axis_iarg_53_tready,
    output ap_axis_iarg_53_tlast,
    output ap_axis_iarg_53_tvalid,
    output [S_AXIS_IARG_53_WIDTH/8-1:0] ap_axis_iarg_53_tkeep,
    output [S_AXIS_IARG_53_WIDTH/8-1:0] ap_axis_iarg_53_tstrb,
    output [S_AXIS_IARG_53_WIDTH-1:0] ap_axis_iarg_53_tdata,
    input ap_axis_iarg_53_tready,
    //input AXI-Stream pass-through interface 54
    input s_axis_iarg_54_aclk,
    input s_axis_iarg_54_aresetn,
    input s_axis_iarg_54_tlast,
    input s_axis_iarg_54_tvalid,
    input [S_AXIS_IARG_54_DMWIDTH/8-1:0] s_axis_iarg_54_tkeep,
    input [S_AXIS_IARG_54_DMWIDTH/8-1:0] s_axis_iarg_54_tstrb,
    input [S_AXIS_IARG_54_DMWIDTH-1:0] s_axis_iarg_54_tdata,
    output s_axis_iarg_54_tready,
    output ap_axis_iarg_54_tlast,
    output ap_axis_iarg_54_tvalid,
    output [S_AXIS_IARG_54_WIDTH/8-1:0] ap_axis_iarg_54_tkeep,
    output [S_AXIS_IARG_54_WIDTH/8-1:0] ap_axis_iarg_54_tstrb,
    output [S_AXIS_IARG_54_WIDTH-1:0] ap_axis_iarg_54_tdata,
    input ap_axis_iarg_54_tready,
    //input AXI-Stream pass-through interface 55
    input s_axis_iarg_55_aclk,
    input s_axis_iarg_55_aresetn,
    input s_axis_iarg_55_tlast,
    input s_axis_iarg_55_tvalid,
    input [S_AXIS_IARG_55_DMWIDTH/8-1:0] s_axis_iarg_55_tkeep,
    input [S_AXIS_IARG_55_DMWIDTH/8-1:0] s_axis_iarg_55_tstrb,
    input [S_AXIS_IARG_55_DMWIDTH-1:0] s_axis_iarg_55_tdata,
    output s_axis_iarg_55_tready,
    output ap_axis_iarg_55_tlast,
    output ap_axis_iarg_55_tvalid,
    output [S_AXIS_IARG_55_WIDTH/8-1:0] ap_axis_iarg_55_tkeep,
    output [S_AXIS_IARG_55_WIDTH/8-1:0] ap_axis_iarg_55_tstrb,
    output [S_AXIS_IARG_55_WIDTH-1:0] ap_axis_iarg_55_tdata,
    input ap_axis_iarg_55_tready,
    //input AXI-Stream pass-through interface 56
    input s_axis_iarg_56_aclk,
    input s_axis_iarg_56_aresetn,
    input s_axis_iarg_56_tlast,
    input s_axis_iarg_56_tvalid,
    input [S_AXIS_IARG_56_DMWIDTH/8-1:0] s_axis_iarg_56_tkeep,
    input [S_AXIS_IARG_56_DMWIDTH/8-1:0] s_axis_iarg_56_tstrb,
    input [S_AXIS_IARG_56_DMWIDTH-1:0] s_axis_iarg_56_tdata,
    output s_axis_iarg_56_tready,
    output ap_axis_iarg_56_tlast,
    output ap_axis_iarg_56_tvalid,
    output [S_AXIS_IARG_56_WIDTH/8-1:0] ap_axis_iarg_56_tkeep,
    output [S_AXIS_IARG_56_WIDTH/8-1:0] ap_axis_iarg_56_tstrb,
    output [S_AXIS_IARG_56_WIDTH-1:0] ap_axis_iarg_56_tdata,
    input ap_axis_iarg_56_tready,
    //input AXI-Stream pass-through interface 57
    input s_axis_iarg_57_aclk,
    input s_axis_iarg_57_aresetn,
    input s_axis_iarg_57_tlast,
    input s_axis_iarg_57_tvalid,
    input [S_AXIS_IARG_57_DMWIDTH/8-1:0] s_axis_iarg_57_tkeep,
    input [S_AXIS_IARG_57_DMWIDTH/8-1:0] s_axis_iarg_57_tstrb,
    input [S_AXIS_IARG_57_DMWIDTH-1:0] s_axis_iarg_57_tdata,
    output s_axis_iarg_57_tready,
    output ap_axis_iarg_57_tlast,
    output ap_axis_iarg_57_tvalid,
    output [S_AXIS_IARG_57_WIDTH/8-1:0] ap_axis_iarg_57_tkeep,
    output [S_AXIS_IARG_57_WIDTH/8-1:0] ap_axis_iarg_57_tstrb,
    output [S_AXIS_IARG_57_WIDTH-1:0] ap_axis_iarg_57_tdata,
    input ap_axis_iarg_57_tready,
    //input AXI-Stream pass-through interface 58
    input s_axis_iarg_58_aclk,
    input s_axis_iarg_58_aresetn,
    input s_axis_iarg_58_tlast,
    input s_axis_iarg_58_tvalid,
    input [S_AXIS_IARG_58_DMWIDTH/8-1:0] s_axis_iarg_58_tkeep,
    input [S_AXIS_IARG_58_DMWIDTH/8-1:0] s_axis_iarg_58_tstrb,
    input [S_AXIS_IARG_58_DMWIDTH-1:0] s_axis_iarg_58_tdata,
    output s_axis_iarg_58_tready,
    output ap_axis_iarg_58_tlast,
    output ap_axis_iarg_58_tvalid,
    output [S_AXIS_IARG_58_WIDTH/8-1:0] ap_axis_iarg_58_tkeep,
    output [S_AXIS_IARG_58_WIDTH/8-1:0] ap_axis_iarg_58_tstrb,
    output [S_AXIS_IARG_58_WIDTH-1:0] ap_axis_iarg_58_tdata,
    input ap_axis_iarg_58_tready,
    //input AXI-Stream pass-through interface 59
    input s_axis_iarg_59_aclk,
    input s_axis_iarg_59_aresetn,
    input s_axis_iarg_59_tlast,
    input s_axis_iarg_59_tvalid,
    input [S_AXIS_IARG_59_DMWIDTH/8-1:0] s_axis_iarg_59_tkeep,
    input [S_AXIS_IARG_59_DMWIDTH/8-1:0] s_axis_iarg_59_tstrb,
    input [S_AXIS_IARG_59_DMWIDTH-1:0] s_axis_iarg_59_tdata,
    output s_axis_iarg_59_tready,
    output ap_axis_iarg_59_tlast,
    output ap_axis_iarg_59_tvalid,
    output [S_AXIS_IARG_59_WIDTH/8-1:0] ap_axis_iarg_59_tkeep,
    output [S_AXIS_IARG_59_WIDTH/8-1:0] ap_axis_iarg_59_tstrb,
    output [S_AXIS_IARG_59_WIDTH-1:0] ap_axis_iarg_59_tdata,
    input ap_axis_iarg_59_tready,
    //input AXI-Stream pass-through interface 60
    input s_axis_iarg_60_aclk,
    input s_axis_iarg_60_aresetn,
    input s_axis_iarg_60_tlast,
    input s_axis_iarg_60_tvalid,
    input [S_AXIS_IARG_60_DMWIDTH/8-1:0] s_axis_iarg_60_tkeep,
    input [S_AXIS_IARG_60_DMWIDTH/8-1:0] s_axis_iarg_60_tstrb,
    input [S_AXIS_IARG_60_DMWIDTH-1:0] s_axis_iarg_60_tdata,
    output s_axis_iarg_60_tready,
    output ap_axis_iarg_60_tlast,
    output ap_axis_iarg_60_tvalid,
    output [S_AXIS_IARG_60_WIDTH/8-1:0] ap_axis_iarg_60_tkeep,
    output [S_AXIS_IARG_60_WIDTH/8-1:0] ap_axis_iarg_60_tstrb,
    output [S_AXIS_IARG_60_WIDTH-1:0] ap_axis_iarg_60_tdata,
    input ap_axis_iarg_60_tready,
    //input AXI-Stream pass-through interface 61
    input s_axis_iarg_61_aclk,
    input s_axis_iarg_61_aresetn,
    input s_axis_iarg_61_tlast,
    input s_axis_iarg_61_tvalid,
    input [S_AXIS_IARG_61_DMWIDTH/8-1:0] s_axis_iarg_61_tkeep,
    input [S_AXIS_IARG_61_DMWIDTH/8-1:0] s_axis_iarg_61_tstrb,
    input [S_AXIS_IARG_61_DMWIDTH-1:0] s_axis_iarg_61_tdata,
    output s_axis_iarg_61_tready,
    output ap_axis_iarg_61_tlast,
    output ap_axis_iarg_61_tvalid,
    output [S_AXIS_IARG_61_WIDTH/8-1:0] ap_axis_iarg_61_tkeep,
    output [S_AXIS_IARG_61_WIDTH/8-1:0] ap_axis_iarg_61_tstrb,
    output [S_AXIS_IARG_61_WIDTH-1:0] ap_axis_iarg_61_tdata,
    input ap_axis_iarg_61_tready,
    //input AXI-Stream pass-through interface 62
    input s_axis_iarg_62_aclk,
    input s_axis_iarg_62_aresetn,
    input s_axis_iarg_62_tlast,
    input s_axis_iarg_62_tvalid,
    input [S_AXIS_IARG_62_DMWIDTH/8-1:0] s_axis_iarg_62_tkeep,
    input [S_AXIS_IARG_62_DMWIDTH/8-1:0] s_axis_iarg_62_tstrb,
    input [S_AXIS_IARG_62_DMWIDTH-1:0] s_axis_iarg_62_tdata,
    output s_axis_iarg_62_tready,
    output ap_axis_iarg_62_tlast,
    output ap_axis_iarg_62_tvalid,
    output [S_AXIS_IARG_62_WIDTH/8-1:0] ap_axis_iarg_62_tkeep,
    output [S_AXIS_IARG_62_WIDTH/8-1:0] ap_axis_iarg_62_tstrb,
    output [S_AXIS_IARG_62_WIDTH-1:0] ap_axis_iarg_62_tdata,
    input ap_axis_iarg_62_tready,
    //input AXI-Stream pass-through interface 63
    input s_axis_iarg_63_aclk,
    input s_axis_iarg_63_aresetn,
    input s_axis_iarg_63_tlast,
    input s_axis_iarg_63_tvalid,
    input [S_AXIS_IARG_63_DMWIDTH/8-1:0] s_axis_iarg_63_tkeep,
    input [S_AXIS_IARG_63_DMWIDTH/8-1:0] s_axis_iarg_63_tstrb,
    input [S_AXIS_IARG_63_DMWIDTH-1:0] s_axis_iarg_63_tdata,
    output s_axis_iarg_63_tready,
    output ap_axis_iarg_63_tlast,
    output ap_axis_iarg_63_tvalid,
    output [S_AXIS_IARG_63_WIDTH/8-1:0] ap_axis_iarg_63_tkeep,
    output [S_AXIS_IARG_63_WIDTH/8-1:0] ap_axis_iarg_63_tstrb,
    output [S_AXIS_IARG_63_WIDTH-1:0] ap_axis_iarg_63_tdata,
    input ap_axis_iarg_63_tready,
    //input AXI-Stream pass-through interface 64
    input s_axis_iarg_64_aclk,
    input s_axis_iarg_64_aresetn,
    input s_axis_iarg_64_tlast,
    input s_axis_iarg_64_tvalid,
    input [S_AXIS_IARG_64_DMWIDTH/8-1:0] s_axis_iarg_64_tkeep,
    input [S_AXIS_IARG_64_DMWIDTH/8-1:0] s_axis_iarg_64_tstrb,
    input [S_AXIS_IARG_64_DMWIDTH-1:0] s_axis_iarg_64_tdata,
    output s_axis_iarg_64_tready,
    output ap_axis_iarg_64_tlast,
    output ap_axis_iarg_64_tvalid,
    output [S_AXIS_IARG_64_WIDTH/8-1:0] ap_axis_iarg_64_tkeep,
    output [S_AXIS_IARG_64_WIDTH/8-1:0] ap_axis_iarg_64_tstrb,
    output [S_AXIS_IARG_64_WIDTH-1:0] ap_axis_iarg_64_tdata,
    input ap_axis_iarg_64_tready,
    //input AXI-Stream pass-through interface 65
    input s_axis_iarg_65_aclk,
    input s_axis_iarg_65_aresetn,
    input s_axis_iarg_65_tlast,
    input s_axis_iarg_65_tvalid,
    input [S_AXIS_IARG_65_DMWIDTH/8-1:0] s_axis_iarg_65_tkeep,
    input [S_AXIS_IARG_65_DMWIDTH/8-1:0] s_axis_iarg_65_tstrb,
    input [S_AXIS_IARG_65_DMWIDTH-1:0] s_axis_iarg_65_tdata,
    output s_axis_iarg_65_tready,
    output ap_axis_iarg_65_tlast,
    output ap_axis_iarg_65_tvalid,
    output [S_AXIS_IARG_65_WIDTH/8-1:0] ap_axis_iarg_65_tkeep,
    output [S_AXIS_IARG_65_WIDTH/8-1:0] ap_axis_iarg_65_tstrb,
    output [S_AXIS_IARG_65_WIDTH-1:0] ap_axis_iarg_65_tdata,
    input ap_axis_iarg_65_tready,
    //input AXI-Stream pass-through interface 66
    input s_axis_iarg_66_aclk,
    input s_axis_iarg_66_aresetn,
    input s_axis_iarg_66_tlast,
    input s_axis_iarg_66_tvalid,
    input [S_AXIS_IARG_66_DMWIDTH/8-1:0] s_axis_iarg_66_tkeep,
    input [S_AXIS_IARG_66_DMWIDTH/8-1:0] s_axis_iarg_66_tstrb,
    input [S_AXIS_IARG_66_DMWIDTH-1:0] s_axis_iarg_66_tdata,
    output s_axis_iarg_66_tready,
    output ap_axis_iarg_66_tlast,
    output ap_axis_iarg_66_tvalid,
    output [S_AXIS_IARG_66_WIDTH/8-1:0] ap_axis_iarg_66_tkeep,
    output [S_AXIS_IARG_66_WIDTH/8-1:0] ap_axis_iarg_66_tstrb,
    output [S_AXIS_IARG_66_WIDTH-1:0] ap_axis_iarg_66_tdata,
    input ap_axis_iarg_66_tready,
    //input AXI-Stream pass-through interface 67
    input s_axis_iarg_67_aclk,
    input s_axis_iarg_67_aresetn,
    input s_axis_iarg_67_tlast,
    input s_axis_iarg_67_tvalid,
    input [S_AXIS_IARG_67_DMWIDTH/8-1:0] s_axis_iarg_67_tkeep,
    input [S_AXIS_IARG_67_DMWIDTH/8-1:0] s_axis_iarg_67_tstrb,
    input [S_AXIS_IARG_67_DMWIDTH-1:0] s_axis_iarg_67_tdata,
    output s_axis_iarg_67_tready,
    output ap_axis_iarg_67_tlast,
    output ap_axis_iarg_67_tvalid,
    output [S_AXIS_IARG_67_WIDTH/8-1:0] ap_axis_iarg_67_tkeep,
    output [S_AXIS_IARG_67_WIDTH/8-1:0] ap_axis_iarg_67_tstrb,
    output [S_AXIS_IARG_67_WIDTH-1:0] ap_axis_iarg_67_tdata,
    input ap_axis_iarg_67_tready,
    //input AXI-Stream pass-through interface 68
    input s_axis_iarg_68_aclk,
    input s_axis_iarg_68_aresetn,
    input s_axis_iarg_68_tlast,
    input s_axis_iarg_68_tvalid,
    input [S_AXIS_IARG_68_DMWIDTH/8-1:0] s_axis_iarg_68_tkeep,
    input [S_AXIS_IARG_68_DMWIDTH/8-1:0] s_axis_iarg_68_tstrb,
    input [S_AXIS_IARG_68_DMWIDTH-1:0] s_axis_iarg_68_tdata,
    output s_axis_iarg_68_tready,
    output ap_axis_iarg_68_tlast,
    output ap_axis_iarg_68_tvalid,
    output [S_AXIS_IARG_68_WIDTH/8-1:0] ap_axis_iarg_68_tkeep,
    output [S_AXIS_IARG_68_WIDTH/8-1:0] ap_axis_iarg_68_tstrb,
    output [S_AXIS_IARG_68_WIDTH-1:0] ap_axis_iarg_68_tdata,
    input ap_axis_iarg_68_tready,
    //input AXI-Stream pass-through interface 69
    input s_axis_iarg_69_aclk,
    input s_axis_iarg_69_aresetn,
    input s_axis_iarg_69_tlast,
    input s_axis_iarg_69_tvalid,
    input [S_AXIS_IARG_69_DMWIDTH/8-1:0] s_axis_iarg_69_tkeep,
    input [S_AXIS_IARG_69_DMWIDTH/8-1:0] s_axis_iarg_69_tstrb,
    input [S_AXIS_IARG_69_DMWIDTH-1:0] s_axis_iarg_69_tdata,
    output s_axis_iarg_69_tready,
    output ap_axis_iarg_69_tlast,
    output ap_axis_iarg_69_tvalid,
    output [S_AXIS_IARG_69_WIDTH/8-1:0] ap_axis_iarg_69_tkeep,
    output [S_AXIS_IARG_69_WIDTH/8-1:0] ap_axis_iarg_69_tstrb,
    output [S_AXIS_IARG_69_WIDTH-1:0] ap_axis_iarg_69_tdata,
    input ap_axis_iarg_69_tready,
    //input AXI-Stream pass-through interface 70
    input s_axis_iarg_70_aclk,
    input s_axis_iarg_70_aresetn,
    input s_axis_iarg_70_tlast,
    input s_axis_iarg_70_tvalid,
    input [S_AXIS_IARG_70_DMWIDTH/8-1:0] s_axis_iarg_70_tkeep,
    input [S_AXIS_IARG_70_DMWIDTH/8-1:0] s_axis_iarg_70_tstrb,
    input [S_AXIS_IARG_70_DMWIDTH-1:0] s_axis_iarg_70_tdata,
    output s_axis_iarg_70_tready,
    output ap_axis_iarg_70_tlast,
    output ap_axis_iarg_70_tvalid,
    output [S_AXIS_IARG_70_WIDTH/8-1:0] ap_axis_iarg_70_tkeep,
    output [S_AXIS_IARG_70_WIDTH/8-1:0] ap_axis_iarg_70_tstrb,
    output [S_AXIS_IARG_70_WIDTH-1:0] ap_axis_iarg_70_tdata,
    input ap_axis_iarg_70_tready,
    //input AXI-Stream pass-through interface 71
    input s_axis_iarg_71_aclk,
    input s_axis_iarg_71_aresetn,
    input s_axis_iarg_71_tlast,
    input s_axis_iarg_71_tvalid,
    input [S_AXIS_IARG_71_DMWIDTH/8-1:0] s_axis_iarg_71_tkeep,
    input [S_AXIS_IARG_71_DMWIDTH/8-1:0] s_axis_iarg_71_tstrb,
    input [S_AXIS_IARG_71_DMWIDTH-1:0] s_axis_iarg_71_tdata,
    output s_axis_iarg_71_tready,
    output ap_axis_iarg_71_tlast,
    output ap_axis_iarg_71_tvalid,
    output [S_AXIS_IARG_71_WIDTH/8-1:0] ap_axis_iarg_71_tkeep,
    output [S_AXIS_IARG_71_WIDTH/8-1:0] ap_axis_iarg_71_tstrb,
    output [S_AXIS_IARG_71_WIDTH-1:0] ap_axis_iarg_71_tdata,
    input ap_axis_iarg_71_tready,
    //input AXI-Stream pass-through interface 72
    input s_axis_iarg_72_aclk,
    input s_axis_iarg_72_aresetn,
    input s_axis_iarg_72_tlast,
    input s_axis_iarg_72_tvalid,
    input [S_AXIS_IARG_72_DMWIDTH/8-1:0] s_axis_iarg_72_tkeep,
    input [S_AXIS_IARG_72_DMWIDTH/8-1:0] s_axis_iarg_72_tstrb,
    input [S_AXIS_IARG_72_DMWIDTH-1:0] s_axis_iarg_72_tdata,
    output s_axis_iarg_72_tready,
    output ap_axis_iarg_72_tlast,
    output ap_axis_iarg_72_tvalid,
    output [S_AXIS_IARG_72_WIDTH/8-1:0] ap_axis_iarg_72_tkeep,
    output [S_AXIS_IARG_72_WIDTH/8-1:0] ap_axis_iarg_72_tstrb,
    output [S_AXIS_IARG_72_WIDTH-1:0] ap_axis_iarg_72_tdata,
    input ap_axis_iarg_72_tready,
    //input AXI-Stream pass-through interface 73
    input s_axis_iarg_73_aclk,
    input s_axis_iarg_73_aresetn,
    input s_axis_iarg_73_tlast,
    input s_axis_iarg_73_tvalid,
    input [S_AXIS_IARG_73_DMWIDTH/8-1:0] s_axis_iarg_73_tkeep,
    input [S_AXIS_IARG_73_DMWIDTH/8-1:0] s_axis_iarg_73_tstrb,
    input [S_AXIS_IARG_73_DMWIDTH-1:0] s_axis_iarg_73_tdata,
    output s_axis_iarg_73_tready,
    output ap_axis_iarg_73_tlast,
    output ap_axis_iarg_73_tvalid,
    output [S_AXIS_IARG_73_WIDTH/8-1:0] ap_axis_iarg_73_tkeep,
    output [S_AXIS_IARG_73_WIDTH/8-1:0] ap_axis_iarg_73_tstrb,
    output [S_AXIS_IARG_73_WIDTH-1:0] ap_axis_iarg_73_tdata,
    input ap_axis_iarg_73_tready,
    //input AXI-Stream pass-through interface 74
    input s_axis_iarg_74_aclk,
    input s_axis_iarg_74_aresetn,
    input s_axis_iarg_74_tlast,
    input s_axis_iarg_74_tvalid,
    input [S_AXIS_IARG_74_DMWIDTH/8-1:0] s_axis_iarg_74_tkeep,
    input [S_AXIS_IARG_74_DMWIDTH/8-1:0] s_axis_iarg_74_tstrb,
    input [S_AXIS_IARG_74_DMWIDTH-1:0] s_axis_iarg_74_tdata,
    output s_axis_iarg_74_tready,
    output ap_axis_iarg_74_tlast,
    output ap_axis_iarg_74_tvalid,
    output [S_AXIS_IARG_74_WIDTH/8-1:0] ap_axis_iarg_74_tkeep,
    output [S_AXIS_IARG_74_WIDTH/8-1:0] ap_axis_iarg_74_tstrb,
    output [S_AXIS_IARG_74_WIDTH-1:0] ap_axis_iarg_74_tdata,
    input ap_axis_iarg_74_tready,
    //input AXI-Stream pass-through interface 75
    input s_axis_iarg_75_aclk,
    input s_axis_iarg_75_aresetn,
    input s_axis_iarg_75_tlast,
    input s_axis_iarg_75_tvalid,
    input [S_AXIS_IARG_75_DMWIDTH/8-1:0] s_axis_iarg_75_tkeep,
    input [S_AXIS_IARG_75_DMWIDTH/8-1:0] s_axis_iarg_75_tstrb,
    input [S_AXIS_IARG_75_DMWIDTH-1:0] s_axis_iarg_75_tdata,
    output s_axis_iarg_75_tready,
    output ap_axis_iarg_75_tlast,
    output ap_axis_iarg_75_tvalid,
    output [S_AXIS_IARG_75_WIDTH/8-1:0] ap_axis_iarg_75_tkeep,
    output [S_AXIS_IARG_75_WIDTH/8-1:0] ap_axis_iarg_75_tstrb,
    output [S_AXIS_IARG_75_WIDTH-1:0] ap_axis_iarg_75_tdata,
    input ap_axis_iarg_75_tready,
    //input AXI-Stream pass-through interface 76
    input s_axis_iarg_76_aclk,
    input s_axis_iarg_76_aresetn,
    input s_axis_iarg_76_tlast,
    input s_axis_iarg_76_tvalid,
    input [S_AXIS_IARG_76_DMWIDTH/8-1:0] s_axis_iarg_76_tkeep,
    input [S_AXIS_IARG_76_DMWIDTH/8-1:0] s_axis_iarg_76_tstrb,
    input [S_AXIS_IARG_76_DMWIDTH-1:0] s_axis_iarg_76_tdata,
    output s_axis_iarg_76_tready,
    output ap_axis_iarg_76_tlast,
    output ap_axis_iarg_76_tvalid,
    output [S_AXIS_IARG_76_WIDTH/8-1:0] ap_axis_iarg_76_tkeep,
    output [S_AXIS_IARG_76_WIDTH/8-1:0] ap_axis_iarg_76_tstrb,
    output [S_AXIS_IARG_76_WIDTH-1:0] ap_axis_iarg_76_tdata,
    input ap_axis_iarg_76_tready,
    //input AXI-Stream pass-through interface 77
    input s_axis_iarg_77_aclk,
    input s_axis_iarg_77_aresetn,
    input s_axis_iarg_77_tlast,
    input s_axis_iarg_77_tvalid,
    input [S_AXIS_IARG_77_DMWIDTH/8-1:0] s_axis_iarg_77_tkeep,
    input [S_AXIS_IARG_77_DMWIDTH/8-1:0] s_axis_iarg_77_tstrb,
    input [S_AXIS_IARG_77_DMWIDTH-1:0] s_axis_iarg_77_tdata,
    output s_axis_iarg_77_tready,
    output ap_axis_iarg_77_tlast,
    output ap_axis_iarg_77_tvalid,
    output [S_AXIS_IARG_77_WIDTH/8-1:0] ap_axis_iarg_77_tkeep,
    output [S_AXIS_IARG_77_WIDTH/8-1:0] ap_axis_iarg_77_tstrb,
    output [S_AXIS_IARG_77_WIDTH-1:0] ap_axis_iarg_77_tdata,
    input ap_axis_iarg_77_tready,
    //input AXI-Stream pass-through interface 78
    input s_axis_iarg_78_aclk,
    input s_axis_iarg_78_aresetn,
    input s_axis_iarg_78_tlast,
    input s_axis_iarg_78_tvalid,
    input [S_AXIS_IARG_78_DMWIDTH/8-1:0] s_axis_iarg_78_tkeep,
    input [S_AXIS_IARG_78_DMWIDTH/8-1:0] s_axis_iarg_78_tstrb,
    input [S_AXIS_IARG_78_DMWIDTH-1:0] s_axis_iarg_78_tdata,
    output s_axis_iarg_78_tready,
    output ap_axis_iarg_78_tlast,
    output ap_axis_iarg_78_tvalid,
    output [S_AXIS_IARG_78_WIDTH/8-1:0] ap_axis_iarg_78_tkeep,
    output [S_AXIS_IARG_78_WIDTH/8-1:0] ap_axis_iarg_78_tstrb,
    output [S_AXIS_IARG_78_WIDTH-1:0] ap_axis_iarg_78_tdata,
    input ap_axis_iarg_78_tready,
    //input AXI-Stream pass-through interface 79
    input s_axis_iarg_79_aclk,
    input s_axis_iarg_79_aresetn,
    input s_axis_iarg_79_tlast,
    input s_axis_iarg_79_tvalid,
    input [S_AXIS_IARG_79_DMWIDTH/8-1:0] s_axis_iarg_79_tkeep,
    input [S_AXIS_IARG_79_DMWIDTH/8-1:0] s_axis_iarg_79_tstrb,
    input [S_AXIS_IARG_79_DMWIDTH-1:0] s_axis_iarg_79_tdata,
    output s_axis_iarg_79_tready,
    output ap_axis_iarg_79_tlast,
    output ap_axis_iarg_79_tvalid,
    output [S_AXIS_IARG_79_WIDTH/8-1:0] ap_axis_iarg_79_tkeep,
    output [S_AXIS_IARG_79_WIDTH/8-1:0] ap_axis_iarg_79_tstrb,
    output [S_AXIS_IARG_79_WIDTH-1:0] ap_axis_iarg_79_tdata,
    input ap_axis_iarg_79_tready,
    //input AXI-Stream pass-through interface 80
    input s_axis_iarg_80_aclk,
    input s_axis_iarg_80_aresetn,
    input s_axis_iarg_80_tlast,
    input s_axis_iarg_80_tvalid,
    input [S_AXIS_IARG_80_DMWIDTH/8-1:0] s_axis_iarg_80_tkeep,
    input [S_AXIS_IARG_80_DMWIDTH/8-1:0] s_axis_iarg_80_tstrb,
    input [S_AXIS_IARG_80_DMWIDTH-1:0] s_axis_iarg_80_tdata,
    output s_axis_iarg_80_tready,
    output ap_axis_iarg_80_tlast,
    output ap_axis_iarg_80_tvalid,
    output [S_AXIS_IARG_80_WIDTH/8-1:0] ap_axis_iarg_80_tkeep,
    output [S_AXIS_IARG_80_WIDTH/8-1:0] ap_axis_iarg_80_tstrb,
    output [S_AXIS_IARG_80_WIDTH-1:0] ap_axis_iarg_80_tdata,
    input ap_axis_iarg_80_tready,
    //input AXI-Stream pass-through interface 81
    input s_axis_iarg_81_aclk,
    input s_axis_iarg_81_aresetn,
    input s_axis_iarg_81_tlast,
    input s_axis_iarg_81_tvalid,
    input [S_AXIS_IARG_81_DMWIDTH/8-1:0] s_axis_iarg_81_tkeep,
    input [S_AXIS_IARG_81_DMWIDTH/8-1:0] s_axis_iarg_81_tstrb,
    input [S_AXIS_IARG_81_DMWIDTH-1:0] s_axis_iarg_81_tdata,
    output s_axis_iarg_81_tready,
    output ap_axis_iarg_81_tlast,
    output ap_axis_iarg_81_tvalid,
    output [S_AXIS_IARG_81_WIDTH/8-1:0] ap_axis_iarg_81_tkeep,
    output [S_AXIS_IARG_81_WIDTH/8-1:0] ap_axis_iarg_81_tstrb,
    output [S_AXIS_IARG_81_WIDTH-1:0] ap_axis_iarg_81_tdata,
    input ap_axis_iarg_81_tready,
    //input AXI-Stream pass-through interface 82
    input s_axis_iarg_82_aclk,
    input s_axis_iarg_82_aresetn,
    input s_axis_iarg_82_tlast,
    input s_axis_iarg_82_tvalid,
    input [S_AXIS_IARG_82_DMWIDTH/8-1:0] s_axis_iarg_82_tkeep,
    input [S_AXIS_IARG_82_DMWIDTH/8-1:0] s_axis_iarg_82_tstrb,
    input [S_AXIS_IARG_82_DMWIDTH-1:0] s_axis_iarg_82_tdata,
    output s_axis_iarg_82_tready,
    output ap_axis_iarg_82_tlast,
    output ap_axis_iarg_82_tvalid,
    output [S_AXIS_IARG_82_WIDTH/8-1:0] ap_axis_iarg_82_tkeep,
    output [S_AXIS_IARG_82_WIDTH/8-1:0] ap_axis_iarg_82_tstrb,
    output [S_AXIS_IARG_82_WIDTH-1:0] ap_axis_iarg_82_tdata,
    input ap_axis_iarg_82_tready,
    //input AXI-Stream pass-through interface 83
    input s_axis_iarg_83_aclk,
    input s_axis_iarg_83_aresetn,
    input s_axis_iarg_83_tlast,
    input s_axis_iarg_83_tvalid,
    input [S_AXIS_IARG_83_DMWIDTH/8-1:0] s_axis_iarg_83_tkeep,
    input [S_AXIS_IARG_83_DMWIDTH/8-1:0] s_axis_iarg_83_tstrb,
    input [S_AXIS_IARG_83_DMWIDTH-1:0] s_axis_iarg_83_tdata,
    output s_axis_iarg_83_tready,
    output ap_axis_iarg_83_tlast,
    output ap_axis_iarg_83_tvalid,
    output [S_AXIS_IARG_83_WIDTH/8-1:0] ap_axis_iarg_83_tkeep,
    output [S_AXIS_IARG_83_WIDTH/8-1:0] ap_axis_iarg_83_tstrb,
    output [S_AXIS_IARG_83_WIDTH-1:0] ap_axis_iarg_83_tdata,
    input ap_axis_iarg_83_tready,
    //input AXI-Stream pass-through interface 84
    input s_axis_iarg_84_aclk,
    input s_axis_iarg_84_aresetn,
    input s_axis_iarg_84_tlast,
    input s_axis_iarg_84_tvalid,
    input [S_AXIS_IARG_84_DMWIDTH/8-1:0] s_axis_iarg_84_tkeep,
    input [S_AXIS_IARG_84_DMWIDTH/8-1:0] s_axis_iarg_84_tstrb,
    input [S_AXIS_IARG_84_DMWIDTH-1:0] s_axis_iarg_84_tdata,
    output s_axis_iarg_84_tready,
    output ap_axis_iarg_84_tlast,
    output ap_axis_iarg_84_tvalid,
    output [S_AXIS_IARG_84_WIDTH/8-1:0] ap_axis_iarg_84_tkeep,
    output [S_AXIS_IARG_84_WIDTH/8-1:0] ap_axis_iarg_84_tstrb,
    output [S_AXIS_IARG_84_WIDTH-1:0] ap_axis_iarg_84_tdata,
    input ap_axis_iarg_84_tready,
    //input AXI-Stream pass-through interface 85
    input s_axis_iarg_85_aclk,
    input s_axis_iarg_85_aresetn,
    input s_axis_iarg_85_tlast,
    input s_axis_iarg_85_tvalid,
    input [S_AXIS_IARG_85_DMWIDTH/8-1:0] s_axis_iarg_85_tkeep,
    input [S_AXIS_IARG_85_DMWIDTH/8-1:0] s_axis_iarg_85_tstrb,
    input [S_AXIS_IARG_85_DMWIDTH-1:0] s_axis_iarg_85_tdata,
    output s_axis_iarg_85_tready,
    output ap_axis_iarg_85_tlast,
    output ap_axis_iarg_85_tvalid,
    output [S_AXIS_IARG_85_WIDTH/8-1:0] ap_axis_iarg_85_tkeep,
    output [S_AXIS_IARG_85_WIDTH/8-1:0] ap_axis_iarg_85_tstrb,
    output [S_AXIS_IARG_85_WIDTH-1:0] ap_axis_iarg_85_tdata,
    input ap_axis_iarg_85_tready,
    //input AXI-Stream pass-through interface 86
    input s_axis_iarg_86_aclk,
    input s_axis_iarg_86_aresetn,
    input s_axis_iarg_86_tlast,
    input s_axis_iarg_86_tvalid,
    input [S_AXIS_IARG_86_DMWIDTH/8-1:0] s_axis_iarg_86_tkeep,
    input [S_AXIS_IARG_86_DMWIDTH/8-1:0] s_axis_iarg_86_tstrb,
    input [S_AXIS_IARG_86_DMWIDTH-1:0] s_axis_iarg_86_tdata,
    output s_axis_iarg_86_tready,
    output ap_axis_iarg_86_tlast,
    output ap_axis_iarg_86_tvalid,
    output [S_AXIS_IARG_86_WIDTH/8-1:0] ap_axis_iarg_86_tkeep,
    output [S_AXIS_IARG_86_WIDTH/8-1:0] ap_axis_iarg_86_tstrb,
    output [S_AXIS_IARG_86_WIDTH-1:0] ap_axis_iarg_86_tdata,
    input ap_axis_iarg_86_tready,
    //input AXI-Stream pass-through interface 87
    input s_axis_iarg_87_aclk,
    input s_axis_iarg_87_aresetn,
    input s_axis_iarg_87_tlast,
    input s_axis_iarg_87_tvalid,
    input [S_AXIS_IARG_87_DMWIDTH/8-1:0] s_axis_iarg_87_tkeep,
    input [S_AXIS_IARG_87_DMWIDTH/8-1:0] s_axis_iarg_87_tstrb,
    input [S_AXIS_IARG_87_DMWIDTH-1:0] s_axis_iarg_87_tdata,
    output s_axis_iarg_87_tready,
    output ap_axis_iarg_87_tlast,
    output ap_axis_iarg_87_tvalid,
    output [S_AXIS_IARG_87_WIDTH/8-1:0] ap_axis_iarg_87_tkeep,
    output [S_AXIS_IARG_87_WIDTH/8-1:0] ap_axis_iarg_87_tstrb,
    output [S_AXIS_IARG_87_WIDTH-1:0] ap_axis_iarg_87_tdata,
    input ap_axis_iarg_87_tready,
    //input AXI-Stream pass-through interface 88
    input s_axis_iarg_88_aclk,
    input s_axis_iarg_88_aresetn,
    input s_axis_iarg_88_tlast,
    input s_axis_iarg_88_tvalid,
    input [S_AXIS_IARG_88_DMWIDTH/8-1:0] s_axis_iarg_88_tkeep,
    input [S_AXIS_IARG_88_DMWIDTH/8-1:0] s_axis_iarg_88_tstrb,
    input [S_AXIS_IARG_88_DMWIDTH-1:0] s_axis_iarg_88_tdata,
    output s_axis_iarg_88_tready,
    output ap_axis_iarg_88_tlast,
    output ap_axis_iarg_88_tvalid,
    output [S_AXIS_IARG_88_WIDTH/8-1:0] ap_axis_iarg_88_tkeep,
    output [S_AXIS_IARG_88_WIDTH/8-1:0] ap_axis_iarg_88_tstrb,
    output [S_AXIS_IARG_88_WIDTH-1:0] ap_axis_iarg_88_tdata,
    input ap_axis_iarg_88_tready,
    //input AXI-Stream pass-through interface 89
    input s_axis_iarg_89_aclk,
    input s_axis_iarg_89_aresetn,
    input s_axis_iarg_89_tlast,
    input s_axis_iarg_89_tvalid,
    input [S_AXIS_IARG_89_DMWIDTH/8-1:0] s_axis_iarg_89_tkeep,
    input [S_AXIS_IARG_89_DMWIDTH/8-1:0] s_axis_iarg_89_tstrb,
    input [S_AXIS_IARG_89_DMWIDTH-1:0] s_axis_iarg_89_tdata,
    output s_axis_iarg_89_tready,
    output ap_axis_iarg_89_tlast,
    output ap_axis_iarg_89_tvalid,
    output [S_AXIS_IARG_89_WIDTH/8-1:0] ap_axis_iarg_89_tkeep,
    output [S_AXIS_IARG_89_WIDTH/8-1:0] ap_axis_iarg_89_tstrb,
    output [S_AXIS_IARG_89_WIDTH-1:0] ap_axis_iarg_89_tdata,
    input ap_axis_iarg_89_tready,
    //input AXI-Stream pass-through interface 90
    input s_axis_iarg_90_aclk,
    input s_axis_iarg_90_aresetn,
    input s_axis_iarg_90_tlast,
    input s_axis_iarg_90_tvalid,
    input [S_AXIS_IARG_90_DMWIDTH/8-1:0] s_axis_iarg_90_tkeep,
    input [S_AXIS_IARG_90_DMWIDTH/8-1:0] s_axis_iarg_90_tstrb,
    input [S_AXIS_IARG_90_DMWIDTH-1:0] s_axis_iarg_90_tdata,
    output s_axis_iarg_90_tready,
    output ap_axis_iarg_90_tlast,
    output ap_axis_iarg_90_tvalid,
    output [S_AXIS_IARG_90_WIDTH/8-1:0] ap_axis_iarg_90_tkeep,
    output [S_AXIS_IARG_90_WIDTH/8-1:0] ap_axis_iarg_90_tstrb,
    output [S_AXIS_IARG_90_WIDTH-1:0] ap_axis_iarg_90_tdata,
    input ap_axis_iarg_90_tready,
    //input AXI-Stream pass-through interface 91
    input s_axis_iarg_91_aclk,
    input s_axis_iarg_91_aresetn,
    input s_axis_iarg_91_tlast,
    input s_axis_iarg_91_tvalid,
    input [S_AXIS_IARG_91_DMWIDTH/8-1:0] s_axis_iarg_91_tkeep,
    input [S_AXIS_IARG_91_DMWIDTH/8-1:0] s_axis_iarg_91_tstrb,
    input [S_AXIS_IARG_91_DMWIDTH-1:0] s_axis_iarg_91_tdata,
    output s_axis_iarg_91_tready,
    output ap_axis_iarg_91_tlast,
    output ap_axis_iarg_91_tvalid,
    output [S_AXIS_IARG_91_WIDTH/8-1:0] ap_axis_iarg_91_tkeep,
    output [S_AXIS_IARG_91_WIDTH/8-1:0] ap_axis_iarg_91_tstrb,
    output [S_AXIS_IARG_91_WIDTH-1:0] ap_axis_iarg_91_tdata,
    input ap_axis_iarg_91_tready,
    //input AXI-Stream pass-through interface 92
    input s_axis_iarg_92_aclk,
    input s_axis_iarg_92_aresetn,
    input s_axis_iarg_92_tlast,
    input s_axis_iarg_92_tvalid,
    input [S_AXIS_IARG_92_DMWIDTH/8-1:0] s_axis_iarg_92_tkeep,
    input [S_AXIS_IARG_92_DMWIDTH/8-1:0] s_axis_iarg_92_tstrb,
    input [S_AXIS_IARG_92_DMWIDTH-1:0] s_axis_iarg_92_tdata,
    output s_axis_iarg_92_tready,
    output ap_axis_iarg_92_tlast,
    output ap_axis_iarg_92_tvalid,
    output [S_AXIS_IARG_92_WIDTH/8-1:0] ap_axis_iarg_92_tkeep,
    output [S_AXIS_IARG_92_WIDTH/8-1:0] ap_axis_iarg_92_tstrb,
    output [S_AXIS_IARG_92_WIDTH-1:0] ap_axis_iarg_92_tdata,
    input ap_axis_iarg_92_tready,
    //input AXI-Stream pass-through interface 93
    input s_axis_iarg_93_aclk,
    input s_axis_iarg_93_aresetn,
    input s_axis_iarg_93_tlast,
    input s_axis_iarg_93_tvalid,
    input [S_AXIS_IARG_93_DMWIDTH/8-1:0] s_axis_iarg_93_tkeep,
    input [S_AXIS_IARG_93_DMWIDTH/8-1:0] s_axis_iarg_93_tstrb,
    input [S_AXIS_IARG_93_DMWIDTH-1:0] s_axis_iarg_93_tdata,
    output s_axis_iarg_93_tready,
    output ap_axis_iarg_93_tlast,
    output ap_axis_iarg_93_tvalid,
    output [S_AXIS_IARG_93_WIDTH/8-1:0] ap_axis_iarg_93_tkeep,
    output [S_AXIS_IARG_93_WIDTH/8-1:0] ap_axis_iarg_93_tstrb,
    output [S_AXIS_IARG_93_WIDTH-1:0] ap_axis_iarg_93_tdata,
    input ap_axis_iarg_93_tready,
    //input AXI-Stream pass-through interface 94
    input s_axis_iarg_94_aclk,
    input s_axis_iarg_94_aresetn,
    input s_axis_iarg_94_tlast,
    input s_axis_iarg_94_tvalid,
    input [S_AXIS_IARG_94_DMWIDTH/8-1:0] s_axis_iarg_94_tkeep,
    input [S_AXIS_IARG_94_DMWIDTH/8-1:0] s_axis_iarg_94_tstrb,
    input [S_AXIS_IARG_94_DMWIDTH-1:0] s_axis_iarg_94_tdata,
    output s_axis_iarg_94_tready,
    output ap_axis_iarg_94_tlast,
    output ap_axis_iarg_94_tvalid,
    output [S_AXIS_IARG_94_WIDTH/8-1:0] ap_axis_iarg_94_tkeep,
    output [S_AXIS_IARG_94_WIDTH/8-1:0] ap_axis_iarg_94_tstrb,
    output [S_AXIS_IARG_94_WIDTH-1:0] ap_axis_iarg_94_tdata,
    input ap_axis_iarg_94_tready,
    //input AXI-Stream pass-through interface 95
    input s_axis_iarg_95_aclk,
    input s_axis_iarg_95_aresetn,
    input s_axis_iarg_95_tlast,
    input s_axis_iarg_95_tvalid,
    input [S_AXIS_IARG_95_DMWIDTH/8-1:0] s_axis_iarg_95_tkeep,
    input [S_AXIS_IARG_95_DMWIDTH/8-1:0] s_axis_iarg_95_tstrb,
    input [S_AXIS_IARG_95_DMWIDTH-1:0] s_axis_iarg_95_tdata,
    output s_axis_iarg_95_tready,
    output ap_axis_iarg_95_tlast,
    output ap_axis_iarg_95_tvalid,
    output [S_AXIS_IARG_95_WIDTH/8-1:0] ap_axis_iarg_95_tkeep,
    output [S_AXIS_IARG_95_WIDTH/8-1:0] ap_axis_iarg_95_tstrb,
    output [S_AXIS_IARG_95_WIDTH-1:0] ap_axis_iarg_95_tdata,
    input ap_axis_iarg_95_tready,
    //input AXI-Stream pass-through interface 96
    input s_axis_iarg_96_aclk,
    input s_axis_iarg_96_aresetn,
    input s_axis_iarg_96_tlast,
    input s_axis_iarg_96_tvalid,
    input [S_AXIS_IARG_96_DMWIDTH/8-1:0] s_axis_iarg_96_tkeep,
    input [S_AXIS_IARG_96_DMWIDTH/8-1:0] s_axis_iarg_96_tstrb,
    input [S_AXIS_IARG_96_DMWIDTH-1:0] s_axis_iarg_96_tdata,
    output s_axis_iarg_96_tready,
    output ap_axis_iarg_96_tlast,
    output ap_axis_iarg_96_tvalid,
    output [S_AXIS_IARG_96_WIDTH/8-1:0] ap_axis_iarg_96_tkeep,
    output [S_AXIS_IARG_96_WIDTH/8-1:0] ap_axis_iarg_96_tstrb,
    output [S_AXIS_IARG_96_WIDTH-1:0] ap_axis_iarg_96_tdata,
    input ap_axis_iarg_96_tready,
    //input AXI-Stream pass-through interface 97
    input s_axis_iarg_97_aclk,
    input s_axis_iarg_97_aresetn,
    input s_axis_iarg_97_tlast,
    input s_axis_iarg_97_tvalid,
    input [S_AXIS_IARG_97_DMWIDTH/8-1:0] s_axis_iarg_97_tkeep,
    input [S_AXIS_IARG_97_DMWIDTH/8-1:0] s_axis_iarg_97_tstrb,
    input [S_AXIS_IARG_97_DMWIDTH-1:0] s_axis_iarg_97_tdata,
    output s_axis_iarg_97_tready,
    output ap_axis_iarg_97_tlast,
    output ap_axis_iarg_97_tvalid,
    output [S_AXIS_IARG_97_WIDTH/8-1:0] ap_axis_iarg_97_tkeep,
    output [S_AXIS_IARG_97_WIDTH/8-1:0] ap_axis_iarg_97_tstrb,
    output [S_AXIS_IARG_97_WIDTH-1:0] ap_axis_iarg_97_tdata,
    input ap_axis_iarg_97_tready,
    //input AXI-Stream pass-through interface 98
    input s_axis_iarg_98_aclk,
    input s_axis_iarg_98_aresetn,
    input s_axis_iarg_98_tlast,
    input s_axis_iarg_98_tvalid,
    input [S_AXIS_IARG_98_DMWIDTH/8-1:0] s_axis_iarg_98_tkeep,
    input [S_AXIS_IARG_98_DMWIDTH/8-1:0] s_axis_iarg_98_tstrb,
    input [S_AXIS_IARG_98_DMWIDTH-1:0] s_axis_iarg_98_tdata,
    output s_axis_iarg_98_tready,
    output ap_axis_iarg_98_tlast,
    output ap_axis_iarg_98_tvalid,
    output [S_AXIS_IARG_98_WIDTH/8-1:0] ap_axis_iarg_98_tkeep,
    output [S_AXIS_IARG_98_WIDTH/8-1:0] ap_axis_iarg_98_tstrb,
    output [S_AXIS_IARG_98_WIDTH-1:0] ap_axis_iarg_98_tdata,
    input ap_axis_iarg_98_tready,
    //input AXI-Stream pass-through interface 99
    input s_axis_iarg_99_aclk,
    input s_axis_iarg_99_aresetn,
    input s_axis_iarg_99_tlast,
    input s_axis_iarg_99_tvalid,
    input [S_AXIS_IARG_99_DMWIDTH/8-1:0] s_axis_iarg_99_tkeep,
    input [S_AXIS_IARG_99_DMWIDTH/8-1:0] s_axis_iarg_99_tstrb,
    input [S_AXIS_IARG_99_DMWIDTH-1:0] s_axis_iarg_99_tdata,
    output s_axis_iarg_99_tready,
    output ap_axis_iarg_99_tlast,
    output ap_axis_iarg_99_tvalid,
    output [S_AXIS_IARG_99_WIDTH/8-1:0] ap_axis_iarg_99_tkeep,
    output [S_AXIS_IARG_99_WIDTH/8-1:0] ap_axis_iarg_99_tstrb,
    output [S_AXIS_IARG_99_WIDTH-1:0] ap_axis_iarg_99_tdata,
    input ap_axis_iarg_99_tready,
    //input AXI-Stream pass-through interface 100
    input s_axis_iarg_100_aclk,
    input s_axis_iarg_100_aresetn,
    input s_axis_iarg_100_tlast,
    input s_axis_iarg_100_tvalid,
    input [S_AXIS_IARG_100_DMWIDTH/8-1:0] s_axis_iarg_100_tkeep,
    input [S_AXIS_IARG_100_DMWIDTH/8-1:0] s_axis_iarg_100_tstrb,
    input [S_AXIS_IARG_100_DMWIDTH-1:0] s_axis_iarg_100_tdata,
    output s_axis_iarg_100_tready,
    output ap_axis_iarg_100_tlast,
    output ap_axis_iarg_100_tvalid,
    output [S_AXIS_IARG_100_WIDTH/8-1:0] ap_axis_iarg_100_tkeep,
    output [S_AXIS_IARG_100_WIDTH/8-1:0] ap_axis_iarg_100_tstrb,
    output [S_AXIS_IARG_100_WIDTH-1:0] ap_axis_iarg_100_tdata,
    input ap_axis_iarg_100_tready,
    //input AXI-Stream pass-through interface 101
    input s_axis_iarg_101_aclk,
    input s_axis_iarg_101_aresetn,
    input s_axis_iarg_101_tlast,
    input s_axis_iarg_101_tvalid,
    input [S_AXIS_IARG_101_DMWIDTH/8-1:0] s_axis_iarg_101_tkeep,
    input [S_AXIS_IARG_101_DMWIDTH/8-1:0] s_axis_iarg_101_tstrb,
    input [S_AXIS_IARG_101_DMWIDTH-1:0] s_axis_iarg_101_tdata,
    output s_axis_iarg_101_tready,
    output ap_axis_iarg_101_tlast,
    output ap_axis_iarg_101_tvalid,
    output [S_AXIS_IARG_101_WIDTH/8-1:0] ap_axis_iarg_101_tkeep,
    output [S_AXIS_IARG_101_WIDTH/8-1:0] ap_axis_iarg_101_tstrb,
    output [S_AXIS_IARG_101_WIDTH-1:0] ap_axis_iarg_101_tdata,
    input ap_axis_iarg_101_tready,
    //input AXI-Stream pass-through interface 102
    input s_axis_iarg_102_aclk,
    input s_axis_iarg_102_aresetn,
    input s_axis_iarg_102_tlast,
    input s_axis_iarg_102_tvalid,
    input [S_AXIS_IARG_102_DMWIDTH/8-1:0] s_axis_iarg_102_tkeep,
    input [S_AXIS_IARG_102_DMWIDTH/8-1:0] s_axis_iarg_102_tstrb,
    input [S_AXIS_IARG_102_DMWIDTH-1:0] s_axis_iarg_102_tdata,
    output s_axis_iarg_102_tready,
    output ap_axis_iarg_102_tlast,
    output ap_axis_iarg_102_tvalid,
    output [S_AXIS_IARG_102_WIDTH/8-1:0] ap_axis_iarg_102_tkeep,
    output [S_AXIS_IARG_102_WIDTH/8-1:0] ap_axis_iarg_102_tstrb,
    output [S_AXIS_IARG_102_WIDTH-1:0] ap_axis_iarg_102_tdata,
    input ap_axis_iarg_102_tready,
    //input AXI-Stream pass-through interface 103
    input s_axis_iarg_103_aclk,
    input s_axis_iarg_103_aresetn,
    input s_axis_iarg_103_tlast,
    input s_axis_iarg_103_tvalid,
    input [S_AXIS_IARG_103_DMWIDTH/8-1:0] s_axis_iarg_103_tkeep,
    input [S_AXIS_IARG_103_DMWIDTH/8-1:0] s_axis_iarg_103_tstrb,
    input [S_AXIS_IARG_103_DMWIDTH-1:0] s_axis_iarg_103_tdata,
    output s_axis_iarg_103_tready,
    output ap_axis_iarg_103_tlast,
    output ap_axis_iarg_103_tvalid,
    output [S_AXIS_IARG_103_WIDTH/8-1:0] ap_axis_iarg_103_tkeep,
    output [S_AXIS_IARG_103_WIDTH/8-1:0] ap_axis_iarg_103_tstrb,
    output [S_AXIS_IARG_103_WIDTH-1:0] ap_axis_iarg_103_tdata,
    input ap_axis_iarg_103_tready,
    //input AXI-Stream pass-through interface 104
    input s_axis_iarg_104_aclk,
    input s_axis_iarg_104_aresetn,
    input s_axis_iarg_104_tlast,
    input s_axis_iarg_104_tvalid,
    input [S_AXIS_IARG_104_DMWIDTH/8-1:0] s_axis_iarg_104_tkeep,
    input [S_AXIS_IARG_104_DMWIDTH/8-1:0] s_axis_iarg_104_tstrb,
    input [S_AXIS_IARG_104_DMWIDTH-1:0] s_axis_iarg_104_tdata,
    output s_axis_iarg_104_tready,
    output ap_axis_iarg_104_tlast,
    output ap_axis_iarg_104_tvalid,
    output [S_AXIS_IARG_104_WIDTH/8-1:0] ap_axis_iarg_104_tkeep,
    output [S_AXIS_IARG_104_WIDTH/8-1:0] ap_axis_iarg_104_tstrb,
    output [S_AXIS_IARG_104_WIDTH-1:0] ap_axis_iarg_104_tdata,
    input ap_axis_iarg_104_tready,
    //input AXI-Stream pass-through interface 105
    input s_axis_iarg_105_aclk,
    input s_axis_iarg_105_aresetn,
    input s_axis_iarg_105_tlast,
    input s_axis_iarg_105_tvalid,
    input [S_AXIS_IARG_105_DMWIDTH/8-1:0] s_axis_iarg_105_tkeep,
    input [S_AXIS_IARG_105_DMWIDTH/8-1:0] s_axis_iarg_105_tstrb,
    input [S_AXIS_IARG_105_DMWIDTH-1:0] s_axis_iarg_105_tdata,
    output s_axis_iarg_105_tready,
    output ap_axis_iarg_105_tlast,
    output ap_axis_iarg_105_tvalid,
    output [S_AXIS_IARG_105_WIDTH/8-1:0] ap_axis_iarg_105_tkeep,
    output [S_AXIS_IARG_105_WIDTH/8-1:0] ap_axis_iarg_105_tstrb,
    output [S_AXIS_IARG_105_WIDTH-1:0] ap_axis_iarg_105_tdata,
    input ap_axis_iarg_105_tready,
    //input AXI-Stream pass-through interface 106
    input s_axis_iarg_106_aclk,
    input s_axis_iarg_106_aresetn,
    input s_axis_iarg_106_tlast,
    input s_axis_iarg_106_tvalid,
    input [S_AXIS_IARG_106_DMWIDTH/8-1:0] s_axis_iarg_106_tkeep,
    input [S_AXIS_IARG_106_DMWIDTH/8-1:0] s_axis_iarg_106_tstrb,
    input [S_AXIS_IARG_106_DMWIDTH-1:0] s_axis_iarg_106_tdata,
    output s_axis_iarg_106_tready,
    output ap_axis_iarg_106_tlast,
    output ap_axis_iarg_106_tvalid,
    output [S_AXIS_IARG_106_WIDTH/8-1:0] ap_axis_iarg_106_tkeep,
    output [S_AXIS_IARG_106_WIDTH/8-1:0] ap_axis_iarg_106_tstrb,
    output [S_AXIS_IARG_106_WIDTH-1:0] ap_axis_iarg_106_tdata,
    input ap_axis_iarg_106_tready,
    //input AXI-Stream pass-through interface 107
    input s_axis_iarg_107_aclk,
    input s_axis_iarg_107_aresetn,
    input s_axis_iarg_107_tlast,
    input s_axis_iarg_107_tvalid,
    input [S_AXIS_IARG_107_DMWIDTH/8-1:0] s_axis_iarg_107_tkeep,
    input [S_AXIS_IARG_107_DMWIDTH/8-1:0] s_axis_iarg_107_tstrb,
    input [S_AXIS_IARG_107_DMWIDTH-1:0] s_axis_iarg_107_tdata,
    output s_axis_iarg_107_tready,
    output ap_axis_iarg_107_tlast,
    output ap_axis_iarg_107_tvalid,
    output [S_AXIS_IARG_107_WIDTH/8-1:0] ap_axis_iarg_107_tkeep,
    output [S_AXIS_IARG_107_WIDTH/8-1:0] ap_axis_iarg_107_tstrb,
    output [S_AXIS_IARG_107_WIDTH-1:0] ap_axis_iarg_107_tdata,
    input ap_axis_iarg_107_tready,
    //input AXI-Stream pass-through interface 108
    input s_axis_iarg_108_aclk,
    input s_axis_iarg_108_aresetn,
    input s_axis_iarg_108_tlast,
    input s_axis_iarg_108_tvalid,
    input [S_AXIS_IARG_108_DMWIDTH/8-1:0] s_axis_iarg_108_tkeep,
    input [S_AXIS_IARG_108_DMWIDTH/8-1:0] s_axis_iarg_108_tstrb,
    input [S_AXIS_IARG_108_DMWIDTH-1:0] s_axis_iarg_108_tdata,
    output s_axis_iarg_108_tready,
    output ap_axis_iarg_108_tlast,
    output ap_axis_iarg_108_tvalid,
    output [S_AXIS_IARG_108_WIDTH/8-1:0] ap_axis_iarg_108_tkeep,
    output [S_AXIS_IARG_108_WIDTH/8-1:0] ap_axis_iarg_108_tstrb,
    output [S_AXIS_IARG_108_WIDTH-1:0] ap_axis_iarg_108_tdata,
    input ap_axis_iarg_108_tready,
    //input AXI-Stream pass-through interface 109
    input s_axis_iarg_109_aclk,
    input s_axis_iarg_109_aresetn,
    input s_axis_iarg_109_tlast,
    input s_axis_iarg_109_tvalid,
    input [S_AXIS_IARG_109_DMWIDTH/8-1:0] s_axis_iarg_109_tkeep,
    input [S_AXIS_IARG_109_DMWIDTH/8-1:0] s_axis_iarg_109_tstrb,
    input [S_AXIS_IARG_109_DMWIDTH-1:0] s_axis_iarg_109_tdata,
    output s_axis_iarg_109_tready,
    output ap_axis_iarg_109_tlast,
    output ap_axis_iarg_109_tvalid,
    output [S_AXIS_IARG_109_WIDTH/8-1:0] ap_axis_iarg_109_tkeep,
    output [S_AXIS_IARG_109_WIDTH/8-1:0] ap_axis_iarg_109_tstrb,
    output [S_AXIS_IARG_109_WIDTH-1:0] ap_axis_iarg_109_tdata,
    input ap_axis_iarg_109_tready,
    //input AXI-Stream pass-through interface 110
    input s_axis_iarg_110_aclk,
    input s_axis_iarg_110_aresetn,
    input s_axis_iarg_110_tlast,
    input s_axis_iarg_110_tvalid,
    input [S_AXIS_IARG_110_DMWIDTH/8-1:0] s_axis_iarg_110_tkeep,
    input [S_AXIS_IARG_110_DMWIDTH/8-1:0] s_axis_iarg_110_tstrb,
    input [S_AXIS_IARG_110_DMWIDTH-1:0] s_axis_iarg_110_tdata,
    output s_axis_iarg_110_tready,
    output ap_axis_iarg_110_tlast,
    output ap_axis_iarg_110_tvalid,
    output [S_AXIS_IARG_110_WIDTH/8-1:0] ap_axis_iarg_110_tkeep,
    output [S_AXIS_IARG_110_WIDTH/8-1:0] ap_axis_iarg_110_tstrb,
    output [S_AXIS_IARG_110_WIDTH-1:0] ap_axis_iarg_110_tdata,
    input ap_axis_iarg_110_tready,
    //input AXI-Stream pass-through interface 111
    input s_axis_iarg_111_aclk,
    input s_axis_iarg_111_aresetn,
    input s_axis_iarg_111_tlast,
    input s_axis_iarg_111_tvalid,
    input [S_AXIS_IARG_111_DMWIDTH/8-1:0] s_axis_iarg_111_tkeep,
    input [S_AXIS_IARG_111_DMWIDTH/8-1:0] s_axis_iarg_111_tstrb,
    input [S_AXIS_IARG_111_DMWIDTH-1:0] s_axis_iarg_111_tdata,
    output s_axis_iarg_111_tready,
    output ap_axis_iarg_111_tlast,
    output ap_axis_iarg_111_tvalid,
    output [S_AXIS_IARG_111_WIDTH/8-1:0] ap_axis_iarg_111_tkeep,
    output [S_AXIS_IARG_111_WIDTH/8-1:0] ap_axis_iarg_111_tstrb,
    output [S_AXIS_IARG_111_WIDTH-1:0] ap_axis_iarg_111_tdata,
    input ap_axis_iarg_111_tready,
    //input AXI-Stream pass-through interface 112
    input s_axis_iarg_112_aclk,
    input s_axis_iarg_112_aresetn,
    input s_axis_iarg_112_tlast,
    input s_axis_iarg_112_tvalid,
    input [S_AXIS_IARG_112_DMWIDTH/8-1:0] s_axis_iarg_112_tkeep,
    input [S_AXIS_IARG_112_DMWIDTH/8-1:0] s_axis_iarg_112_tstrb,
    input [S_AXIS_IARG_112_DMWIDTH-1:0] s_axis_iarg_112_tdata,
    output s_axis_iarg_112_tready,
    output ap_axis_iarg_112_tlast,
    output ap_axis_iarg_112_tvalid,
    output [S_AXIS_IARG_112_WIDTH/8-1:0] ap_axis_iarg_112_tkeep,
    output [S_AXIS_IARG_112_WIDTH/8-1:0] ap_axis_iarg_112_tstrb,
    output [S_AXIS_IARG_112_WIDTH-1:0] ap_axis_iarg_112_tdata,
    input ap_axis_iarg_112_tready,
    //input AXI-Stream pass-through interface 113
    input s_axis_iarg_113_aclk,
    input s_axis_iarg_113_aresetn,
    input s_axis_iarg_113_tlast,
    input s_axis_iarg_113_tvalid,
    input [S_AXIS_IARG_113_DMWIDTH/8-1:0] s_axis_iarg_113_tkeep,
    input [S_AXIS_IARG_113_DMWIDTH/8-1:0] s_axis_iarg_113_tstrb,
    input [S_AXIS_IARG_113_DMWIDTH-1:0] s_axis_iarg_113_tdata,
    output s_axis_iarg_113_tready,
    output ap_axis_iarg_113_tlast,
    output ap_axis_iarg_113_tvalid,
    output [S_AXIS_IARG_113_WIDTH/8-1:0] ap_axis_iarg_113_tkeep,
    output [S_AXIS_IARG_113_WIDTH/8-1:0] ap_axis_iarg_113_tstrb,
    output [S_AXIS_IARG_113_WIDTH-1:0] ap_axis_iarg_113_tdata,
    input ap_axis_iarg_113_tready,
    //input AXI-Stream pass-through interface 114
    input s_axis_iarg_114_aclk,
    input s_axis_iarg_114_aresetn,
    input s_axis_iarg_114_tlast,
    input s_axis_iarg_114_tvalid,
    input [S_AXIS_IARG_114_DMWIDTH/8-1:0] s_axis_iarg_114_tkeep,
    input [S_AXIS_IARG_114_DMWIDTH/8-1:0] s_axis_iarg_114_tstrb,
    input [S_AXIS_IARG_114_DMWIDTH-1:0] s_axis_iarg_114_tdata,
    output s_axis_iarg_114_tready,
    output ap_axis_iarg_114_tlast,
    output ap_axis_iarg_114_tvalid,
    output [S_AXIS_IARG_114_WIDTH/8-1:0] ap_axis_iarg_114_tkeep,
    output [S_AXIS_IARG_114_WIDTH/8-1:0] ap_axis_iarg_114_tstrb,
    output [S_AXIS_IARG_114_WIDTH-1:0] ap_axis_iarg_114_tdata,
    input ap_axis_iarg_114_tready,
    //input AXI-Stream pass-through interface 115
    input s_axis_iarg_115_aclk,
    input s_axis_iarg_115_aresetn,
    input s_axis_iarg_115_tlast,
    input s_axis_iarg_115_tvalid,
    input [S_AXIS_IARG_115_DMWIDTH/8-1:0] s_axis_iarg_115_tkeep,
    input [S_AXIS_IARG_115_DMWIDTH/8-1:0] s_axis_iarg_115_tstrb,
    input [S_AXIS_IARG_115_DMWIDTH-1:0] s_axis_iarg_115_tdata,
    output s_axis_iarg_115_tready,
    output ap_axis_iarg_115_tlast,
    output ap_axis_iarg_115_tvalid,
    output [S_AXIS_IARG_115_WIDTH/8-1:0] ap_axis_iarg_115_tkeep,
    output [S_AXIS_IARG_115_WIDTH/8-1:0] ap_axis_iarg_115_tstrb,
    output [S_AXIS_IARG_115_WIDTH-1:0] ap_axis_iarg_115_tdata,
    input ap_axis_iarg_115_tready,
    //input AXI-Stream pass-through interface 116
    input s_axis_iarg_116_aclk,
    input s_axis_iarg_116_aresetn,
    input s_axis_iarg_116_tlast,
    input s_axis_iarg_116_tvalid,
    input [S_AXIS_IARG_116_DMWIDTH/8-1:0] s_axis_iarg_116_tkeep,
    input [S_AXIS_IARG_116_DMWIDTH/8-1:0] s_axis_iarg_116_tstrb,
    input [S_AXIS_IARG_116_DMWIDTH-1:0] s_axis_iarg_116_tdata,
    output s_axis_iarg_116_tready,
    output ap_axis_iarg_116_tlast,
    output ap_axis_iarg_116_tvalid,
    output [S_AXIS_IARG_116_WIDTH/8-1:0] ap_axis_iarg_116_tkeep,
    output [S_AXIS_IARG_116_WIDTH/8-1:0] ap_axis_iarg_116_tstrb,
    output [S_AXIS_IARG_116_WIDTH-1:0] ap_axis_iarg_116_tdata,
    input ap_axis_iarg_116_tready,
    //input AXI-Stream pass-through interface 117
    input s_axis_iarg_117_aclk,
    input s_axis_iarg_117_aresetn,
    input s_axis_iarg_117_tlast,
    input s_axis_iarg_117_tvalid,
    input [S_AXIS_IARG_117_DMWIDTH/8-1:0] s_axis_iarg_117_tkeep,
    input [S_AXIS_IARG_117_DMWIDTH/8-1:0] s_axis_iarg_117_tstrb,
    input [S_AXIS_IARG_117_DMWIDTH-1:0] s_axis_iarg_117_tdata,
    output s_axis_iarg_117_tready,
    output ap_axis_iarg_117_tlast,
    output ap_axis_iarg_117_tvalid,
    output [S_AXIS_IARG_117_WIDTH/8-1:0] ap_axis_iarg_117_tkeep,
    output [S_AXIS_IARG_117_WIDTH/8-1:0] ap_axis_iarg_117_tstrb,
    output [S_AXIS_IARG_117_WIDTH-1:0] ap_axis_iarg_117_tdata,
    input ap_axis_iarg_117_tready,
    //input AXI-Stream pass-through interface 118
    input s_axis_iarg_118_aclk,
    input s_axis_iarg_118_aresetn,
    input s_axis_iarg_118_tlast,
    input s_axis_iarg_118_tvalid,
    input [S_AXIS_IARG_118_DMWIDTH/8-1:0] s_axis_iarg_118_tkeep,
    input [S_AXIS_IARG_118_DMWIDTH/8-1:0] s_axis_iarg_118_tstrb,
    input [S_AXIS_IARG_118_DMWIDTH-1:0] s_axis_iarg_118_tdata,
    output s_axis_iarg_118_tready,
    output ap_axis_iarg_118_tlast,
    output ap_axis_iarg_118_tvalid,
    output [S_AXIS_IARG_118_WIDTH/8-1:0] ap_axis_iarg_118_tkeep,
    output [S_AXIS_IARG_118_WIDTH/8-1:0] ap_axis_iarg_118_tstrb,
    output [S_AXIS_IARG_118_WIDTH-1:0] ap_axis_iarg_118_tdata,
    input ap_axis_iarg_118_tready,
    //input AXI-Stream pass-through interface 119
    input s_axis_iarg_119_aclk,
    input s_axis_iarg_119_aresetn,
    input s_axis_iarg_119_tlast,
    input s_axis_iarg_119_tvalid,
    input [S_AXIS_IARG_119_DMWIDTH/8-1:0] s_axis_iarg_119_tkeep,
    input [S_AXIS_IARG_119_DMWIDTH/8-1:0] s_axis_iarg_119_tstrb,
    input [S_AXIS_IARG_119_DMWIDTH-1:0] s_axis_iarg_119_tdata,
    output s_axis_iarg_119_tready,
    output ap_axis_iarg_119_tlast,
    output ap_axis_iarg_119_tvalid,
    output [S_AXIS_IARG_119_WIDTH/8-1:0] ap_axis_iarg_119_tkeep,
    output [S_AXIS_IARG_119_WIDTH/8-1:0] ap_axis_iarg_119_tstrb,
    output [S_AXIS_IARG_119_WIDTH-1:0] ap_axis_iarg_119_tdata,
    input ap_axis_iarg_119_tready,
    //input AXI-Stream pass-through interface 120
    input s_axis_iarg_120_aclk,
    input s_axis_iarg_120_aresetn,
    input s_axis_iarg_120_tlast,
    input s_axis_iarg_120_tvalid,
    input [S_AXIS_IARG_120_DMWIDTH/8-1:0] s_axis_iarg_120_tkeep,
    input [S_AXIS_IARG_120_DMWIDTH/8-1:0] s_axis_iarg_120_tstrb,
    input [S_AXIS_IARG_120_DMWIDTH-1:0] s_axis_iarg_120_tdata,
    output s_axis_iarg_120_tready,
    output ap_axis_iarg_120_tlast,
    output ap_axis_iarg_120_tvalid,
    output [S_AXIS_IARG_120_WIDTH/8-1:0] ap_axis_iarg_120_tkeep,
    output [S_AXIS_IARG_120_WIDTH/8-1:0] ap_axis_iarg_120_tstrb,
    output [S_AXIS_IARG_120_WIDTH-1:0] ap_axis_iarg_120_tdata,
    input ap_axis_iarg_120_tready,
    //input AXI-Stream pass-through interface 121
    input s_axis_iarg_121_aclk,
    input s_axis_iarg_121_aresetn,
    input s_axis_iarg_121_tlast,
    input s_axis_iarg_121_tvalid,
    input [S_AXIS_IARG_121_DMWIDTH/8-1:0] s_axis_iarg_121_tkeep,
    input [S_AXIS_IARG_121_DMWIDTH/8-1:0] s_axis_iarg_121_tstrb,
    input [S_AXIS_IARG_121_DMWIDTH-1:0] s_axis_iarg_121_tdata,
    output s_axis_iarg_121_tready,
    output ap_axis_iarg_121_tlast,
    output ap_axis_iarg_121_tvalid,
    output [S_AXIS_IARG_121_WIDTH/8-1:0] ap_axis_iarg_121_tkeep,
    output [S_AXIS_IARG_121_WIDTH/8-1:0] ap_axis_iarg_121_tstrb,
    output [S_AXIS_IARG_121_WIDTH-1:0] ap_axis_iarg_121_tdata,
    input ap_axis_iarg_121_tready,
    //input AXI-Stream pass-through interface 122
    input s_axis_iarg_122_aclk,
    input s_axis_iarg_122_aresetn,
    input s_axis_iarg_122_tlast,
    input s_axis_iarg_122_tvalid,
    input [S_AXIS_IARG_122_DMWIDTH/8-1:0] s_axis_iarg_122_tkeep,
    input [S_AXIS_IARG_122_DMWIDTH/8-1:0] s_axis_iarg_122_tstrb,
    input [S_AXIS_IARG_122_DMWIDTH-1:0] s_axis_iarg_122_tdata,
    output s_axis_iarg_122_tready,
    output ap_axis_iarg_122_tlast,
    output ap_axis_iarg_122_tvalid,
    output [S_AXIS_IARG_122_WIDTH/8-1:0] ap_axis_iarg_122_tkeep,
    output [S_AXIS_IARG_122_WIDTH/8-1:0] ap_axis_iarg_122_tstrb,
    output [S_AXIS_IARG_122_WIDTH-1:0] ap_axis_iarg_122_tdata,
    input ap_axis_iarg_122_tready,
    //input AXI-Stream pass-through interface 123
    input s_axis_iarg_123_aclk,
    input s_axis_iarg_123_aresetn,
    input s_axis_iarg_123_tlast,
    input s_axis_iarg_123_tvalid,
    input [S_AXIS_IARG_123_DMWIDTH/8-1:0] s_axis_iarg_123_tkeep,
    input [S_AXIS_IARG_123_DMWIDTH/8-1:0] s_axis_iarg_123_tstrb,
    input [S_AXIS_IARG_123_DMWIDTH-1:0] s_axis_iarg_123_tdata,
    output s_axis_iarg_123_tready,
    output ap_axis_iarg_123_tlast,
    output ap_axis_iarg_123_tvalid,
    output [S_AXIS_IARG_123_WIDTH/8-1:0] ap_axis_iarg_123_tkeep,
    output [S_AXIS_IARG_123_WIDTH/8-1:0] ap_axis_iarg_123_tstrb,
    output [S_AXIS_IARG_123_WIDTH-1:0] ap_axis_iarg_123_tdata,
    input ap_axis_iarg_123_tready,
    //input AXI-Stream pass-through interface 124
    input s_axis_iarg_124_aclk,
    input s_axis_iarg_124_aresetn,
    input s_axis_iarg_124_tlast,
    input s_axis_iarg_124_tvalid,
    input [S_AXIS_IARG_124_DMWIDTH/8-1:0] s_axis_iarg_124_tkeep,
    input [S_AXIS_IARG_124_DMWIDTH/8-1:0] s_axis_iarg_124_tstrb,
    input [S_AXIS_IARG_124_DMWIDTH-1:0] s_axis_iarg_124_tdata,
    output s_axis_iarg_124_tready,
    output ap_axis_iarg_124_tlast,
    output ap_axis_iarg_124_tvalid,
    output [S_AXIS_IARG_124_WIDTH/8-1:0] ap_axis_iarg_124_tkeep,
    output [S_AXIS_IARG_124_WIDTH/8-1:0] ap_axis_iarg_124_tstrb,
    output [S_AXIS_IARG_124_WIDTH-1:0] ap_axis_iarg_124_tdata,
    input ap_axis_iarg_124_tready,
    //input AXI-Stream pass-through interface 125
    input s_axis_iarg_125_aclk,
    input s_axis_iarg_125_aresetn,
    input s_axis_iarg_125_tlast,
    input s_axis_iarg_125_tvalid,
    input [S_AXIS_IARG_125_DMWIDTH/8-1:0] s_axis_iarg_125_tkeep,
    input [S_AXIS_IARG_125_DMWIDTH/8-1:0] s_axis_iarg_125_tstrb,
    input [S_AXIS_IARG_125_DMWIDTH-1:0] s_axis_iarg_125_tdata,
    output s_axis_iarg_125_tready,
    output ap_axis_iarg_125_tlast,
    output ap_axis_iarg_125_tvalid,
    output [S_AXIS_IARG_125_WIDTH/8-1:0] ap_axis_iarg_125_tkeep,
    output [S_AXIS_IARG_125_WIDTH/8-1:0] ap_axis_iarg_125_tstrb,
    output [S_AXIS_IARG_125_WIDTH-1:0] ap_axis_iarg_125_tdata,
    input ap_axis_iarg_125_tready,
    //input AXI-Stream pass-through interface 126
    input s_axis_iarg_126_aclk,
    input s_axis_iarg_126_aresetn,
    input s_axis_iarg_126_tlast,
    input s_axis_iarg_126_tvalid,
    input [S_AXIS_IARG_126_DMWIDTH/8-1:0] s_axis_iarg_126_tkeep,
    input [S_AXIS_IARG_126_DMWIDTH/8-1:0] s_axis_iarg_126_tstrb,
    input [S_AXIS_IARG_126_DMWIDTH-1:0] s_axis_iarg_126_tdata,
    output s_axis_iarg_126_tready,
    output ap_axis_iarg_126_tlast,
    output ap_axis_iarg_126_tvalid,
    output [S_AXIS_IARG_126_WIDTH/8-1:0] ap_axis_iarg_126_tkeep,
    output [S_AXIS_IARG_126_WIDTH/8-1:0] ap_axis_iarg_126_tstrb,
    output [S_AXIS_IARG_126_WIDTH-1:0] ap_axis_iarg_126_tdata,
    input ap_axis_iarg_126_tready,
    //input AXI-Stream pass-through interface 127
    input s_axis_iarg_127_aclk,
    input s_axis_iarg_127_aresetn,
    input s_axis_iarg_127_tlast,
    input s_axis_iarg_127_tvalid,
    input [S_AXIS_IARG_127_DMWIDTH/8-1:0] s_axis_iarg_127_tkeep,
    input [S_AXIS_IARG_127_DMWIDTH/8-1:0] s_axis_iarg_127_tstrb,
    input [S_AXIS_IARG_127_DMWIDTH-1:0] s_axis_iarg_127_tdata,
    output s_axis_iarg_127_tready,
    output ap_axis_iarg_127_tlast,
    output ap_axis_iarg_127_tvalid,
    output [S_AXIS_IARG_127_WIDTH/8-1:0] ap_axis_iarg_127_tkeep,
    output [S_AXIS_IARG_127_WIDTH/8-1:0] ap_axis_iarg_127_tstrb,
    output [S_AXIS_IARG_127_WIDTH-1:0] ap_axis_iarg_127_tdata,
    input ap_axis_iarg_127_tready
    );
    

    localparam C_MAX_INPUT_AXISs = 128;
    localparam C_MAX_BIT_WIDTH = 1024;
    localparam [(C_MAX_INPUT_AXISs*32)-1:0] C_INAXIS_BIT_ARRAY = {S_AXIS_IARG_127_WIDTH,S_AXIS_IARG_126_WIDTH,S_AXIS_IARG_125_WIDTH,S_AXIS_IARG_124_WIDTH,S_AXIS_IARG_123_WIDTH,S_AXIS_IARG_122_WIDTH,S_AXIS_IARG_121_WIDTH,S_AXIS_IARG_120_WIDTH,S_AXIS_IARG_119_WIDTH,S_AXIS_IARG_118_WIDTH,S_AXIS_IARG_117_WIDTH,S_AXIS_IARG_116_WIDTH,S_AXIS_IARG_115_WIDTH,S_AXIS_IARG_114_WIDTH,S_AXIS_IARG_113_WIDTH,S_AXIS_IARG_112_WIDTH,S_AXIS_IARG_111_WIDTH,S_AXIS_IARG_110_WIDTH,S_AXIS_IARG_109_WIDTH,S_AXIS_IARG_108_WIDTH,S_AXIS_IARG_107_WIDTH,S_AXIS_IARG_106_WIDTH,S_AXIS_IARG_105_WIDTH,S_AXIS_IARG_104_WIDTH,S_AXIS_IARG_103_WIDTH,S_AXIS_IARG_102_WIDTH,S_AXIS_IARG_101_WIDTH,S_AXIS_IARG_100_WIDTH,S_AXIS_IARG_99_WIDTH,S_AXIS_IARG_98_WIDTH,S_AXIS_IARG_97_WIDTH,S_AXIS_IARG_96_WIDTH,S_AXIS_IARG_95_WIDTH,S_AXIS_IARG_94_WIDTH,S_AXIS_IARG_93_WIDTH,S_AXIS_IARG_92_WIDTH,S_AXIS_IARG_91_WIDTH,S_AXIS_IARG_90_WIDTH,S_AXIS_IARG_89_WIDTH,S_AXIS_IARG_88_WIDTH,S_AXIS_IARG_87_WIDTH,S_AXIS_IARG_86_WIDTH,S_AXIS_IARG_85_WIDTH,S_AXIS_IARG_84_WIDTH,S_AXIS_IARG_83_WIDTH,S_AXIS_IARG_82_WIDTH,S_AXIS_IARG_81_WIDTH,S_AXIS_IARG_80_WIDTH,S_AXIS_IARG_79_WIDTH,S_AXIS_IARG_78_WIDTH,S_AXIS_IARG_77_WIDTH,S_AXIS_IARG_76_WIDTH,S_AXIS_IARG_75_WIDTH,S_AXIS_IARG_74_WIDTH,S_AXIS_IARG_73_WIDTH,S_AXIS_IARG_72_WIDTH,S_AXIS_IARG_71_WIDTH,S_AXIS_IARG_70_WIDTH,S_AXIS_IARG_69_WIDTH,S_AXIS_IARG_68_WIDTH,S_AXIS_IARG_67_WIDTH,S_AXIS_IARG_66_WIDTH,S_AXIS_IARG_65_WIDTH,S_AXIS_IARG_64_WIDTH,S_AXIS_IARG_63_WIDTH,S_AXIS_IARG_62_WIDTH,S_AXIS_IARG_61_WIDTH,S_AXIS_IARG_60_WIDTH,S_AXIS_IARG_59_WIDTH,S_AXIS_IARG_58_WIDTH,S_AXIS_IARG_57_WIDTH,S_AXIS_IARG_56_WIDTH,S_AXIS_IARG_55_WIDTH,S_AXIS_IARG_54_WIDTH,S_AXIS_IARG_53_WIDTH,S_AXIS_IARG_52_WIDTH,S_AXIS_IARG_51_WIDTH,S_AXIS_IARG_50_WIDTH,S_AXIS_IARG_49_WIDTH,S_AXIS_IARG_48_WIDTH,S_AXIS_IARG_47_WIDTH,S_AXIS_IARG_46_WIDTH,S_AXIS_IARG_45_WIDTH,S_AXIS_IARG_44_WIDTH,S_AXIS_IARG_43_WIDTH,S_AXIS_IARG_42_WIDTH,S_AXIS_IARG_41_WIDTH,S_AXIS_IARG_40_WIDTH,S_AXIS_IARG_39_WIDTH,S_AXIS_IARG_38_WIDTH,S_AXIS_IARG_37_WIDTH,S_AXIS_IARG_36_WIDTH,S_AXIS_IARG_35_WIDTH,S_AXIS_IARG_34_WIDTH,S_AXIS_IARG_33_WIDTH,S_AXIS_IARG_32_WIDTH,S_AXIS_IARG_31_WIDTH,S_AXIS_IARG_30_WIDTH,S_AXIS_IARG_29_WIDTH,S_AXIS_IARG_28_WIDTH,S_AXIS_IARG_27_WIDTH,S_AXIS_IARG_26_WIDTH,S_AXIS_IARG_25_WIDTH,S_AXIS_IARG_24_WIDTH,S_AXIS_IARG_23_WIDTH,S_AXIS_IARG_22_WIDTH,S_AXIS_IARG_21_WIDTH,S_AXIS_IARG_20_WIDTH,S_AXIS_IARG_19_WIDTH,S_AXIS_IARG_18_WIDTH,S_AXIS_IARG_17_WIDTH,S_AXIS_IARG_16_WIDTH,S_AXIS_IARG_15_WIDTH,S_AXIS_IARG_14_WIDTH,S_AXIS_IARG_13_WIDTH,S_AXIS_IARG_12_WIDTH,S_AXIS_IARG_11_WIDTH,S_AXIS_IARG_10_WIDTH,S_AXIS_IARG_9_WIDTH,S_AXIS_IARG_8_WIDTH,S_AXIS_IARG_7_WIDTH,S_AXIS_IARG_6_WIDTH,S_AXIS_IARG_5_WIDTH,S_AXIS_IARG_4_WIDTH,S_AXIS_IARG_3_WIDTH,S_AXIS_IARG_2_WIDTH,S_AXIS_IARG_1_WIDTH,S_AXIS_IARG_0_WIDTH};
    localparam [(C_MAX_INPUT_AXISs*32)-1:0] C_DEPTH_BIT_ARRAY = {S_AXIS_IARG_127_DEPTH,S_AXIS_IARG_126_DEPTH,S_AXIS_IARG_125_DEPTH,S_AXIS_IARG_124_DEPTH,S_AXIS_IARG_123_DEPTH,S_AXIS_IARG_122_DEPTH,S_AXIS_IARG_121_DEPTH,S_AXIS_IARG_120_DEPTH,S_AXIS_IARG_119_DEPTH,S_AXIS_IARG_118_DEPTH,S_AXIS_IARG_117_DEPTH,S_AXIS_IARG_116_DEPTH,S_AXIS_IARG_115_DEPTH,S_AXIS_IARG_114_DEPTH,S_AXIS_IARG_113_DEPTH,S_AXIS_IARG_112_DEPTH,S_AXIS_IARG_111_DEPTH,S_AXIS_IARG_110_DEPTH,S_AXIS_IARG_109_DEPTH,S_AXIS_IARG_108_DEPTH,S_AXIS_IARG_107_DEPTH,S_AXIS_IARG_106_DEPTH,S_AXIS_IARG_105_DEPTH,S_AXIS_IARG_104_DEPTH,S_AXIS_IARG_103_DEPTH,S_AXIS_IARG_102_DEPTH,S_AXIS_IARG_101_DEPTH,S_AXIS_IARG_100_DEPTH,S_AXIS_IARG_99_DEPTH,S_AXIS_IARG_98_DEPTH,S_AXIS_IARG_97_DEPTH,S_AXIS_IARG_96_DEPTH,S_AXIS_IARG_95_DEPTH,S_AXIS_IARG_94_DEPTH,S_AXIS_IARG_93_DEPTH,S_AXIS_IARG_92_DEPTH,S_AXIS_IARG_91_DEPTH,S_AXIS_IARG_90_DEPTH,S_AXIS_IARG_89_DEPTH,S_AXIS_IARG_88_DEPTH,S_AXIS_IARG_87_DEPTH,S_AXIS_IARG_86_DEPTH,S_AXIS_IARG_85_DEPTH,S_AXIS_IARG_84_DEPTH,S_AXIS_IARG_83_DEPTH,S_AXIS_IARG_82_DEPTH,S_AXIS_IARG_81_DEPTH,S_AXIS_IARG_80_DEPTH,S_AXIS_IARG_79_DEPTH,S_AXIS_IARG_78_DEPTH,S_AXIS_IARG_77_DEPTH,S_AXIS_IARG_76_DEPTH,S_AXIS_IARG_75_DEPTH,S_AXIS_IARG_74_DEPTH,S_AXIS_IARG_73_DEPTH,S_AXIS_IARG_72_DEPTH,S_AXIS_IARG_71_DEPTH,S_AXIS_IARG_70_DEPTH,S_AXIS_IARG_69_DEPTH,S_AXIS_IARG_68_DEPTH,S_AXIS_IARG_67_DEPTH,S_AXIS_IARG_66_DEPTH,S_AXIS_IARG_65_DEPTH,S_AXIS_IARG_64_DEPTH,S_AXIS_IARG_63_DEPTH,S_AXIS_IARG_62_DEPTH,S_AXIS_IARG_61_DEPTH,S_AXIS_IARG_60_DEPTH,S_AXIS_IARG_59_DEPTH,S_AXIS_IARG_58_DEPTH,S_AXIS_IARG_57_DEPTH,S_AXIS_IARG_56_DEPTH,S_AXIS_IARG_55_DEPTH,S_AXIS_IARG_54_DEPTH,S_AXIS_IARG_53_DEPTH,S_AXIS_IARG_52_DEPTH,S_AXIS_IARG_51_DEPTH,S_AXIS_IARG_50_DEPTH,S_AXIS_IARG_49_DEPTH,S_AXIS_IARG_48_DEPTH,S_AXIS_IARG_47_DEPTH,S_AXIS_IARG_46_DEPTH,S_AXIS_IARG_45_DEPTH,S_AXIS_IARG_44_DEPTH,S_AXIS_IARG_43_DEPTH,S_AXIS_IARG_42_DEPTH,S_AXIS_IARG_41_DEPTH,S_AXIS_IARG_40_DEPTH,S_AXIS_IARG_39_DEPTH,S_AXIS_IARG_38_DEPTH,S_AXIS_IARG_37_DEPTH,S_AXIS_IARG_36_DEPTH,S_AXIS_IARG_35_DEPTH,S_AXIS_IARG_34_DEPTH,S_AXIS_IARG_33_DEPTH,S_AXIS_IARG_32_DEPTH,S_AXIS_IARG_31_DEPTH,S_AXIS_IARG_30_DEPTH,S_AXIS_IARG_29_DEPTH,S_AXIS_IARG_28_DEPTH,S_AXIS_IARG_27_DEPTH,S_AXIS_IARG_26_DEPTH,S_AXIS_IARG_25_DEPTH,S_AXIS_IARG_24_DEPTH,S_AXIS_IARG_23_DEPTH,S_AXIS_IARG_22_DEPTH,S_AXIS_IARG_21_DEPTH,S_AXIS_IARG_20_DEPTH,S_AXIS_IARG_19_DEPTH,S_AXIS_IARG_18_DEPTH,S_AXIS_IARG_17_DEPTH,S_AXIS_IARG_16_DEPTH,S_AXIS_IARG_15_DEPTH,S_AXIS_IARG_14_DEPTH,S_AXIS_IARG_13_DEPTH,S_AXIS_IARG_12_DEPTH,S_AXIS_IARG_11_DEPTH,S_AXIS_IARG_10_DEPTH,S_AXIS_IARG_9_DEPTH,S_AXIS_IARG_8_DEPTH,S_AXIS_IARG_7_DEPTH,S_AXIS_IARG_6_DEPTH,S_AXIS_IARG_5_DEPTH,S_AXIS_IARG_4_DEPTH,S_AXIS_IARG_3_DEPTH,S_AXIS_IARG_2_DEPTH,S_AXIS_IARG_1_DEPTH,S_AXIS_IARG_0_DEPTH};
    localparam [(C_MAX_INPUT_AXISs*32)-1:0] C_DMWIDTH_BIT_ARRAY = {S_AXIS_IARG_127_DMWIDTH,S_AXIS_IARG_126_DMWIDTH,S_AXIS_IARG_125_DMWIDTH,S_AXIS_IARG_124_DMWIDTH,S_AXIS_IARG_123_DMWIDTH,S_AXIS_IARG_122_DMWIDTH,S_AXIS_IARG_121_DMWIDTH,S_AXIS_IARG_120_DMWIDTH,S_AXIS_IARG_119_DMWIDTH,S_AXIS_IARG_118_DMWIDTH,S_AXIS_IARG_117_DMWIDTH,S_AXIS_IARG_116_DMWIDTH,S_AXIS_IARG_115_DMWIDTH,S_AXIS_IARG_114_DMWIDTH,S_AXIS_IARG_113_DMWIDTH,S_AXIS_IARG_112_DMWIDTH,S_AXIS_IARG_111_DMWIDTH,S_AXIS_IARG_110_DMWIDTH,S_AXIS_IARG_109_DMWIDTH,S_AXIS_IARG_108_DMWIDTH,S_AXIS_IARG_107_DMWIDTH,S_AXIS_IARG_106_DMWIDTH,S_AXIS_IARG_105_DMWIDTH,S_AXIS_IARG_104_DMWIDTH,S_AXIS_IARG_103_DMWIDTH,S_AXIS_IARG_102_DMWIDTH,S_AXIS_IARG_101_DMWIDTH,S_AXIS_IARG_100_DMWIDTH,S_AXIS_IARG_99_DMWIDTH,S_AXIS_IARG_98_DMWIDTH,S_AXIS_IARG_97_DMWIDTH,S_AXIS_IARG_96_DMWIDTH,S_AXIS_IARG_95_DMWIDTH,S_AXIS_IARG_94_DMWIDTH,S_AXIS_IARG_93_DMWIDTH,S_AXIS_IARG_92_DMWIDTH,S_AXIS_IARG_91_DMWIDTH,S_AXIS_IARG_90_DMWIDTH,S_AXIS_IARG_89_DMWIDTH,S_AXIS_IARG_88_DMWIDTH,S_AXIS_IARG_87_DMWIDTH,S_AXIS_IARG_86_DMWIDTH,S_AXIS_IARG_85_DMWIDTH,S_AXIS_IARG_84_DMWIDTH,S_AXIS_IARG_83_DMWIDTH,S_AXIS_IARG_82_DMWIDTH,S_AXIS_IARG_81_DMWIDTH,S_AXIS_IARG_80_DMWIDTH,S_AXIS_IARG_79_DMWIDTH,S_AXIS_IARG_78_DMWIDTH,S_AXIS_IARG_77_DMWIDTH,S_AXIS_IARG_76_DMWIDTH,S_AXIS_IARG_75_DMWIDTH,S_AXIS_IARG_74_DMWIDTH,S_AXIS_IARG_73_DMWIDTH,S_AXIS_IARG_72_DMWIDTH,S_AXIS_IARG_71_DMWIDTH,S_AXIS_IARG_70_DMWIDTH,S_AXIS_IARG_69_DMWIDTH,S_AXIS_IARG_68_DMWIDTH,S_AXIS_IARG_67_DMWIDTH,S_AXIS_IARG_66_DMWIDTH,S_AXIS_IARG_65_DMWIDTH,S_AXIS_IARG_64_DMWIDTH,S_AXIS_IARG_63_DMWIDTH,S_AXIS_IARG_62_DMWIDTH,S_AXIS_IARG_61_DMWIDTH,S_AXIS_IARG_60_DMWIDTH,S_AXIS_IARG_59_DMWIDTH,S_AXIS_IARG_58_DMWIDTH,S_AXIS_IARG_57_DMWIDTH,S_AXIS_IARG_56_DMWIDTH,S_AXIS_IARG_55_DMWIDTH,S_AXIS_IARG_54_DMWIDTH,S_AXIS_IARG_53_DMWIDTH,S_AXIS_IARG_52_DMWIDTH,S_AXIS_IARG_51_DMWIDTH,S_AXIS_IARG_50_DMWIDTH,S_AXIS_IARG_49_DMWIDTH,S_AXIS_IARG_48_DMWIDTH,S_AXIS_IARG_47_DMWIDTH,S_AXIS_IARG_46_DMWIDTH,S_AXIS_IARG_45_DMWIDTH,S_AXIS_IARG_44_DMWIDTH,S_AXIS_IARG_43_DMWIDTH,S_AXIS_IARG_42_DMWIDTH,S_AXIS_IARG_41_DMWIDTH,S_AXIS_IARG_40_DMWIDTH,S_AXIS_IARG_39_DMWIDTH,S_AXIS_IARG_38_DMWIDTH,S_AXIS_IARG_37_DMWIDTH,S_AXIS_IARG_36_DMWIDTH,S_AXIS_IARG_35_DMWIDTH,S_AXIS_IARG_34_DMWIDTH,S_AXIS_IARG_33_DMWIDTH,S_AXIS_IARG_32_DMWIDTH,S_AXIS_IARG_31_DMWIDTH,S_AXIS_IARG_30_DMWIDTH,S_AXIS_IARG_29_DMWIDTH,S_AXIS_IARG_28_DMWIDTH,S_AXIS_IARG_27_DMWIDTH,S_AXIS_IARG_26_DMWIDTH,S_AXIS_IARG_25_DMWIDTH,S_AXIS_IARG_24_DMWIDTH,S_AXIS_IARG_23_DMWIDTH,S_AXIS_IARG_22_DMWIDTH,S_AXIS_IARG_21_DMWIDTH,S_AXIS_IARG_20_DMWIDTH,S_AXIS_IARG_19_DMWIDTH,S_AXIS_IARG_18_DMWIDTH,S_AXIS_IARG_17_DMWIDTH,S_AXIS_IARG_16_DMWIDTH,S_AXIS_IARG_15_DMWIDTH,S_AXIS_IARG_14_DMWIDTH,S_AXIS_IARG_13_DMWIDTH,S_AXIS_IARG_12_DMWIDTH,S_AXIS_IARG_11_DMWIDTH,S_AXIS_IARG_10_DMWIDTH,S_AXIS_IARG_9_DMWIDTH,S_AXIS_IARG_8_DMWIDTH,S_AXIS_IARG_7_DMWIDTH,S_AXIS_IARG_6_DMWIDTH,S_AXIS_IARG_5_DMWIDTH,S_AXIS_IARG_4_DMWIDTH,S_AXIS_IARG_3_DMWIDTH,S_AXIS_IARG_2_DMWIDTH,S_AXIS_IARG_1_DMWIDTH,S_AXIS_IARG_0_DMWIDTH};
    localparam [(C_MAX_INPUT_AXISs*32)-1:0] C_IS_ASYNC_BIT_ARRAY = {S_AXIS_IARG_127_IS_ASYNC,S_AXIS_IARG_126_IS_ASYNC,S_AXIS_IARG_125_IS_ASYNC,S_AXIS_IARG_124_IS_ASYNC,S_AXIS_IARG_123_IS_ASYNC,S_AXIS_IARG_122_IS_ASYNC,S_AXIS_IARG_121_IS_ASYNC,S_AXIS_IARG_120_IS_ASYNC,S_AXIS_IARG_119_IS_ASYNC,S_AXIS_IARG_118_IS_ASYNC,S_AXIS_IARG_117_IS_ASYNC,S_AXIS_IARG_116_IS_ASYNC,S_AXIS_IARG_115_IS_ASYNC,S_AXIS_IARG_114_IS_ASYNC,S_AXIS_IARG_113_IS_ASYNC,S_AXIS_IARG_112_IS_ASYNC,S_AXIS_IARG_111_IS_ASYNC,S_AXIS_IARG_110_IS_ASYNC,S_AXIS_IARG_109_IS_ASYNC,S_AXIS_IARG_108_IS_ASYNC,S_AXIS_IARG_107_IS_ASYNC,S_AXIS_IARG_106_IS_ASYNC,S_AXIS_IARG_105_IS_ASYNC,S_AXIS_IARG_104_IS_ASYNC,S_AXIS_IARG_103_IS_ASYNC,S_AXIS_IARG_102_IS_ASYNC,S_AXIS_IARG_101_IS_ASYNC,S_AXIS_IARG_100_IS_ASYNC,S_AXIS_IARG_99_IS_ASYNC,S_AXIS_IARG_98_IS_ASYNC,S_AXIS_IARG_97_IS_ASYNC,S_AXIS_IARG_96_IS_ASYNC,S_AXIS_IARG_95_IS_ASYNC,S_AXIS_IARG_94_IS_ASYNC,S_AXIS_IARG_93_IS_ASYNC,S_AXIS_IARG_92_IS_ASYNC,S_AXIS_IARG_91_IS_ASYNC,S_AXIS_IARG_90_IS_ASYNC,S_AXIS_IARG_89_IS_ASYNC,S_AXIS_IARG_88_IS_ASYNC,S_AXIS_IARG_87_IS_ASYNC,S_AXIS_IARG_86_IS_ASYNC,S_AXIS_IARG_85_IS_ASYNC,S_AXIS_IARG_84_IS_ASYNC,S_AXIS_IARG_83_IS_ASYNC,S_AXIS_IARG_82_IS_ASYNC,S_AXIS_IARG_81_IS_ASYNC,S_AXIS_IARG_80_IS_ASYNC,S_AXIS_IARG_79_IS_ASYNC,S_AXIS_IARG_78_IS_ASYNC,S_AXIS_IARG_77_IS_ASYNC,S_AXIS_IARG_76_IS_ASYNC,S_AXIS_IARG_75_IS_ASYNC,S_AXIS_IARG_74_IS_ASYNC,S_AXIS_IARG_73_IS_ASYNC,S_AXIS_IARG_72_IS_ASYNC,S_AXIS_IARG_71_IS_ASYNC,S_AXIS_IARG_70_IS_ASYNC,S_AXIS_IARG_69_IS_ASYNC,S_AXIS_IARG_68_IS_ASYNC,S_AXIS_IARG_67_IS_ASYNC,S_AXIS_IARG_66_IS_ASYNC,S_AXIS_IARG_65_IS_ASYNC,S_AXIS_IARG_64_IS_ASYNC,S_AXIS_IARG_63_IS_ASYNC,S_AXIS_IARG_62_IS_ASYNC,S_AXIS_IARG_61_IS_ASYNC,S_AXIS_IARG_60_IS_ASYNC,S_AXIS_IARG_59_IS_ASYNC,S_AXIS_IARG_58_IS_ASYNC,S_AXIS_IARG_57_IS_ASYNC,S_AXIS_IARG_56_IS_ASYNC,S_AXIS_IARG_55_IS_ASYNC,S_AXIS_IARG_54_IS_ASYNC,S_AXIS_IARG_53_IS_ASYNC,S_AXIS_IARG_52_IS_ASYNC,S_AXIS_IARG_51_IS_ASYNC,S_AXIS_IARG_50_IS_ASYNC,S_AXIS_IARG_49_IS_ASYNC,S_AXIS_IARG_48_IS_ASYNC,S_AXIS_IARG_47_IS_ASYNC,S_AXIS_IARG_46_IS_ASYNC,S_AXIS_IARG_45_IS_ASYNC,S_AXIS_IARG_44_IS_ASYNC,S_AXIS_IARG_43_IS_ASYNC,S_AXIS_IARG_42_IS_ASYNC,S_AXIS_IARG_41_IS_ASYNC,S_AXIS_IARG_40_IS_ASYNC,S_AXIS_IARG_39_IS_ASYNC,S_AXIS_IARG_38_IS_ASYNC,S_AXIS_IARG_37_IS_ASYNC,S_AXIS_IARG_36_IS_ASYNC,S_AXIS_IARG_35_IS_ASYNC,S_AXIS_IARG_34_IS_ASYNC,S_AXIS_IARG_33_IS_ASYNC,S_AXIS_IARG_32_IS_ASYNC,S_AXIS_IARG_31_IS_ASYNC,S_AXIS_IARG_30_IS_ASYNC,S_AXIS_IARG_29_IS_ASYNC,S_AXIS_IARG_28_IS_ASYNC,S_AXIS_IARG_27_IS_ASYNC,S_AXIS_IARG_26_IS_ASYNC,S_AXIS_IARG_25_IS_ASYNC,S_AXIS_IARG_24_IS_ASYNC,S_AXIS_IARG_23_IS_ASYNC,S_AXIS_IARG_22_IS_ASYNC,S_AXIS_IARG_21_IS_ASYNC,S_AXIS_IARG_20_IS_ASYNC,S_AXIS_IARG_19_IS_ASYNC,S_AXIS_IARG_18_IS_ASYNC,S_AXIS_IARG_17_IS_ASYNC,S_AXIS_IARG_16_IS_ASYNC,S_AXIS_IARG_15_IS_ASYNC,S_AXIS_IARG_14_IS_ASYNC,S_AXIS_IARG_13_IS_ASYNC,S_AXIS_IARG_12_IS_ASYNC,S_AXIS_IARG_11_IS_ASYNC,S_AXIS_IARG_10_IS_ASYNC,S_AXIS_IARG_9_IS_ASYNC,S_AXIS_IARG_8_IS_ASYNC,S_AXIS_IARG_7_IS_ASYNC,S_AXIS_IARG_6_IS_ASYNC,S_AXIS_IARG_5_IS_ASYNC,S_AXIS_IARG_4_IS_ASYNC,S_AXIS_IARG_3_IS_ASYNC,S_AXIS_IARG_2_IS_ASYNC,S_AXIS_IARG_1_IS_ASYNC,S_AXIS_IARG_0_IS_ASYNC};
    
    wire [C_NUM_INPUT_AXISs-1:0] axis_clk;
    wire [C_NUM_INPUT_AXISs-1:0] axis_rst;
    
    wire [C_NUM_INPUT_AXISs-1:0] dm_tlast;
    wire [C_NUM_INPUT_AXISs-1:0] dm_tvalid;
    wire [C_MAX_BIT_WIDTH/8-1:0] dm_tkeep [C_NUM_INPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] dm_tstrb [C_NUM_INPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0]   dm_tdata [C_NUM_INPUT_AXISs-1:0];
    wire [C_NUM_INPUT_AXISs-1:0] dm_tready;
    
    wire [C_NUM_INPUT_AXISs-1:0] dwconv_tlast;
    wire [C_NUM_INPUT_AXISs-1:0] dwconv_tvalid;
    wire [C_MAX_BIT_WIDTH-1:0] dwconv_tdata [C_NUM_INPUT_AXISs-1:0];
    wire [C_NUM_INPUT_AXISs-1:0] dwconv_tready;
    
    wire [C_NUM_INPUT_AXISs-1:0] buf_tlast;
    wire [C_NUM_INPUT_AXISs-1:0] buf_tvalid;
    wire [C_MAX_BIT_WIDTH-1:0] buf_tdata [C_NUM_INPUT_AXISs-1:0];
    wire [C_NUM_INPUT_AXISs-1:0] buf_tready;
    
    wire [C_NUM_INPUT_AXISs-1:0] ap_tlast;
    wire [C_NUM_INPUT_AXISs-1:0] ap_tvalid;
    wire [C_MAX_BIT_WIDTH/8-1:0] ap_tkeep [C_NUM_INPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] ap_tstrb [C_NUM_INPUT_AXISs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0]   ap_tdata [C_NUM_INPUT_AXISs-1:0];
    wire [C_NUM_INPUT_AXISs-1:0] ap_tready;
    
    //assign inputs to buses, and buses to outputs
    generate
        if(C_NUM_INPUT_AXISs > 0) begin
            assign axis_clk[0] = s_axis_iarg_0_aclk;
            assign axis_rst[0] = s_axis_iarg_0_aresetn;
            assign dm_tlast[0] = s_axis_iarg_0_tlast;
            assign dm_tvalid[0] = s_axis_iarg_0_tvalid;
            assign dm_tkeep[0][S_AXIS_IARG_0_DMWIDTH/8-1:0] = s_axis_iarg_0_tkeep;
            assign dm_tstrb[0][S_AXIS_IARG_0_DMWIDTH/8-1:0] = s_axis_iarg_0_tstrb;
            assign dm_tdata[0][S_AXIS_IARG_0_DMWIDTH-1:0] = s_axis_iarg_0_tdata;
            assign s_axis_iarg_0_tready = dm_tready[0];
            assign ap_axis_iarg_0_tlast = ap_tlast[0];
            assign ap_axis_iarg_0_tvalid = ap_tvalid[0];
            assign ap_axis_iarg_0_tkeep = ap_tkeep[0][S_AXIS_IARG_0_WIDTH/8-1:0];
            assign ap_axis_iarg_0_tstrb = ap_tstrb[0][S_AXIS_IARG_0_WIDTH/8-1:0];
            assign ap_axis_iarg_0_tdata = ap_tdata[0][S_AXIS_IARG_0_WIDTH-1:0];
            assign ap_tready[0] = ap_axis_iarg_0_tready;
        end
        if(C_NUM_INPUT_AXISs > 1) begin
            assign axis_clk[1] = s_axis_iarg_1_aclk;
            assign axis_rst[1] = s_axis_iarg_1_aresetn;
            assign dm_tlast[1] = s_axis_iarg_1_tlast;
            assign dm_tvalid[1] = s_axis_iarg_1_tvalid;
            assign dm_tkeep[1][S_AXIS_IARG_1_DMWIDTH/8-1:0] = s_axis_iarg_1_tkeep;
            assign dm_tstrb[1][S_AXIS_IARG_1_DMWIDTH/8-1:0] = s_axis_iarg_1_tstrb;
            assign dm_tdata[1][S_AXIS_IARG_1_DMWIDTH-1:0] = s_axis_iarg_1_tdata;
            assign s_axis_iarg_1_tready = dm_tready[1];
            assign ap_axis_iarg_1_tlast = ap_tlast[1];
            assign ap_axis_iarg_1_tvalid = ap_tvalid[1];
            assign ap_axis_iarg_1_tkeep = ap_tkeep[1][S_AXIS_IARG_1_WIDTH/8-1:0];
            assign ap_axis_iarg_1_tstrb = ap_tstrb[1][S_AXIS_IARG_1_WIDTH/8-1:0];
            assign ap_axis_iarg_1_tdata = ap_tdata[1][S_AXIS_IARG_1_WIDTH-1:0];
            assign ap_tready[1] = ap_axis_iarg_1_tready;
        end
        if(C_NUM_INPUT_AXISs > 2) begin
            assign axis_clk[2] = s_axis_iarg_2_aclk;
            assign axis_rst[2] = s_axis_iarg_2_aresetn;
            assign dm_tlast[2] = s_axis_iarg_2_tlast;
            assign dm_tvalid[2] = s_axis_iarg_2_tvalid;
            assign dm_tkeep[2][S_AXIS_IARG_2_DMWIDTH/8-1:0] = s_axis_iarg_2_tkeep;
            assign dm_tstrb[2][S_AXIS_IARG_2_DMWIDTH/8-1:0] = s_axis_iarg_2_tstrb;
            assign dm_tdata[2][S_AXIS_IARG_2_DMWIDTH-1:0] = s_axis_iarg_2_tdata;
            assign s_axis_iarg_2_tready = dm_tready[2];
            assign ap_axis_iarg_2_tlast = ap_tlast[2];
            assign ap_axis_iarg_2_tvalid = ap_tvalid[2];
            assign ap_axis_iarg_2_tkeep = ap_tkeep[2][S_AXIS_IARG_2_WIDTH/8-1:0];
            assign ap_axis_iarg_2_tstrb = ap_tstrb[2][S_AXIS_IARG_2_WIDTH/8-1:0];
            assign ap_axis_iarg_2_tdata = ap_tdata[2][S_AXIS_IARG_2_WIDTH-1:0];
            assign ap_tready[2] = ap_axis_iarg_2_tready;
        end
        if(C_NUM_INPUT_AXISs > 3) begin
            assign axis_clk[3] = s_axis_iarg_3_aclk;
            assign axis_rst[3] = s_axis_iarg_3_aresetn;
            assign dm_tlast[3] = s_axis_iarg_3_tlast;
            assign dm_tvalid[3] = s_axis_iarg_3_tvalid;
            assign dm_tkeep[3][S_AXIS_IARG_3_DMWIDTH/8-1:0] = s_axis_iarg_3_tkeep;
            assign dm_tstrb[3][S_AXIS_IARG_3_DMWIDTH/8-1:0] = s_axis_iarg_3_tstrb;
            assign dm_tdata[3][S_AXIS_IARG_3_DMWIDTH-1:0] = s_axis_iarg_3_tdata;
            assign s_axis_iarg_3_tready = dm_tready[3];
            assign ap_axis_iarg_3_tlast = ap_tlast[3];
            assign ap_axis_iarg_3_tvalid = ap_tvalid[3];
            assign ap_axis_iarg_3_tkeep = ap_tkeep[3][S_AXIS_IARG_3_WIDTH/8-1:0];
            assign ap_axis_iarg_3_tstrb = ap_tstrb[3][S_AXIS_IARG_3_WIDTH/8-1:0];
            assign ap_axis_iarg_3_tdata = ap_tdata[3][S_AXIS_IARG_3_WIDTH-1:0];
            assign ap_tready[3] = ap_axis_iarg_3_tready;
        end
        if(C_NUM_INPUT_AXISs > 4) begin
            assign axis_clk[4] = s_axis_iarg_4_aclk;
            assign axis_rst[4] = s_axis_iarg_4_aresetn;
            assign dm_tlast[4] = s_axis_iarg_4_tlast;
            assign dm_tvalid[4] = s_axis_iarg_4_tvalid;
            assign dm_tkeep[4][S_AXIS_IARG_4_DMWIDTH/8-1:0] = s_axis_iarg_4_tkeep;
            assign dm_tstrb[4][S_AXIS_IARG_4_DMWIDTH/8-1:0] = s_axis_iarg_4_tstrb;
            assign dm_tdata[4][S_AXIS_IARG_4_DMWIDTH-1:0] = s_axis_iarg_4_tdata;
            assign s_axis_iarg_4_tready = dm_tready[4];
            assign ap_axis_iarg_4_tlast = ap_tlast[4];
            assign ap_axis_iarg_4_tvalid = ap_tvalid[4];
            assign ap_axis_iarg_4_tkeep = ap_tkeep[4][S_AXIS_IARG_4_WIDTH/8-1:0];
            assign ap_axis_iarg_4_tstrb = ap_tstrb[4][S_AXIS_IARG_4_WIDTH/8-1:0];
            assign ap_axis_iarg_4_tdata = ap_tdata[4][S_AXIS_IARG_4_WIDTH-1:0];
            assign ap_tready[4] = ap_axis_iarg_4_tready;
        end
        if(C_NUM_INPUT_AXISs > 5) begin
            assign axis_clk[5] = s_axis_iarg_5_aclk;
            assign axis_rst[5] = s_axis_iarg_5_aresetn;
            assign dm_tlast[5] = s_axis_iarg_5_tlast;
            assign dm_tvalid[5] = s_axis_iarg_5_tvalid;
            assign dm_tkeep[5][S_AXIS_IARG_5_DMWIDTH/8-1:0] = s_axis_iarg_5_tkeep;
            assign dm_tstrb[5][S_AXIS_IARG_5_DMWIDTH/8-1:0] = s_axis_iarg_5_tstrb;
            assign dm_tdata[5][S_AXIS_IARG_5_DMWIDTH-1:0] = s_axis_iarg_5_tdata;
            assign s_axis_iarg_5_tready = dm_tready[5];
            assign ap_axis_iarg_5_tlast = ap_tlast[5];
            assign ap_axis_iarg_5_tvalid = ap_tvalid[5];
            assign ap_axis_iarg_5_tkeep = ap_tkeep[5][S_AXIS_IARG_5_WIDTH/8-1:0];
            assign ap_axis_iarg_5_tstrb = ap_tstrb[5][S_AXIS_IARG_5_WIDTH/8-1:0];
            assign ap_axis_iarg_5_tdata = ap_tdata[5][S_AXIS_IARG_5_WIDTH-1:0];
            assign ap_tready[5] = ap_axis_iarg_5_tready;
        end
        if(C_NUM_INPUT_AXISs > 6) begin
            assign axis_clk[6] = s_axis_iarg_6_aclk;
            assign axis_rst[6] = s_axis_iarg_6_aresetn;
            assign dm_tlast[6] = s_axis_iarg_6_tlast;
            assign dm_tvalid[6] = s_axis_iarg_6_tvalid;
            assign dm_tkeep[6][S_AXIS_IARG_6_DMWIDTH/8-1:0] = s_axis_iarg_6_tkeep;
            assign dm_tstrb[6][S_AXIS_IARG_6_DMWIDTH/8-1:0] = s_axis_iarg_6_tstrb;
            assign dm_tdata[6][S_AXIS_IARG_6_DMWIDTH-1:0] = s_axis_iarg_6_tdata;
            assign s_axis_iarg_6_tready = dm_tready[6];
            assign ap_axis_iarg_6_tlast = ap_tlast[6];
            assign ap_axis_iarg_6_tvalid = ap_tvalid[6];
            assign ap_axis_iarg_6_tkeep = ap_tkeep[6][S_AXIS_IARG_6_WIDTH/8-1:0];
            assign ap_axis_iarg_6_tstrb = ap_tstrb[6][S_AXIS_IARG_6_WIDTH/8-1:0];
            assign ap_axis_iarg_6_tdata = ap_tdata[6][S_AXIS_IARG_6_WIDTH-1:0];
            assign ap_tready[6] = ap_axis_iarg_6_tready;
        end
        if(C_NUM_INPUT_AXISs > 7) begin
            assign axis_clk[7] = s_axis_iarg_7_aclk;
            assign axis_rst[7] = s_axis_iarg_7_aresetn;
            assign dm_tlast[7] = s_axis_iarg_7_tlast;
            assign dm_tvalid[7] = s_axis_iarg_7_tvalid;
            assign dm_tkeep[7][S_AXIS_IARG_7_DMWIDTH/8-1:0] = s_axis_iarg_7_tkeep;
            assign dm_tstrb[7][S_AXIS_IARG_7_DMWIDTH/8-1:0] = s_axis_iarg_7_tstrb;
            assign dm_tdata[7][S_AXIS_IARG_7_DMWIDTH-1:0] = s_axis_iarg_7_tdata;
            assign s_axis_iarg_7_tready = dm_tready[7];
            assign ap_axis_iarg_7_tlast = ap_tlast[7];
            assign ap_axis_iarg_7_tvalid = ap_tvalid[7];
            assign ap_axis_iarg_7_tkeep = ap_tkeep[7][S_AXIS_IARG_7_WIDTH/8-1:0];
            assign ap_axis_iarg_7_tstrb = ap_tstrb[7][S_AXIS_IARG_7_WIDTH/8-1:0];
            assign ap_axis_iarg_7_tdata = ap_tdata[7][S_AXIS_IARG_7_WIDTH-1:0];
            assign ap_tready[7] = ap_axis_iarg_7_tready;
        end
        if(C_NUM_INPUT_AXISs > 8) begin
            assign axis_clk[8] = s_axis_iarg_8_aclk;
            assign axis_rst[8] = s_axis_iarg_8_aresetn;
            assign dm_tlast[8] = s_axis_iarg_8_tlast;
            assign dm_tvalid[8] = s_axis_iarg_8_tvalid;
            assign dm_tkeep[8][S_AXIS_IARG_8_DMWIDTH/8-1:0] = s_axis_iarg_8_tkeep;
            assign dm_tstrb[8][S_AXIS_IARG_8_DMWIDTH/8-1:0] = s_axis_iarg_8_tstrb;
            assign dm_tdata[8][S_AXIS_IARG_8_DMWIDTH-1:0] = s_axis_iarg_8_tdata;
            assign s_axis_iarg_8_tready = dm_tready[8];
            assign ap_axis_iarg_8_tlast = ap_tlast[8];
            assign ap_axis_iarg_8_tvalid = ap_tvalid[8];
            assign ap_axis_iarg_8_tkeep = ap_tkeep[8][S_AXIS_IARG_8_WIDTH/8-1:0];
            assign ap_axis_iarg_8_tstrb = ap_tstrb[8][S_AXIS_IARG_8_WIDTH/8-1:0];
            assign ap_axis_iarg_8_tdata = ap_tdata[8][S_AXIS_IARG_8_WIDTH-1:0];
            assign ap_tready[8] = ap_axis_iarg_8_tready;
        end
        if(C_NUM_INPUT_AXISs > 9) begin
            assign axis_clk[9] = s_axis_iarg_9_aclk;
            assign axis_rst[9] = s_axis_iarg_9_aresetn;
            assign dm_tlast[9] = s_axis_iarg_9_tlast;
            assign dm_tvalid[9] = s_axis_iarg_9_tvalid;
            assign dm_tkeep[9][S_AXIS_IARG_9_DMWIDTH/8-1:0] = s_axis_iarg_9_tkeep;
            assign dm_tstrb[9][S_AXIS_IARG_9_DMWIDTH/8-1:0] = s_axis_iarg_9_tstrb;
            assign dm_tdata[9][S_AXIS_IARG_9_DMWIDTH-1:0] = s_axis_iarg_9_tdata;
            assign s_axis_iarg_9_tready = dm_tready[9];
            assign ap_axis_iarg_9_tlast = ap_tlast[9];
            assign ap_axis_iarg_9_tvalid = ap_tvalid[9];
            assign ap_axis_iarg_9_tkeep = ap_tkeep[9][S_AXIS_IARG_9_WIDTH/8-1:0];
            assign ap_axis_iarg_9_tstrb = ap_tstrb[9][S_AXIS_IARG_9_WIDTH/8-1:0];
            assign ap_axis_iarg_9_tdata = ap_tdata[9][S_AXIS_IARG_9_WIDTH-1:0];
            assign ap_tready[9] = ap_axis_iarg_9_tready;
        end
        if(C_NUM_INPUT_AXISs > 10) begin
            assign axis_clk[10] = s_axis_iarg_10_aclk;
            assign axis_rst[10] = s_axis_iarg_10_aresetn;
            assign dm_tlast[10] = s_axis_iarg_10_tlast;
            assign dm_tvalid[10] = s_axis_iarg_10_tvalid;
            assign dm_tkeep[10][S_AXIS_IARG_10_DMWIDTH/8-1:0] = s_axis_iarg_10_tkeep;
            assign dm_tstrb[10][S_AXIS_IARG_10_DMWIDTH/8-1:0] = s_axis_iarg_10_tstrb;
            assign dm_tdata[10][S_AXIS_IARG_10_DMWIDTH-1:0] = s_axis_iarg_10_tdata;
            assign s_axis_iarg_10_tready = dm_tready[10];
            assign ap_axis_iarg_10_tlast = ap_tlast[10];
            assign ap_axis_iarg_10_tvalid = ap_tvalid[10];
            assign ap_axis_iarg_10_tkeep = ap_tkeep[10][S_AXIS_IARG_10_WIDTH/8-1:0];
            assign ap_axis_iarg_10_tstrb = ap_tstrb[10][S_AXIS_IARG_10_WIDTH/8-1:0];
            assign ap_axis_iarg_10_tdata = ap_tdata[10][S_AXIS_IARG_10_WIDTH-1:0];
            assign ap_tready[10] = ap_axis_iarg_10_tready;
        end
        if(C_NUM_INPUT_AXISs > 11) begin
            assign axis_clk[11] = s_axis_iarg_11_aclk;
            assign axis_rst[11] = s_axis_iarg_11_aresetn;
            assign dm_tlast[11] = s_axis_iarg_11_tlast;
            assign dm_tvalid[11] = s_axis_iarg_11_tvalid;
            assign dm_tkeep[11][S_AXIS_IARG_11_DMWIDTH/8-1:0] = s_axis_iarg_11_tkeep;
            assign dm_tstrb[11][S_AXIS_IARG_11_DMWIDTH/8-1:0] = s_axis_iarg_11_tstrb;
            assign dm_tdata[11][S_AXIS_IARG_11_DMWIDTH-1:0] = s_axis_iarg_11_tdata;
            assign s_axis_iarg_11_tready = dm_tready[11];
            assign ap_axis_iarg_11_tlast = ap_tlast[11];
            assign ap_axis_iarg_11_tvalid = ap_tvalid[11];
            assign ap_axis_iarg_11_tkeep = ap_tkeep[11][S_AXIS_IARG_11_WIDTH/8-1:0];
            assign ap_axis_iarg_11_tstrb = ap_tstrb[11][S_AXIS_IARG_11_WIDTH/8-1:0];
            assign ap_axis_iarg_11_tdata = ap_tdata[11][S_AXIS_IARG_11_WIDTH-1:0];
            assign ap_tready[11] = ap_axis_iarg_11_tready;
        end
        if(C_NUM_INPUT_AXISs > 12) begin
            assign axis_clk[12] = s_axis_iarg_12_aclk;
            assign axis_rst[12] = s_axis_iarg_12_aresetn;
            assign dm_tlast[12] = s_axis_iarg_12_tlast;
            assign dm_tvalid[12] = s_axis_iarg_12_tvalid;
            assign dm_tkeep[12][S_AXIS_IARG_12_DMWIDTH/8-1:0] = s_axis_iarg_12_tkeep;
            assign dm_tstrb[12][S_AXIS_IARG_12_DMWIDTH/8-1:0] = s_axis_iarg_12_tstrb;
            assign dm_tdata[12][S_AXIS_IARG_12_DMWIDTH-1:0] = s_axis_iarg_12_tdata;
            assign s_axis_iarg_12_tready = dm_tready[12];
            assign ap_axis_iarg_12_tlast = ap_tlast[12];
            assign ap_axis_iarg_12_tvalid = ap_tvalid[12];
            assign ap_axis_iarg_12_tkeep = ap_tkeep[12][S_AXIS_IARG_12_WIDTH/8-1:0];
            assign ap_axis_iarg_12_tstrb = ap_tstrb[12][S_AXIS_IARG_12_WIDTH/8-1:0];
            assign ap_axis_iarg_12_tdata = ap_tdata[12][S_AXIS_IARG_12_WIDTH-1:0];
            assign ap_tready[12] = ap_axis_iarg_12_tready;
        end
        if(C_NUM_INPUT_AXISs > 13) begin
            assign axis_clk[13] = s_axis_iarg_13_aclk;
            assign axis_rst[13] = s_axis_iarg_13_aresetn;
            assign dm_tlast[13] = s_axis_iarg_13_tlast;
            assign dm_tvalid[13] = s_axis_iarg_13_tvalid;
            assign dm_tkeep[13][S_AXIS_IARG_13_DMWIDTH/8-1:0] = s_axis_iarg_13_tkeep;
            assign dm_tstrb[13][S_AXIS_IARG_13_DMWIDTH/8-1:0] = s_axis_iarg_13_tstrb;
            assign dm_tdata[13][S_AXIS_IARG_13_DMWIDTH-1:0] = s_axis_iarg_13_tdata;
            assign s_axis_iarg_13_tready = dm_tready[13];
            assign ap_axis_iarg_13_tlast = ap_tlast[13];
            assign ap_axis_iarg_13_tvalid = ap_tvalid[13];
            assign ap_axis_iarg_13_tkeep = ap_tkeep[13][S_AXIS_IARG_13_WIDTH/8-1:0];
            assign ap_axis_iarg_13_tstrb = ap_tstrb[13][S_AXIS_IARG_13_WIDTH/8-1:0];
            assign ap_axis_iarg_13_tdata = ap_tdata[13][S_AXIS_IARG_13_WIDTH-1:0];
            assign ap_tready[13] = ap_axis_iarg_13_tready;
        end
        if(C_NUM_INPUT_AXISs > 14) begin
            assign axis_clk[14] = s_axis_iarg_14_aclk;
            assign axis_rst[14] = s_axis_iarg_14_aresetn;
            assign dm_tlast[14] = s_axis_iarg_14_tlast;
            assign dm_tvalid[14] = s_axis_iarg_14_tvalid;
            assign dm_tkeep[14][S_AXIS_IARG_14_DMWIDTH/8-1:0] = s_axis_iarg_14_tkeep;
            assign dm_tstrb[14][S_AXIS_IARG_14_DMWIDTH/8-1:0] = s_axis_iarg_14_tstrb;
            assign dm_tdata[14][S_AXIS_IARG_14_DMWIDTH-1:0] = s_axis_iarg_14_tdata;
            assign s_axis_iarg_14_tready = dm_tready[14];
            assign ap_axis_iarg_14_tlast = ap_tlast[14];
            assign ap_axis_iarg_14_tvalid = ap_tvalid[14];
            assign ap_axis_iarg_14_tkeep = ap_tkeep[14][S_AXIS_IARG_14_WIDTH/8-1:0];
            assign ap_axis_iarg_14_tstrb = ap_tstrb[14][S_AXIS_IARG_14_WIDTH/8-1:0];
            assign ap_axis_iarg_14_tdata = ap_tdata[14][S_AXIS_IARG_14_WIDTH-1:0];
            assign ap_tready[14] = ap_axis_iarg_14_tready;
        end
        if(C_NUM_INPUT_AXISs > 15) begin
            assign axis_clk[15] = s_axis_iarg_15_aclk;
            assign axis_rst[15] = s_axis_iarg_15_aresetn;
            assign dm_tlast[15] = s_axis_iarg_15_tlast;
            assign dm_tvalid[15] = s_axis_iarg_15_tvalid;
            assign dm_tkeep[15][S_AXIS_IARG_15_DMWIDTH/8-1:0] = s_axis_iarg_15_tkeep;
            assign dm_tstrb[15][S_AXIS_IARG_15_DMWIDTH/8-1:0] = s_axis_iarg_15_tstrb;
            assign dm_tdata[15][S_AXIS_IARG_15_DMWIDTH-1:0] = s_axis_iarg_15_tdata;
            assign s_axis_iarg_15_tready = dm_tready[15];
            assign ap_axis_iarg_15_tlast = ap_tlast[15];
            assign ap_axis_iarg_15_tvalid = ap_tvalid[15];
            assign ap_axis_iarg_15_tkeep = ap_tkeep[15][S_AXIS_IARG_15_WIDTH/8-1:0];
            assign ap_axis_iarg_15_tstrb = ap_tstrb[15][S_AXIS_IARG_15_WIDTH/8-1:0];
            assign ap_axis_iarg_15_tdata = ap_tdata[15][S_AXIS_IARG_15_WIDTH-1:0];
            assign ap_tready[15] = ap_axis_iarg_15_tready;
        end
        if(C_NUM_INPUT_AXISs > 16) begin
            assign axis_clk[16] = s_axis_iarg_16_aclk;
            assign axis_rst[16] = s_axis_iarg_16_aresetn;
            assign dm_tlast[16] = s_axis_iarg_16_tlast;
            assign dm_tvalid[16] = s_axis_iarg_16_tvalid;
            assign dm_tkeep[16][S_AXIS_IARG_16_DMWIDTH/8-1:0] = s_axis_iarg_16_tkeep;
            assign dm_tstrb[16][S_AXIS_IARG_16_DMWIDTH/8-1:0] = s_axis_iarg_16_tstrb;
            assign dm_tdata[16][S_AXIS_IARG_16_DMWIDTH-1:0] = s_axis_iarg_16_tdata;
            assign s_axis_iarg_16_tready = dm_tready[16];
            assign ap_axis_iarg_16_tlast = ap_tlast[16];
            assign ap_axis_iarg_16_tvalid = ap_tvalid[16];
            assign ap_axis_iarg_16_tkeep = ap_tkeep[16][S_AXIS_IARG_16_WIDTH/8-1:0];
            assign ap_axis_iarg_16_tstrb = ap_tstrb[16][S_AXIS_IARG_16_WIDTH/8-1:0];
            assign ap_axis_iarg_16_tdata = ap_tdata[16][S_AXIS_IARG_16_WIDTH-1:0];
            assign ap_tready[16] = ap_axis_iarg_16_tready;
        end
        if(C_NUM_INPUT_AXISs > 17) begin
            assign axis_clk[17] = s_axis_iarg_17_aclk;
            assign axis_rst[17] = s_axis_iarg_17_aresetn;
            assign dm_tlast[17] = s_axis_iarg_17_tlast;
            assign dm_tvalid[17] = s_axis_iarg_17_tvalid;
            assign dm_tkeep[17][S_AXIS_IARG_17_DMWIDTH/8-1:0] = s_axis_iarg_17_tkeep;
            assign dm_tstrb[17][S_AXIS_IARG_17_DMWIDTH/8-1:0] = s_axis_iarg_17_tstrb;
            assign dm_tdata[17][S_AXIS_IARG_17_DMWIDTH-1:0] = s_axis_iarg_17_tdata;
            assign s_axis_iarg_17_tready = dm_tready[17];
            assign ap_axis_iarg_17_tlast = ap_tlast[17];
            assign ap_axis_iarg_17_tvalid = ap_tvalid[17];
            assign ap_axis_iarg_17_tkeep = ap_tkeep[17][S_AXIS_IARG_17_WIDTH/8-1:0];
            assign ap_axis_iarg_17_tstrb = ap_tstrb[17][S_AXIS_IARG_17_WIDTH/8-1:0];
            assign ap_axis_iarg_17_tdata = ap_tdata[17][S_AXIS_IARG_17_WIDTH-1:0];
            assign ap_tready[17] = ap_axis_iarg_17_tready;
        end
        if(C_NUM_INPUT_AXISs > 18) begin
            assign axis_clk[18] = s_axis_iarg_18_aclk;
            assign axis_rst[18] = s_axis_iarg_18_aresetn;
            assign dm_tlast[18] = s_axis_iarg_18_tlast;
            assign dm_tvalid[18] = s_axis_iarg_18_tvalid;
            assign dm_tkeep[18][S_AXIS_IARG_18_DMWIDTH/8-1:0] = s_axis_iarg_18_tkeep;
            assign dm_tstrb[18][S_AXIS_IARG_18_DMWIDTH/8-1:0] = s_axis_iarg_18_tstrb;
            assign dm_tdata[18][S_AXIS_IARG_18_DMWIDTH-1:0] = s_axis_iarg_18_tdata;
            assign s_axis_iarg_18_tready = dm_tready[18];
            assign ap_axis_iarg_18_tlast = ap_tlast[18];
            assign ap_axis_iarg_18_tvalid = ap_tvalid[18];
            assign ap_axis_iarg_18_tkeep = ap_tkeep[18][S_AXIS_IARG_18_WIDTH/8-1:0];
            assign ap_axis_iarg_18_tstrb = ap_tstrb[18][S_AXIS_IARG_18_WIDTH/8-1:0];
            assign ap_axis_iarg_18_tdata = ap_tdata[18][S_AXIS_IARG_18_WIDTH-1:0];
            assign ap_tready[18] = ap_axis_iarg_18_tready;
        end
        if(C_NUM_INPUT_AXISs > 19) begin
            assign axis_clk[19] = s_axis_iarg_19_aclk;
            assign axis_rst[19] = s_axis_iarg_19_aresetn;
            assign dm_tlast[19] = s_axis_iarg_19_tlast;
            assign dm_tvalid[19] = s_axis_iarg_19_tvalid;
            assign dm_tkeep[19][S_AXIS_IARG_19_DMWIDTH/8-1:0] = s_axis_iarg_19_tkeep;
            assign dm_tstrb[19][S_AXIS_IARG_19_DMWIDTH/8-1:0] = s_axis_iarg_19_tstrb;
            assign dm_tdata[19][S_AXIS_IARG_19_DMWIDTH-1:0] = s_axis_iarg_19_tdata;
            assign s_axis_iarg_19_tready = dm_tready[19];
            assign ap_axis_iarg_19_tlast = ap_tlast[19];
            assign ap_axis_iarg_19_tvalid = ap_tvalid[19];
            assign ap_axis_iarg_19_tkeep = ap_tkeep[19][S_AXIS_IARG_19_WIDTH/8-1:0];
            assign ap_axis_iarg_19_tstrb = ap_tstrb[19][S_AXIS_IARG_19_WIDTH/8-1:0];
            assign ap_axis_iarg_19_tdata = ap_tdata[19][S_AXIS_IARG_19_WIDTH-1:0];
            assign ap_tready[19] = ap_axis_iarg_19_tready;
        end
        if(C_NUM_INPUT_AXISs > 20) begin
            assign axis_clk[20] = s_axis_iarg_20_aclk;
            assign axis_rst[20] = s_axis_iarg_20_aresetn;
            assign dm_tlast[20] = s_axis_iarg_20_tlast;
            assign dm_tvalid[20] = s_axis_iarg_20_tvalid;
            assign dm_tkeep[20][S_AXIS_IARG_20_DMWIDTH/8-1:0] = s_axis_iarg_20_tkeep;
            assign dm_tstrb[20][S_AXIS_IARG_20_DMWIDTH/8-1:0] = s_axis_iarg_20_tstrb;
            assign dm_tdata[20][S_AXIS_IARG_20_DMWIDTH-1:0] = s_axis_iarg_20_tdata;
            assign s_axis_iarg_20_tready = dm_tready[20];
            assign ap_axis_iarg_20_tlast = ap_tlast[20];
            assign ap_axis_iarg_20_tvalid = ap_tvalid[20];
            assign ap_axis_iarg_20_tkeep = ap_tkeep[20][S_AXIS_IARG_20_WIDTH/8-1:0];
            assign ap_axis_iarg_20_tstrb = ap_tstrb[20][S_AXIS_IARG_20_WIDTH/8-1:0];
            assign ap_axis_iarg_20_tdata = ap_tdata[20][S_AXIS_IARG_20_WIDTH-1:0];
            assign ap_tready[20] = ap_axis_iarg_20_tready;
        end
        if(C_NUM_INPUT_AXISs > 21) begin
            assign axis_clk[21] = s_axis_iarg_21_aclk;
            assign axis_rst[21] = s_axis_iarg_21_aresetn;
            assign dm_tlast[21] = s_axis_iarg_21_tlast;
            assign dm_tvalid[21] = s_axis_iarg_21_tvalid;
            assign dm_tkeep[21][S_AXIS_IARG_21_DMWIDTH/8-1:0] = s_axis_iarg_21_tkeep;
            assign dm_tstrb[21][S_AXIS_IARG_21_DMWIDTH/8-1:0] = s_axis_iarg_21_tstrb;
            assign dm_tdata[21][S_AXIS_IARG_21_DMWIDTH-1:0] = s_axis_iarg_21_tdata;
            assign s_axis_iarg_21_tready = dm_tready[21];
            assign ap_axis_iarg_21_tlast = ap_tlast[21];
            assign ap_axis_iarg_21_tvalid = ap_tvalid[21];
            assign ap_axis_iarg_21_tkeep = ap_tkeep[21][S_AXIS_IARG_21_WIDTH/8-1:0];
            assign ap_axis_iarg_21_tstrb = ap_tstrb[21][S_AXIS_IARG_21_WIDTH/8-1:0];
            assign ap_axis_iarg_21_tdata = ap_tdata[21][S_AXIS_IARG_21_WIDTH-1:0];
            assign ap_tready[21] = ap_axis_iarg_21_tready;
        end
        if(C_NUM_INPUT_AXISs > 22) begin
            assign axis_clk[22] = s_axis_iarg_22_aclk;
            assign axis_rst[22] = s_axis_iarg_22_aresetn;
            assign dm_tlast[22] = s_axis_iarg_22_tlast;
            assign dm_tvalid[22] = s_axis_iarg_22_tvalid;
            assign dm_tkeep[22][S_AXIS_IARG_22_DMWIDTH/8-1:0] = s_axis_iarg_22_tkeep;
            assign dm_tstrb[22][S_AXIS_IARG_22_DMWIDTH/8-1:0] = s_axis_iarg_22_tstrb;
            assign dm_tdata[22][S_AXIS_IARG_22_DMWIDTH-1:0] = s_axis_iarg_22_tdata;
            assign s_axis_iarg_22_tready = dm_tready[22];
            assign ap_axis_iarg_22_tlast = ap_tlast[22];
            assign ap_axis_iarg_22_tvalid = ap_tvalid[22];
            assign ap_axis_iarg_22_tkeep = ap_tkeep[22][S_AXIS_IARG_22_WIDTH/8-1:0];
            assign ap_axis_iarg_22_tstrb = ap_tstrb[22][S_AXIS_IARG_22_WIDTH/8-1:0];
            assign ap_axis_iarg_22_tdata = ap_tdata[22][S_AXIS_IARG_22_WIDTH-1:0];
            assign ap_tready[22] = ap_axis_iarg_22_tready;
        end
        if(C_NUM_INPUT_AXISs > 23) begin
            assign axis_clk[23] = s_axis_iarg_23_aclk;
            assign axis_rst[23] = s_axis_iarg_23_aresetn;
            assign dm_tlast[23] = s_axis_iarg_23_tlast;
            assign dm_tvalid[23] = s_axis_iarg_23_tvalid;
            assign dm_tkeep[23][S_AXIS_IARG_23_DMWIDTH/8-1:0] = s_axis_iarg_23_tkeep;
            assign dm_tstrb[23][S_AXIS_IARG_23_DMWIDTH/8-1:0] = s_axis_iarg_23_tstrb;
            assign dm_tdata[23][S_AXIS_IARG_23_DMWIDTH-1:0] = s_axis_iarg_23_tdata;
            assign s_axis_iarg_23_tready = dm_tready[23];
            assign ap_axis_iarg_23_tlast = ap_tlast[23];
            assign ap_axis_iarg_23_tvalid = ap_tvalid[23];
            assign ap_axis_iarg_23_tkeep = ap_tkeep[23][S_AXIS_IARG_23_WIDTH/8-1:0];
            assign ap_axis_iarg_23_tstrb = ap_tstrb[23][S_AXIS_IARG_23_WIDTH/8-1:0];
            assign ap_axis_iarg_23_tdata = ap_tdata[23][S_AXIS_IARG_23_WIDTH-1:0];
            assign ap_tready[23] = ap_axis_iarg_23_tready;
        end
        if(C_NUM_INPUT_AXISs > 24) begin
            assign axis_clk[24] = s_axis_iarg_24_aclk;
            assign axis_rst[24] = s_axis_iarg_24_aresetn;
            assign dm_tlast[24] = s_axis_iarg_24_tlast;
            assign dm_tvalid[24] = s_axis_iarg_24_tvalid;
            assign dm_tkeep[24][S_AXIS_IARG_24_DMWIDTH/8-1:0] = s_axis_iarg_24_tkeep;
            assign dm_tstrb[24][S_AXIS_IARG_24_DMWIDTH/8-1:0] = s_axis_iarg_24_tstrb;
            assign dm_tdata[24][S_AXIS_IARG_24_DMWIDTH-1:0] = s_axis_iarg_24_tdata;
            assign s_axis_iarg_24_tready = dm_tready[24];
            assign ap_axis_iarg_24_tlast = ap_tlast[24];
            assign ap_axis_iarg_24_tvalid = ap_tvalid[24];
            assign ap_axis_iarg_24_tkeep = ap_tkeep[24][S_AXIS_IARG_24_WIDTH/8-1:0];
            assign ap_axis_iarg_24_tstrb = ap_tstrb[24][S_AXIS_IARG_24_WIDTH/8-1:0];
            assign ap_axis_iarg_24_tdata = ap_tdata[24][S_AXIS_IARG_24_WIDTH-1:0];
            assign ap_tready[24] = ap_axis_iarg_24_tready;
        end
        if(C_NUM_INPUT_AXISs > 25) begin
            assign axis_clk[25] = s_axis_iarg_25_aclk;
            assign axis_rst[25] = s_axis_iarg_25_aresetn;
            assign dm_tlast[25] = s_axis_iarg_25_tlast;
            assign dm_tvalid[25] = s_axis_iarg_25_tvalid;
            assign dm_tkeep[25][S_AXIS_IARG_25_DMWIDTH/8-1:0] = s_axis_iarg_25_tkeep;
            assign dm_tstrb[25][S_AXIS_IARG_25_DMWIDTH/8-1:0] = s_axis_iarg_25_tstrb;
            assign dm_tdata[25][S_AXIS_IARG_25_DMWIDTH-1:0] = s_axis_iarg_25_tdata;
            assign s_axis_iarg_25_tready = dm_tready[25];
            assign ap_axis_iarg_25_tlast = ap_tlast[25];
            assign ap_axis_iarg_25_tvalid = ap_tvalid[25];
            assign ap_axis_iarg_25_tkeep = ap_tkeep[25][S_AXIS_IARG_25_WIDTH/8-1:0];
            assign ap_axis_iarg_25_tstrb = ap_tstrb[25][S_AXIS_IARG_25_WIDTH/8-1:0];
            assign ap_axis_iarg_25_tdata = ap_tdata[25][S_AXIS_IARG_25_WIDTH-1:0];
            assign ap_tready[25] = ap_axis_iarg_25_tready;
        end
        if(C_NUM_INPUT_AXISs > 26) begin
            assign axis_clk[26] = s_axis_iarg_26_aclk;
            assign axis_rst[26] = s_axis_iarg_26_aresetn;
            assign dm_tlast[26] = s_axis_iarg_26_tlast;
            assign dm_tvalid[26] = s_axis_iarg_26_tvalid;
            assign dm_tkeep[26][S_AXIS_IARG_26_DMWIDTH/8-1:0] = s_axis_iarg_26_tkeep;
            assign dm_tstrb[26][S_AXIS_IARG_26_DMWIDTH/8-1:0] = s_axis_iarg_26_tstrb;
            assign dm_tdata[26][S_AXIS_IARG_26_DMWIDTH-1:0] = s_axis_iarg_26_tdata;
            assign s_axis_iarg_26_tready = dm_tready[26];
            assign ap_axis_iarg_26_tlast = ap_tlast[26];
            assign ap_axis_iarg_26_tvalid = ap_tvalid[26];
            assign ap_axis_iarg_26_tkeep = ap_tkeep[26][S_AXIS_IARG_26_WIDTH/8-1:0];
            assign ap_axis_iarg_26_tstrb = ap_tstrb[26][S_AXIS_IARG_26_WIDTH/8-1:0];
            assign ap_axis_iarg_26_tdata = ap_tdata[26][S_AXIS_IARG_26_WIDTH-1:0];
            assign ap_tready[26] = ap_axis_iarg_26_tready;
        end
        if(C_NUM_INPUT_AXISs > 27) begin
            assign axis_clk[27] = s_axis_iarg_27_aclk;
            assign axis_rst[27] = s_axis_iarg_27_aresetn;
            assign dm_tlast[27] = s_axis_iarg_27_tlast;
            assign dm_tvalid[27] = s_axis_iarg_27_tvalid;
            assign dm_tkeep[27][S_AXIS_IARG_27_DMWIDTH/8-1:0] = s_axis_iarg_27_tkeep;
            assign dm_tstrb[27][S_AXIS_IARG_27_DMWIDTH/8-1:0] = s_axis_iarg_27_tstrb;
            assign dm_tdata[27][S_AXIS_IARG_27_DMWIDTH-1:0] = s_axis_iarg_27_tdata;
            assign s_axis_iarg_27_tready = dm_tready[27];
            assign ap_axis_iarg_27_tlast = ap_tlast[27];
            assign ap_axis_iarg_27_tvalid = ap_tvalid[27];
            assign ap_axis_iarg_27_tkeep = ap_tkeep[27][S_AXIS_IARG_27_WIDTH/8-1:0];
            assign ap_axis_iarg_27_tstrb = ap_tstrb[27][S_AXIS_IARG_27_WIDTH/8-1:0];
            assign ap_axis_iarg_27_tdata = ap_tdata[27][S_AXIS_IARG_27_WIDTH-1:0];
            assign ap_tready[27] = ap_axis_iarg_27_tready;
        end
        if(C_NUM_INPUT_AXISs > 28) begin
            assign axis_clk[28] = s_axis_iarg_28_aclk;
            assign axis_rst[28] = s_axis_iarg_28_aresetn;
            assign dm_tlast[28] = s_axis_iarg_28_tlast;
            assign dm_tvalid[28] = s_axis_iarg_28_tvalid;
            assign dm_tkeep[28][S_AXIS_IARG_28_DMWIDTH/8-1:0] = s_axis_iarg_28_tkeep;
            assign dm_tstrb[28][S_AXIS_IARG_28_DMWIDTH/8-1:0] = s_axis_iarg_28_tstrb;
            assign dm_tdata[28][S_AXIS_IARG_28_DMWIDTH-1:0] = s_axis_iarg_28_tdata;
            assign s_axis_iarg_28_tready = dm_tready[28];
            assign ap_axis_iarg_28_tlast = ap_tlast[28];
            assign ap_axis_iarg_28_tvalid = ap_tvalid[28];
            assign ap_axis_iarg_28_tkeep = ap_tkeep[28][S_AXIS_IARG_28_WIDTH/8-1:0];
            assign ap_axis_iarg_28_tstrb = ap_tstrb[28][S_AXIS_IARG_28_WIDTH/8-1:0];
            assign ap_axis_iarg_28_tdata = ap_tdata[28][S_AXIS_IARG_28_WIDTH-1:0];
            assign ap_tready[28] = ap_axis_iarg_28_tready;
        end
        if(C_NUM_INPUT_AXISs > 29) begin
            assign axis_clk[29] = s_axis_iarg_29_aclk;
            assign axis_rst[29] = s_axis_iarg_29_aresetn;
            assign dm_tlast[29] = s_axis_iarg_29_tlast;
            assign dm_tvalid[29] = s_axis_iarg_29_tvalid;
            assign dm_tkeep[29][S_AXIS_IARG_29_DMWIDTH/8-1:0] = s_axis_iarg_29_tkeep;
            assign dm_tstrb[29][S_AXIS_IARG_29_DMWIDTH/8-1:0] = s_axis_iarg_29_tstrb;
            assign dm_tdata[29][S_AXIS_IARG_29_DMWIDTH-1:0] = s_axis_iarg_29_tdata;
            assign s_axis_iarg_29_tready = dm_tready[29];
            assign ap_axis_iarg_29_tlast = ap_tlast[29];
            assign ap_axis_iarg_29_tvalid = ap_tvalid[29];
            assign ap_axis_iarg_29_tkeep = ap_tkeep[29][S_AXIS_IARG_29_WIDTH/8-1:0];
            assign ap_axis_iarg_29_tstrb = ap_tstrb[29][S_AXIS_IARG_29_WIDTH/8-1:0];
            assign ap_axis_iarg_29_tdata = ap_tdata[29][S_AXIS_IARG_29_WIDTH-1:0];
            assign ap_tready[29] = ap_axis_iarg_29_tready;
        end
        if(C_NUM_INPUT_AXISs > 30) begin
            assign axis_clk[30] = s_axis_iarg_30_aclk;
            assign axis_rst[30] = s_axis_iarg_30_aresetn;
            assign dm_tlast[30] = s_axis_iarg_30_tlast;
            assign dm_tvalid[30] = s_axis_iarg_30_tvalid;
            assign dm_tkeep[30][S_AXIS_IARG_30_DMWIDTH/8-1:0] = s_axis_iarg_30_tkeep;
            assign dm_tstrb[30][S_AXIS_IARG_30_DMWIDTH/8-1:0] = s_axis_iarg_30_tstrb;
            assign dm_tdata[30][S_AXIS_IARG_30_DMWIDTH-1:0] = s_axis_iarg_30_tdata;
            assign s_axis_iarg_30_tready = dm_tready[30];
            assign ap_axis_iarg_30_tlast = ap_tlast[30];
            assign ap_axis_iarg_30_tvalid = ap_tvalid[30];
            assign ap_axis_iarg_30_tkeep = ap_tkeep[30][S_AXIS_IARG_30_WIDTH/8-1:0];
            assign ap_axis_iarg_30_tstrb = ap_tstrb[30][S_AXIS_IARG_30_WIDTH/8-1:0];
            assign ap_axis_iarg_30_tdata = ap_tdata[30][S_AXIS_IARG_30_WIDTH-1:0];
            assign ap_tready[30] = ap_axis_iarg_30_tready;
        end
        if(C_NUM_INPUT_AXISs > 31) begin
            assign axis_clk[31] = s_axis_iarg_31_aclk;
            assign axis_rst[31] = s_axis_iarg_31_aresetn;
            assign dm_tlast[31] = s_axis_iarg_31_tlast;
            assign dm_tvalid[31] = s_axis_iarg_31_tvalid;
            assign dm_tkeep[31][S_AXIS_IARG_31_DMWIDTH/8-1:0] = s_axis_iarg_31_tkeep;
            assign dm_tstrb[31][S_AXIS_IARG_31_DMWIDTH/8-1:0] = s_axis_iarg_31_tstrb;
            assign dm_tdata[31][S_AXIS_IARG_31_DMWIDTH-1:0] = s_axis_iarg_31_tdata;
            assign s_axis_iarg_31_tready = dm_tready[31];
            assign ap_axis_iarg_31_tlast = ap_tlast[31];
            assign ap_axis_iarg_31_tvalid = ap_tvalid[31];
            assign ap_axis_iarg_31_tkeep = ap_tkeep[31][S_AXIS_IARG_31_WIDTH/8-1:0];
            assign ap_axis_iarg_31_tstrb = ap_tstrb[31][S_AXIS_IARG_31_WIDTH/8-1:0];
            assign ap_axis_iarg_31_tdata = ap_tdata[31][S_AXIS_IARG_31_WIDTH-1:0];
            assign ap_tready[31] = ap_axis_iarg_31_tready;
        end
        if(C_NUM_INPUT_AXISs > 32) begin
            assign axis_clk[32] = s_axis_iarg_32_aclk;
            assign axis_rst[32] = s_axis_iarg_32_aresetn;
            assign dm_tlast[32] = s_axis_iarg_32_tlast;
            assign dm_tvalid[32] = s_axis_iarg_32_tvalid;
            assign dm_tkeep[32][S_AXIS_IARG_32_DMWIDTH/8-1:0] = s_axis_iarg_32_tkeep;
            assign dm_tstrb[32][S_AXIS_IARG_32_DMWIDTH/8-1:0] = s_axis_iarg_32_tstrb;
            assign dm_tdata[32][S_AXIS_IARG_32_DMWIDTH-1:0] = s_axis_iarg_32_tdata;
            assign s_axis_iarg_32_tready = dm_tready[32];
            assign ap_axis_iarg_32_tlast = ap_tlast[32];
            assign ap_axis_iarg_32_tvalid = ap_tvalid[32];
            assign ap_axis_iarg_32_tkeep = ap_tkeep[32][S_AXIS_IARG_32_WIDTH/8-1:0];
            assign ap_axis_iarg_32_tstrb = ap_tstrb[32][S_AXIS_IARG_32_WIDTH/8-1:0];
            assign ap_axis_iarg_32_tdata = ap_tdata[32][S_AXIS_IARG_32_WIDTH-1:0];
            assign ap_tready[32] = ap_axis_iarg_32_tready;
        end
        if(C_NUM_INPUT_AXISs > 33) begin
            assign axis_clk[33] = s_axis_iarg_33_aclk;
            assign axis_rst[33] = s_axis_iarg_33_aresetn;
            assign dm_tlast[33] = s_axis_iarg_33_tlast;
            assign dm_tvalid[33] = s_axis_iarg_33_tvalid;
            assign dm_tkeep[33][S_AXIS_IARG_33_DMWIDTH/8-1:0] = s_axis_iarg_33_tkeep;
            assign dm_tstrb[33][S_AXIS_IARG_33_DMWIDTH/8-1:0] = s_axis_iarg_33_tstrb;
            assign dm_tdata[33][S_AXIS_IARG_33_DMWIDTH-1:0] = s_axis_iarg_33_tdata;
            assign s_axis_iarg_33_tready = dm_tready[33];
            assign ap_axis_iarg_33_tlast = ap_tlast[33];
            assign ap_axis_iarg_33_tvalid = ap_tvalid[33];
            assign ap_axis_iarg_33_tkeep = ap_tkeep[33][S_AXIS_IARG_33_WIDTH/8-1:0];
            assign ap_axis_iarg_33_tstrb = ap_tstrb[33][S_AXIS_IARG_33_WIDTH/8-1:0];
            assign ap_axis_iarg_33_tdata = ap_tdata[33][S_AXIS_IARG_33_WIDTH-1:0];
            assign ap_tready[33] = ap_axis_iarg_33_tready;
        end
        if(C_NUM_INPUT_AXISs > 34) begin
            assign axis_clk[34] = s_axis_iarg_34_aclk;
            assign axis_rst[34] = s_axis_iarg_34_aresetn;
            assign dm_tlast[34] = s_axis_iarg_34_tlast;
            assign dm_tvalid[34] = s_axis_iarg_34_tvalid;
            assign dm_tkeep[34][S_AXIS_IARG_34_DMWIDTH/8-1:0] = s_axis_iarg_34_tkeep;
            assign dm_tstrb[34][S_AXIS_IARG_34_DMWIDTH/8-1:0] = s_axis_iarg_34_tstrb;
            assign dm_tdata[34][S_AXIS_IARG_34_DMWIDTH-1:0] = s_axis_iarg_34_tdata;
            assign s_axis_iarg_34_tready = dm_tready[34];
            assign ap_axis_iarg_34_tlast = ap_tlast[34];
            assign ap_axis_iarg_34_tvalid = ap_tvalid[34];
            assign ap_axis_iarg_34_tkeep = ap_tkeep[34][S_AXIS_IARG_34_WIDTH/8-1:0];
            assign ap_axis_iarg_34_tstrb = ap_tstrb[34][S_AXIS_IARG_34_WIDTH/8-1:0];
            assign ap_axis_iarg_34_tdata = ap_tdata[34][S_AXIS_IARG_34_WIDTH-1:0];
            assign ap_tready[34] = ap_axis_iarg_34_tready;
        end
        if(C_NUM_INPUT_AXISs > 35) begin
            assign axis_clk[35] = s_axis_iarg_35_aclk;
            assign axis_rst[35] = s_axis_iarg_35_aresetn;
            assign dm_tlast[35] = s_axis_iarg_35_tlast;
            assign dm_tvalid[35] = s_axis_iarg_35_tvalid;
            assign dm_tkeep[35][S_AXIS_IARG_35_DMWIDTH/8-1:0] = s_axis_iarg_35_tkeep;
            assign dm_tstrb[35][S_AXIS_IARG_35_DMWIDTH/8-1:0] = s_axis_iarg_35_tstrb;
            assign dm_tdata[35][S_AXIS_IARG_35_DMWIDTH-1:0] = s_axis_iarg_35_tdata;
            assign s_axis_iarg_35_tready = dm_tready[35];
            assign ap_axis_iarg_35_tlast = ap_tlast[35];
            assign ap_axis_iarg_35_tvalid = ap_tvalid[35];
            assign ap_axis_iarg_35_tkeep = ap_tkeep[35][S_AXIS_IARG_35_WIDTH/8-1:0];
            assign ap_axis_iarg_35_tstrb = ap_tstrb[35][S_AXIS_IARG_35_WIDTH/8-1:0];
            assign ap_axis_iarg_35_tdata = ap_tdata[35][S_AXIS_IARG_35_WIDTH-1:0];
            assign ap_tready[35] = ap_axis_iarg_35_tready;
        end
        if(C_NUM_INPUT_AXISs > 36) begin
            assign axis_clk[36] = s_axis_iarg_36_aclk;
            assign axis_rst[36] = s_axis_iarg_36_aresetn;
            assign dm_tlast[36] = s_axis_iarg_36_tlast;
            assign dm_tvalid[36] = s_axis_iarg_36_tvalid;
            assign dm_tkeep[36][S_AXIS_IARG_36_DMWIDTH/8-1:0] = s_axis_iarg_36_tkeep;
            assign dm_tstrb[36][S_AXIS_IARG_36_DMWIDTH/8-1:0] = s_axis_iarg_36_tstrb;
            assign dm_tdata[36][S_AXIS_IARG_36_DMWIDTH-1:0] = s_axis_iarg_36_tdata;
            assign s_axis_iarg_36_tready = dm_tready[36];
            assign ap_axis_iarg_36_tlast = ap_tlast[36];
            assign ap_axis_iarg_36_tvalid = ap_tvalid[36];
            assign ap_axis_iarg_36_tkeep = ap_tkeep[36][S_AXIS_IARG_36_WIDTH/8-1:0];
            assign ap_axis_iarg_36_tstrb = ap_tstrb[36][S_AXIS_IARG_36_WIDTH/8-1:0];
            assign ap_axis_iarg_36_tdata = ap_tdata[36][S_AXIS_IARG_36_WIDTH-1:0];
            assign ap_tready[36] = ap_axis_iarg_36_tready;
        end
        if(C_NUM_INPUT_AXISs > 37) begin
            assign axis_clk[37] = s_axis_iarg_37_aclk;
            assign axis_rst[37] = s_axis_iarg_37_aresetn;
            assign dm_tlast[37] = s_axis_iarg_37_tlast;
            assign dm_tvalid[37] = s_axis_iarg_37_tvalid;
            assign dm_tkeep[37][S_AXIS_IARG_37_DMWIDTH/8-1:0] = s_axis_iarg_37_tkeep;
            assign dm_tstrb[37][S_AXIS_IARG_37_DMWIDTH/8-1:0] = s_axis_iarg_37_tstrb;
            assign dm_tdata[37][S_AXIS_IARG_37_DMWIDTH-1:0] = s_axis_iarg_37_tdata;
            assign s_axis_iarg_37_tready = dm_tready[37];
            assign ap_axis_iarg_37_tlast = ap_tlast[37];
            assign ap_axis_iarg_37_tvalid = ap_tvalid[37];
            assign ap_axis_iarg_37_tkeep = ap_tkeep[37][S_AXIS_IARG_37_WIDTH/8-1:0];
            assign ap_axis_iarg_37_tstrb = ap_tstrb[37][S_AXIS_IARG_37_WIDTH/8-1:0];
            assign ap_axis_iarg_37_tdata = ap_tdata[37][S_AXIS_IARG_37_WIDTH-1:0];
            assign ap_tready[37] = ap_axis_iarg_37_tready;
        end
        if(C_NUM_INPUT_AXISs > 38) begin
            assign axis_clk[38] = s_axis_iarg_38_aclk;
            assign axis_rst[38] = s_axis_iarg_38_aresetn;
            assign dm_tlast[38] = s_axis_iarg_38_tlast;
            assign dm_tvalid[38] = s_axis_iarg_38_tvalid;
            assign dm_tkeep[38][S_AXIS_IARG_38_DMWIDTH/8-1:0] = s_axis_iarg_38_tkeep;
            assign dm_tstrb[38][S_AXIS_IARG_38_DMWIDTH/8-1:0] = s_axis_iarg_38_tstrb;
            assign dm_tdata[38][S_AXIS_IARG_38_DMWIDTH-1:0] = s_axis_iarg_38_tdata;
            assign s_axis_iarg_38_tready = dm_tready[38];
            assign ap_axis_iarg_38_tlast = ap_tlast[38];
            assign ap_axis_iarg_38_tvalid = ap_tvalid[38];
            assign ap_axis_iarg_38_tkeep = ap_tkeep[38][S_AXIS_IARG_38_WIDTH/8-1:0];
            assign ap_axis_iarg_38_tstrb = ap_tstrb[38][S_AXIS_IARG_38_WIDTH/8-1:0];
            assign ap_axis_iarg_38_tdata = ap_tdata[38][S_AXIS_IARG_38_WIDTH-1:0];
            assign ap_tready[38] = ap_axis_iarg_38_tready;
        end
        if(C_NUM_INPUT_AXISs > 39) begin
            assign axis_clk[39] = s_axis_iarg_39_aclk;
            assign axis_rst[39] = s_axis_iarg_39_aresetn;
            assign dm_tlast[39] = s_axis_iarg_39_tlast;
            assign dm_tvalid[39] = s_axis_iarg_39_tvalid;
            assign dm_tkeep[39][S_AXIS_IARG_39_DMWIDTH/8-1:0] = s_axis_iarg_39_tkeep;
            assign dm_tstrb[39][S_AXIS_IARG_39_DMWIDTH/8-1:0] = s_axis_iarg_39_tstrb;
            assign dm_tdata[39][S_AXIS_IARG_39_DMWIDTH-1:0] = s_axis_iarg_39_tdata;
            assign s_axis_iarg_39_tready = dm_tready[39];
            assign ap_axis_iarg_39_tlast = ap_tlast[39];
            assign ap_axis_iarg_39_tvalid = ap_tvalid[39];
            assign ap_axis_iarg_39_tkeep = ap_tkeep[39][S_AXIS_IARG_39_WIDTH/8-1:0];
            assign ap_axis_iarg_39_tstrb = ap_tstrb[39][S_AXIS_IARG_39_WIDTH/8-1:0];
            assign ap_axis_iarg_39_tdata = ap_tdata[39][S_AXIS_IARG_39_WIDTH-1:0];
            assign ap_tready[39] = ap_axis_iarg_39_tready;
        end
        if(C_NUM_INPUT_AXISs > 40) begin
            assign axis_clk[40] = s_axis_iarg_40_aclk;
            assign axis_rst[40] = s_axis_iarg_40_aresetn;
            assign dm_tlast[40] = s_axis_iarg_40_tlast;
            assign dm_tvalid[40] = s_axis_iarg_40_tvalid;
            assign dm_tkeep[40][S_AXIS_IARG_40_DMWIDTH/8-1:0] = s_axis_iarg_40_tkeep;
            assign dm_tstrb[40][S_AXIS_IARG_40_DMWIDTH/8-1:0] = s_axis_iarg_40_tstrb;
            assign dm_tdata[40][S_AXIS_IARG_40_DMWIDTH-1:0] = s_axis_iarg_40_tdata;
            assign s_axis_iarg_40_tready = dm_tready[40];
            assign ap_axis_iarg_40_tlast = ap_tlast[40];
            assign ap_axis_iarg_40_tvalid = ap_tvalid[40];
            assign ap_axis_iarg_40_tkeep = ap_tkeep[40][S_AXIS_IARG_40_WIDTH/8-1:0];
            assign ap_axis_iarg_40_tstrb = ap_tstrb[40][S_AXIS_IARG_40_WIDTH/8-1:0];
            assign ap_axis_iarg_40_tdata = ap_tdata[40][S_AXIS_IARG_40_WIDTH-1:0];
            assign ap_tready[40] = ap_axis_iarg_40_tready;
        end
        if(C_NUM_INPUT_AXISs > 41) begin
            assign axis_clk[41] = s_axis_iarg_41_aclk;
            assign axis_rst[41] = s_axis_iarg_41_aresetn;
            assign dm_tlast[41] = s_axis_iarg_41_tlast;
            assign dm_tvalid[41] = s_axis_iarg_41_tvalid;
            assign dm_tkeep[41][S_AXIS_IARG_41_DMWIDTH/8-1:0] = s_axis_iarg_41_tkeep;
            assign dm_tstrb[41][S_AXIS_IARG_41_DMWIDTH/8-1:0] = s_axis_iarg_41_tstrb;
            assign dm_tdata[41][S_AXIS_IARG_41_DMWIDTH-1:0] = s_axis_iarg_41_tdata;
            assign s_axis_iarg_41_tready = dm_tready[41];
            assign ap_axis_iarg_41_tlast = ap_tlast[41];
            assign ap_axis_iarg_41_tvalid = ap_tvalid[41];
            assign ap_axis_iarg_41_tkeep = ap_tkeep[41][S_AXIS_IARG_41_WIDTH/8-1:0];
            assign ap_axis_iarg_41_tstrb = ap_tstrb[41][S_AXIS_IARG_41_WIDTH/8-1:0];
            assign ap_axis_iarg_41_tdata = ap_tdata[41][S_AXIS_IARG_41_WIDTH-1:0];
            assign ap_tready[41] = ap_axis_iarg_41_tready;
        end
        if(C_NUM_INPUT_AXISs > 42) begin
            assign axis_clk[42] = s_axis_iarg_42_aclk;
            assign axis_rst[42] = s_axis_iarg_42_aresetn;
            assign dm_tlast[42] = s_axis_iarg_42_tlast;
            assign dm_tvalid[42] = s_axis_iarg_42_tvalid;
            assign dm_tkeep[42][S_AXIS_IARG_42_DMWIDTH/8-1:0] = s_axis_iarg_42_tkeep;
            assign dm_tstrb[42][S_AXIS_IARG_42_DMWIDTH/8-1:0] = s_axis_iarg_42_tstrb;
            assign dm_tdata[42][S_AXIS_IARG_42_DMWIDTH-1:0] = s_axis_iarg_42_tdata;
            assign s_axis_iarg_42_tready = dm_tready[42];
            assign ap_axis_iarg_42_tlast = ap_tlast[42];
            assign ap_axis_iarg_42_tvalid = ap_tvalid[42];
            assign ap_axis_iarg_42_tkeep = ap_tkeep[42][S_AXIS_IARG_42_WIDTH/8-1:0];
            assign ap_axis_iarg_42_tstrb = ap_tstrb[42][S_AXIS_IARG_42_WIDTH/8-1:0];
            assign ap_axis_iarg_42_tdata = ap_tdata[42][S_AXIS_IARG_42_WIDTH-1:0];
            assign ap_tready[42] = ap_axis_iarg_42_tready;
        end
        if(C_NUM_INPUT_AXISs > 43) begin
            assign axis_clk[43] = s_axis_iarg_43_aclk;
            assign axis_rst[43] = s_axis_iarg_43_aresetn;
            assign dm_tlast[43] = s_axis_iarg_43_tlast;
            assign dm_tvalid[43] = s_axis_iarg_43_tvalid;
            assign dm_tkeep[43][S_AXIS_IARG_43_DMWIDTH/8-1:0] = s_axis_iarg_43_tkeep;
            assign dm_tstrb[43][S_AXIS_IARG_43_DMWIDTH/8-1:0] = s_axis_iarg_43_tstrb;
            assign dm_tdata[43][S_AXIS_IARG_43_DMWIDTH-1:0] = s_axis_iarg_43_tdata;
            assign s_axis_iarg_43_tready = dm_tready[43];
            assign ap_axis_iarg_43_tlast = ap_tlast[43];
            assign ap_axis_iarg_43_tvalid = ap_tvalid[43];
            assign ap_axis_iarg_43_tkeep = ap_tkeep[43][S_AXIS_IARG_43_WIDTH/8-1:0];
            assign ap_axis_iarg_43_tstrb = ap_tstrb[43][S_AXIS_IARG_43_WIDTH/8-1:0];
            assign ap_axis_iarg_43_tdata = ap_tdata[43][S_AXIS_IARG_43_WIDTH-1:0];
            assign ap_tready[43] = ap_axis_iarg_43_tready;
        end
        if(C_NUM_INPUT_AXISs > 44) begin
            assign axis_clk[44] = s_axis_iarg_44_aclk;
            assign axis_rst[44] = s_axis_iarg_44_aresetn;
            assign dm_tlast[44] = s_axis_iarg_44_tlast;
            assign dm_tvalid[44] = s_axis_iarg_44_tvalid;
            assign dm_tkeep[44][S_AXIS_IARG_44_DMWIDTH/8-1:0] = s_axis_iarg_44_tkeep;
            assign dm_tstrb[44][S_AXIS_IARG_44_DMWIDTH/8-1:0] = s_axis_iarg_44_tstrb;
            assign dm_tdata[44][S_AXIS_IARG_44_DMWIDTH-1:0] = s_axis_iarg_44_tdata;
            assign s_axis_iarg_44_tready = dm_tready[44];
            assign ap_axis_iarg_44_tlast = ap_tlast[44];
            assign ap_axis_iarg_44_tvalid = ap_tvalid[44];
            assign ap_axis_iarg_44_tkeep = ap_tkeep[44][S_AXIS_IARG_44_WIDTH/8-1:0];
            assign ap_axis_iarg_44_tstrb = ap_tstrb[44][S_AXIS_IARG_44_WIDTH/8-1:0];
            assign ap_axis_iarg_44_tdata = ap_tdata[44][S_AXIS_IARG_44_WIDTH-1:0];
            assign ap_tready[44] = ap_axis_iarg_44_tready;
        end
        if(C_NUM_INPUT_AXISs > 45) begin
            assign axis_clk[45] = s_axis_iarg_45_aclk;
            assign axis_rst[45] = s_axis_iarg_45_aresetn;
            assign dm_tlast[45] = s_axis_iarg_45_tlast;
            assign dm_tvalid[45] = s_axis_iarg_45_tvalid;
            assign dm_tkeep[45][S_AXIS_IARG_45_DMWIDTH/8-1:0] = s_axis_iarg_45_tkeep;
            assign dm_tstrb[45][S_AXIS_IARG_45_DMWIDTH/8-1:0] = s_axis_iarg_45_tstrb;
            assign dm_tdata[45][S_AXIS_IARG_45_DMWIDTH-1:0] = s_axis_iarg_45_tdata;
            assign s_axis_iarg_45_tready = dm_tready[45];
            assign ap_axis_iarg_45_tlast = ap_tlast[45];
            assign ap_axis_iarg_45_tvalid = ap_tvalid[45];
            assign ap_axis_iarg_45_tkeep = ap_tkeep[45][S_AXIS_IARG_45_WIDTH/8-1:0];
            assign ap_axis_iarg_45_tstrb = ap_tstrb[45][S_AXIS_IARG_45_WIDTH/8-1:0];
            assign ap_axis_iarg_45_tdata = ap_tdata[45][S_AXIS_IARG_45_WIDTH-1:0];
            assign ap_tready[45] = ap_axis_iarg_45_tready;
        end
        if(C_NUM_INPUT_AXISs > 46) begin
            assign axis_clk[46] = s_axis_iarg_46_aclk;
            assign axis_rst[46] = s_axis_iarg_46_aresetn;
            assign dm_tlast[46] = s_axis_iarg_46_tlast;
            assign dm_tvalid[46] = s_axis_iarg_46_tvalid;
            assign dm_tkeep[46][S_AXIS_IARG_46_DMWIDTH/8-1:0] = s_axis_iarg_46_tkeep;
            assign dm_tstrb[46][S_AXIS_IARG_46_DMWIDTH/8-1:0] = s_axis_iarg_46_tstrb;
            assign dm_tdata[46][S_AXIS_IARG_46_DMWIDTH-1:0] = s_axis_iarg_46_tdata;
            assign s_axis_iarg_46_tready = dm_tready[46];
            assign ap_axis_iarg_46_tlast = ap_tlast[46];
            assign ap_axis_iarg_46_tvalid = ap_tvalid[46];
            assign ap_axis_iarg_46_tkeep = ap_tkeep[46][S_AXIS_IARG_46_WIDTH/8-1:0];
            assign ap_axis_iarg_46_tstrb = ap_tstrb[46][S_AXIS_IARG_46_WIDTH/8-1:0];
            assign ap_axis_iarg_46_tdata = ap_tdata[46][S_AXIS_IARG_46_WIDTH-1:0];
            assign ap_tready[46] = ap_axis_iarg_46_tready;
        end
        if(C_NUM_INPUT_AXISs > 47) begin
            assign axis_clk[47] = s_axis_iarg_47_aclk;
            assign axis_rst[47] = s_axis_iarg_47_aresetn;
            assign dm_tlast[47] = s_axis_iarg_47_tlast;
            assign dm_tvalid[47] = s_axis_iarg_47_tvalid;
            assign dm_tkeep[47][S_AXIS_IARG_47_DMWIDTH/8-1:0] = s_axis_iarg_47_tkeep;
            assign dm_tstrb[47][S_AXIS_IARG_47_DMWIDTH/8-1:0] = s_axis_iarg_47_tstrb;
            assign dm_tdata[47][S_AXIS_IARG_47_DMWIDTH-1:0] = s_axis_iarg_47_tdata;
            assign s_axis_iarg_47_tready = dm_tready[47];
            assign ap_axis_iarg_47_tlast = ap_tlast[47];
            assign ap_axis_iarg_47_tvalid = ap_tvalid[47];
            assign ap_axis_iarg_47_tkeep = ap_tkeep[47][S_AXIS_IARG_47_WIDTH/8-1:0];
            assign ap_axis_iarg_47_tstrb = ap_tstrb[47][S_AXIS_IARG_47_WIDTH/8-1:0];
            assign ap_axis_iarg_47_tdata = ap_tdata[47][S_AXIS_IARG_47_WIDTH-1:0];
            assign ap_tready[47] = ap_axis_iarg_47_tready;
        end
        if(C_NUM_INPUT_AXISs > 48) begin
            assign axis_clk[48] = s_axis_iarg_48_aclk;
            assign axis_rst[48] = s_axis_iarg_48_aresetn;
            assign dm_tlast[48] = s_axis_iarg_48_tlast;
            assign dm_tvalid[48] = s_axis_iarg_48_tvalid;
            assign dm_tkeep[48][S_AXIS_IARG_48_DMWIDTH/8-1:0] = s_axis_iarg_48_tkeep;
            assign dm_tstrb[48][S_AXIS_IARG_48_DMWIDTH/8-1:0] = s_axis_iarg_48_tstrb;
            assign dm_tdata[48][S_AXIS_IARG_48_DMWIDTH-1:0] = s_axis_iarg_48_tdata;
            assign s_axis_iarg_48_tready = dm_tready[48];
            assign ap_axis_iarg_48_tlast = ap_tlast[48];
            assign ap_axis_iarg_48_tvalid = ap_tvalid[48];
            assign ap_axis_iarg_48_tkeep = ap_tkeep[48][S_AXIS_IARG_48_WIDTH/8-1:0];
            assign ap_axis_iarg_48_tstrb = ap_tstrb[48][S_AXIS_IARG_48_WIDTH/8-1:0];
            assign ap_axis_iarg_48_tdata = ap_tdata[48][S_AXIS_IARG_48_WIDTH-1:0];
            assign ap_tready[48] = ap_axis_iarg_48_tready;
        end
        if(C_NUM_INPUT_AXISs > 49) begin
            assign axis_clk[49] = s_axis_iarg_49_aclk;
            assign axis_rst[49] = s_axis_iarg_49_aresetn;
            assign dm_tlast[49] = s_axis_iarg_49_tlast;
            assign dm_tvalid[49] = s_axis_iarg_49_tvalid;
            assign dm_tkeep[49][S_AXIS_IARG_49_DMWIDTH/8-1:0] = s_axis_iarg_49_tkeep;
            assign dm_tstrb[49][S_AXIS_IARG_49_DMWIDTH/8-1:0] = s_axis_iarg_49_tstrb;
            assign dm_tdata[49][S_AXIS_IARG_49_DMWIDTH-1:0] = s_axis_iarg_49_tdata;
            assign s_axis_iarg_49_tready = dm_tready[49];
            assign ap_axis_iarg_49_tlast = ap_tlast[49];
            assign ap_axis_iarg_49_tvalid = ap_tvalid[49];
            assign ap_axis_iarg_49_tkeep = ap_tkeep[49][S_AXIS_IARG_49_WIDTH/8-1:0];
            assign ap_axis_iarg_49_tstrb = ap_tstrb[49][S_AXIS_IARG_49_WIDTH/8-1:0];
            assign ap_axis_iarg_49_tdata = ap_tdata[49][S_AXIS_IARG_49_WIDTH-1:0];
            assign ap_tready[49] = ap_axis_iarg_49_tready;
        end
        if(C_NUM_INPUT_AXISs > 50) begin
            assign axis_clk[50] = s_axis_iarg_50_aclk;
            assign axis_rst[50] = s_axis_iarg_50_aresetn;
            assign dm_tlast[50] = s_axis_iarg_50_tlast;
            assign dm_tvalid[50] = s_axis_iarg_50_tvalid;
            assign dm_tkeep[50][S_AXIS_IARG_50_DMWIDTH/8-1:0] = s_axis_iarg_50_tkeep;
            assign dm_tstrb[50][S_AXIS_IARG_50_DMWIDTH/8-1:0] = s_axis_iarg_50_tstrb;
            assign dm_tdata[50][S_AXIS_IARG_50_DMWIDTH-1:0] = s_axis_iarg_50_tdata;
            assign s_axis_iarg_50_tready = dm_tready[50];
            assign ap_axis_iarg_50_tlast = ap_tlast[50];
            assign ap_axis_iarg_50_tvalid = ap_tvalid[50];
            assign ap_axis_iarg_50_tkeep = ap_tkeep[50][S_AXIS_IARG_50_WIDTH/8-1:0];
            assign ap_axis_iarg_50_tstrb = ap_tstrb[50][S_AXIS_IARG_50_WIDTH/8-1:0];
            assign ap_axis_iarg_50_tdata = ap_tdata[50][S_AXIS_IARG_50_WIDTH-1:0];
            assign ap_tready[50] = ap_axis_iarg_50_tready;
        end
        if(C_NUM_INPUT_AXISs > 51) begin
            assign axis_clk[51] = s_axis_iarg_51_aclk;
            assign axis_rst[51] = s_axis_iarg_51_aresetn;
            assign dm_tlast[51] = s_axis_iarg_51_tlast;
            assign dm_tvalid[51] = s_axis_iarg_51_tvalid;
            assign dm_tkeep[51][S_AXIS_IARG_51_DMWIDTH/8-1:0] = s_axis_iarg_51_tkeep;
            assign dm_tstrb[51][S_AXIS_IARG_51_DMWIDTH/8-1:0] = s_axis_iarg_51_tstrb;
            assign dm_tdata[51][S_AXIS_IARG_51_DMWIDTH-1:0] = s_axis_iarg_51_tdata;
            assign s_axis_iarg_51_tready = dm_tready[51];
            assign ap_axis_iarg_51_tlast = ap_tlast[51];
            assign ap_axis_iarg_51_tvalid = ap_tvalid[51];
            assign ap_axis_iarg_51_tkeep = ap_tkeep[51][S_AXIS_IARG_51_WIDTH/8-1:0];
            assign ap_axis_iarg_51_tstrb = ap_tstrb[51][S_AXIS_IARG_51_WIDTH/8-1:0];
            assign ap_axis_iarg_51_tdata = ap_tdata[51][S_AXIS_IARG_51_WIDTH-1:0];
            assign ap_tready[51] = ap_axis_iarg_51_tready;
        end
        if(C_NUM_INPUT_AXISs > 52) begin
            assign axis_clk[52] = s_axis_iarg_52_aclk;
            assign axis_rst[52] = s_axis_iarg_52_aresetn;
            assign dm_tlast[52] = s_axis_iarg_52_tlast;
            assign dm_tvalid[52] = s_axis_iarg_52_tvalid;
            assign dm_tkeep[52][S_AXIS_IARG_52_DMWIDTH/8-1:0] = s_axis_iarg_52_tkeep;
            assign dm_tstrb[52][S_AXIS_IARG_52_DMWIDTH/8-1:0] = s_axis_iarg_52_tstrb;
            assign dm_tdata[52][S_AXIS_IARG_52_DMWIDTH-1:0] = s_axis_iarg_52_tdata;
            assign s_axis_iarg_52_tready = dm_tready[52];
            assign ap_axis_iarg_52_tlast = ap_tlast[52];
            assign ap_axis_iarg_52_tvalid = ap_tvalid[52];
            assign ap_axis_iarg_52_tkeep = ap_tkeep[52][S_AXIS_IARG_52_WIDTH/8-1:0];
            assign ap_axis_iarg_52_tstrb = ap_tstrb[52][S_AXIS_IARG_52_WIDTH/8-1:0];
            assign ap_axis_iarg_52_tdata = ap_tdata[52][S_AXIS_IARG_52_WIDTH-1:0];
            assign ap_tready[52] = ap_axis_iarg_52_tready;
        end
        if(C_NUM_INPUT_AXISs > 53) begin
            assign axis_clk[53] = s_axis_iarg_53_aclk;
            assign axis_rst[53] = s_axis_iarg_53_aresetn;
            assign dm_tlast[53] = s_axis_iarg_53_tlast;
            assign dm_tvalid[53] = s_axis_iarg_53_tvalid;
            assign dm_tkeep[53][S_AXIS_IARG_53_DMWIDTH/8-1:0] = s_axis_iarg_53_tkeep;
            assign dm_tstrb[53][S_AXIS_IARG_53_DMWIDTH/8-1:0] = s_axis_iarg_53_tstrb;
            assign dm_tdata[53][S_AXIS_IARG_53_DMWIDTH-1:0] = s_axis_iarg_53_tdata;
            assign s_axis_iarg_53_tready = dm_tready[53];
            assign ap_axis_iarg_53_tlast = ap_tlast[53];
            assign ap_axis_iarg_53_tvalid = ap_tvalid[53];
            assign ap_axis_iarg_53_tkeep = ap_tkeep[53][S_AXIS_IARG_53_WIDTH/8-1:0];
            assign ap_axis_iarg_53_tstrb = ap_tstrb[53][S_AXIS_IARG_53_WIDTH/8-1:0];
            assign ap_axis_iarg_53_tdata = ap_tdata[53][S_AXIS_IARG_53_WIDTH-1:0];
            assign ap_tready[53] = ap_axis_iarg_53_tready;
        end
        if(C_NUM_INPUT_AXISs > 54) begin
            assign axis_clk[54] = s_axis_iarg_54_aclk;
            assign axis_rst[54] = s_axis_iarg_54_aresetn;
            assign dm_tlast[54] = s_axis_iarg_54_tlast;
            assign dm_tvalid[54] = s_axis_iarg_54_tvalid;
            assign dm_tkeep[54][S_AXIS_IARG_54_DMWIDTH/8-1:0] = s_axis_iarg_54_tkeep;
            assign dm_tstrb[54][S_AXIS_IARG_54_DMWIDTH/8-1:0] = s_axis_iarg_54_tstrb;
            assign dm_tdata[54][S_AXIS_IARG_54_DMWIDTH-1:0] = s_axis_iarg_54_tdata;
            assign s_axis_iarg_54_tready = dm_tready[54];
            assign ap_axis_iarg_54_tlast = ap_tlast[54];
            assign ap_axis_iarg_54_tvalid = ap_tvalid[54];
            assign ap_axis_iarg_54_tkeep = ap_tkeep[54][S_AXIS_IARG_54_WIDTH/8-1:0];
            assign ap_axis_iarg_54_tstrb = ap_tstrb[54][S_AXIS_IARG_54_WIDTH/8-1:0];
            assign ap_axis_iarg_54_tdata = ap_tdata[54][S_AXIS_IARG_54_WIDTH-1:0];
            assign ap_tready[54] = ap_axis_iarg_54_tready;
        end
        if(C_NUM_INPUT_AXISs > 55) begin
            assign axis_clk[55] = s_axis_iarg_55_aclk;
            assign axis_rst[55] = s_axis_iarg_55_aresetn;
            assign dm_tlast[55] = s_axis_iarg_55_tlast;
            assign dm_tvalid[55] = s_axis_iarg_55_tvalid;
            assign dm_tkeep[55][S_AXIS_IARG_55_DMWIDTH/8-1:0] = s_axis_iarg_55_tkeep;
            assign dm_tstrb[55][S_AXIS_IARG_55_DMWIDTH/8-1:0] = s_axis_iarg_55_tstrb;
            assign dm_tdata[55][S_AXIS_IARG_55_DMWIDTH-1:0] = s_axis_iarg_55_tdata;
            assign s_axis_iarg_55_tready = dm_tready[55];
            assign ap_axis_iarg_55_tlast = ap_tlast[55];
            assign ap_axis_iarg_55_tvalid = ap_tvalid[55];
            assign ap_axis_iarg_55_tkeep = ap_tkeep[55][S_AXIS_IARG_55_WIDTH/8-1:0];
            assign ap_axis_iarg_55_tstrb = ap_tstrb[55][S_AXIS_IARG_55_WIDTH/8-1:0];
            assign ap_axis_iarg_55_tdata = ap_tdata[55][S_AXIS_IARG_55_WIDTH-1:0];
            assign ap_tready[55] = ap_axis_iarg_55_tready;
        end
        if(C_NUM_INPUT_AXISs > 56) begin
            assign axis_clk[56] = s_axis_iarg_56_aclk;
            assign axis_rst[56] = s_axis_iarg_56_aresetn;
            assign dm_tlast[56] = s_axis_iarg_56_tlast;
            assign dm_tvalid[56] = s_axis_iarg_56_tvalid;
            assign dm_tkeep[56][S_AXIS_IARG_56_DMWIDTH/8-1:0] = s_axis_iarg_56_tkeep;
            assign dm_tstrb[56][S_AXIS_IARG_56_DMWIDTH/8-1:0] = s_axis_iarg_56_tstrb;
            assign dm_tdata[56][S_AXIS_IARG_56_DMWIDTH-1:0] = s_axis_iarg_56_tdata;
            assign s_axis_iarg_56_tready = dm_tready[56];
            assign ap_axis_iarg_56_tlast = ap_tlast[56];
            assign ap_axis_iarg_56_tvalid = ap_tvalid[56];
            assign ap_axis_iarg_56_tkeep = ap_tkeep[56][S_AXIS_IARG_56_WIDTH/8-1:0];
            assign ap_axis_iarg_56_tstrb = ap_tstrb[56][S_AXIS_IARG_56_WIDTH/8-1:0];
            assign ap_axis_iarg_56_tdata = ap_tdata[56][S_AXIS_IARG_56_WIDTH-1:0];
            assign ap_tready[56] = ap_axis_iarg_56_tready;
        end
        if(C_NUM_INPUT_AXISs > 57) begin
            assign axis_clk[57] = s_axis_iarg_57_aclk;
            assign axis_rst[57] = s_axis_iarg_57_aresetn;
            assign dm_tlast[57] = s_axis_iarg_57_tlast;
            assign dm_tvalid[57] = s_axis_iarg_57_tvalid;
            assign dm_tkeep[57][S_AXIS_IARG_57_DMWIDTH/8-1:0] = s_axis_iarg_57_tkeep;
            assign dm_tstrb[57][S_AXIS_IARG_57_DMWIDTH/8-1:0] = s_axis_iarg_57_tstrb;
            assign dm_tdata[57][S_AXIS_IARG_57_DMWIDTH-1:0] = s_axis_iarg_57_tdata;
            assign s_axis_iarg_57_tready = dm_tready[57];
            assign ap_axis_iarg_57_tlast = ap_tlast[57];
            assign ap_axis_iarg_57_tvalid = ap_tvalid[57];
            assign ap_axis_iarg_57_tkeep = ap_tkeep[57][S_AXIS_IARG_57_WIDTH/8-1:0];
            assign ap_axis_iarg_57_tstrb = ap_tstrb[57][S_AXIS_IARG_57_WIDTH/8-1:0];
            assign ap_axis_iarg_57_tdata = ap_tdata[57][S_AXIS_IARG_57_WIDTH-1:0];
            assign ap_tready[57] = ap_axis_iarg_57_tready;
        end
        if(C_NUM_INPUT_AXISs > 58) begin
            assign axis_clk[58] = s_axis_iarg_58_aclk;
            assign axis_rst[58] = s_axis_iarg_58_aresetn;
            assign dm_tlast[58] = s_axis_iarg_58_tlast;
            assign dm_tvalid[58] = s_axis_iarg_58_tvalid;
            assign dm_tkeep[58][S_AXIS_IARG_58_DMWIDTH/8-1:0] = s_axis_iarg_58_tkeep;
            assign dm_tstrb[58][S_AXIS_IARG_58_DMWIDTH/8-1:0] = s_axis_iarg_58_tstrb;
            assign dm_tdata[58][S_AXIS_IARG_58_DMWIDTH-1:0] = s_axis_iarg_58_tdata;
            assign s_axis_iarg_58_tready = dm_tready[58];
            assign ap_axis_iarg_58_tlast = ap_tlast[58];
            assign ap_axis_iarg_58_tvalid = ap_tvalid[58];
            assign ap_axis_iarg_58_tkeep = ap_tkeep[58][S_AXIS_IARG_58_WIDTH/8-1:0];
            assign ap_axis_iarg_58_tstrb = ap_tstrb[58][S_AXIS_IARG_58_WIDTH/8-1:0];
            assign ap_axis_iarg_58_tdata = ap_tdata[58][S_AXIS_IARG_58_WIDTH-1:0];
            assign ap_tready[58] = ap_axis_iarg_58_tready;
        end
        if(C_NUM_INPUT_AXISs > 59) begin
            assign axis_clk[59] = s_axis_iarg_59_aclk;
            assign axis_rst[59] = s_axis_iarg_59_aresetn;
            assign dm_tlast[59] = s_axis_iarg_59_tlast;
            assign dm_tvalid[59] = s_axis_iarg_59_tvalid;
            assign dm_tkeep[59][S_AXIS_IARG_59_DMWIDTH/8-1:0] = s_axis_iarg_59_tkeep;
            assign dm_tstrb[59][S_AXIS_IARG_59_DMWIDTH/8-1:0] = s_axis_iarg_59_tstrb;
            assign dm_tdata[59][S_AXIS_IARG_59_DMWIDTH-1:0] = s_axis_iarg_59_tdata;
            assign s_axis_iarg_59_tready = dm_tready[59];
            assign ap_axis_iarg_59_tlast = ap_tlast[59];
            assign ap_axis_iarg_59_tvalid = ap_tvalid[59];
            assign ap_axis_iarg_59_tkeep = ap_tkeep[59][S_AXIS_IARG_59_WIDTH/8-1:0];
            assign ap_axis_iarg_59_tstrb = ap_tstrb[59][S_AXIS_IARG_59_WIDTH/8-1:0];
            assign ap_axis_iarg_59_tdata = ap_tdata[59][S_AXIS_IARG_59_WIDTH-1:0];
            assign ap_tready[59] = ap_axis_iarg_59_tready;
        end
        if(C_NUM_INPUT_AXISs > 60) begin
            assign axis_clk[60] = s_axis_iarg_60_aclk;
            assign axis_rst[60] = s_axis_iarg_60_aresetn;
            assign dm_tlast[60] = s_axis_iarg_60_tlast;
            assign dm_tvalid[60] = s_axis_iarg_60_tvalid;
            assign dm_tkeep[60][S_AXIS_IARG_60_DMWIDTH/8-1:0] = s_axis_iarg_60_tkeep;
            assign dm_tstrb[60][S_AXIS_IARG_60_DMWIDTH/8-1:0] = s_axis_iarg_60_tstrb;
            assign dm_tdata[60][S_AXIS_IARG_60_DMWIDTH-1:0] = s_axis_iarg_60_tdata;
            assign s_axis_iarg_60_tready = dm_tready[60];
            assign ap_axis_iarg_60_tlast = ap_tlast[60];
            assign ap_axis_iarg_60_tvalid = ap_tvalid[60];
            assign ap_axis_iarg_60_tkeep = ap_tkeep[60][S_AXIS_IARG_60_WIDTH/8-1:0];
            assign ap_axis_iarg_60_tstrb = ap_tstrb[60][S_AXIS_IARG_60_WIDTH/8-1:0];
            assign ap_axis_iarg_60_tdata = ap_tdata[60][S_AXIS_IARG_60_WIDTH-1:0];
            assign ap_tready[60] = ap_axis_iarg_60_tready;
        end
        if(C_NUM_INPUT_AXISs > 61) begin
            assign axis_clk[61] = s_axis_iarg_61_aclk;
            assign axis_rst[61] = s_axis_iarg_61_aresetn;
            assign dm_tlast[61] = s_axis_iarg_61_tlast;
            assign dm_tvalid[61] = s_axis_iarg_61_tvalid;
            assign dm_tkeep[61][S_AXIS_IARG_61_DMWIDTH/8-1:0] = s_axis_iarg_61_tkeep;
            assign dm_tstrb[61][S_AXIS_IARG_61_DMWIDTH/8-1:0] = s_axis_iarg_61_tstrb;
            assign dm_tdata[61][S_AXIS_IARG_61_DMWIDTH-1:0] = s_axis_iarg_61_tdata;
            assign s_axis_iarg_61_tready = dm_tready[61];
            assign ap_axis_iarg_61_tlast = ap_tlast[61];
            assign ap_axis_iarg_61_tvalid = ap_tvalid[61];
            assign ap_axis_iarg_61_tkeep = ap_tkeep[61][S_AXIS_IARG_61_WIDTH/8-1:0];
            assign ap_axis_iarg_61_tstrb = ap_tstrb[61][S_AXIS_IARG_61_WIDTH/8-1:0];
            assign ap_axis_iarg_61_tdata = ap_tdata[61][S_AXIS_IARG_61_WIDTH-1:0];
            assign ap_tready[61] = ap_axis_iarg_61_tready;
        end
        if(C_NUM_INPUT_AXISs > 62) begin
            assign axis_clk[62] = s_axis_iarg_62_aclk;
            assign axis_rst[62] = s_axis_iarg_62_aresetn;
            assign dm_tlast[62] = s_axis_iarg_62_tlast;
            assign dm_tvalid[62] = s_axis_iarg_62_tvalid;
            assign dm_tkeep[62][S_AXIS_IARG_62_DMWIDTH/8-1:0] = s_axis_iarg_62_tkeep;
            assign dm_tstrb[62][S_AXIS_IARG_62_DMWIDTH/8-1:0] = s_axis_iarg_62_tstrb;
            assign dm_tdata[62][S_AXIS_IARG_62_DMWIDTH-1:0] = s_axis_iarg_62_tdata;
            assign s_axis_iarg_62_tready = dm_tready[62];
            assign ap_axis_iarg_62_tlast = ap_tlast[62];
            assign ap_axis_iarg_62_tvalid = ap_tvalid[62];
            assign ap_axis_iarg_62_tkeep = ap_tkeep[62][S_AXIS_IARG_62_WIDTH/8-1:0];
            assign ap_axis_iarg_62_tstrb = ap_tstrb[62][S_AXIS_IARG_62_WIDTH/8-1:0];
            assign ap_axis_iarg_62_tdata = ap_tdata[62][S_AXIS_IARG_62_WIDTH-1:0];
            assign ap_tready[62] = ap_axis_iarg_62_tready;
        end
        if(C_NUM_INPUT_AXISs > 63) begin
            assign axis_clk[63] = s_axis_iarg_63_aclk;
            assign axis_rst[63] = s_axis_iarg_63_aresetn;
            assign dm_tlast[63] = s_axis_iarg_63_tlast;
            assign dm_tvalid[63] = s_axis_iarg_63_tvalid;
            assign dm_tkeep[63][S_AXIS_IARG_63_DMWIDTH/8-1:0] = s_axis_iarg_63_tkeep;
            assign dm_tstrb[63][S_AXIS_IARG_63_DMWIDTH/8-1:0] = s_axis_iarg_63_tstrb;
            assign dm_tdata[63][S_AXIS_IARG_63_DMWIDTH-1:0] = s_axis_iarg_63_tdata;
            assign s_axis_iarg_63_tready = dm_tready[63];
            assign ap_axis_iarg_63_tlast = ap_tlast[63];
            assign ap_axis_iarg_63_tvalid = ap_tvalid[63];
            assign ap_axis_iarg_63_tkeep = ap_tkeep[63][S_AXIS_IARG_63_WIDTH/8-1:0];
            assign ap_axis_iarg_63_tstrb = ap_tstrb[63][S_AXIS_IARG_63_WIDTH/8-1:0];
            assign ap_axis_iarg_63_tdata = ap_tdata[63][S_AXIS_IARG_63_WIDTH-1:0];
            assign ap_tready[63] = ap_axis_iarg_63_tready;
        end
        if(C_NUM_INPUT_AXISs > 64) begin
            assign axis_clk[64] = s_axis_iarg_64_aclk;
            assign axis_rst[64] = s_axis_iarg_64_aresetn;
            assign dm_tlast[64] = s_axis_iarg_64_tlast;
            assign dm_tvalid[64] = s_axis_iarg_64_tvalid;
            assign dm_tkeep[64][S_AXIS_IARG_64_DMWIDTH/8-1:0] = s_axis_iarg_64_tkeep;
            assign dm_tstrb[64][S_AXIS_IARG_64_DMWIDTH/8-1:0] = s_axis_iarg_64_tstrb;
            assign dm_tdata[64][S_AXIS_IARG_64_DMWIDTH-1:0] = s_axis_iarg_64_tdata;
            assign s_axis_iarg_64_tready = dm_tready[64];
            assign ap_axis_iarg_64_tlast = ap_tlast[64];
            assign ap_axis_iarg_64_tvalid = ap_tvalid[64];
            assign ap_axis_iarg_64_tkeep = ap_tkeep[64][S_AXIS_IARG_64_WIDTH/8-1:0];
            assign ap_axis_iarg_64_tstrb = ap_tstrb[64][S_AXIS_IARG_64_WIDTH/8-1:0];
            assign ap_axis_iarg_64_tdata = ap_tdata[64][S_AXIS_IARG_64_WIDTH-1:0];
            assign ap_tready[64] = ap_axis_iarg_64_tready;
        end
        if(C_NUM_INPUT_AXISs > 65) begin
            assign axis_clk[65] = s_axis_iarg_65_aclk;
            assign axis_rst[65] = s_axis_iarg_65_aresetn;
            assign dm_tlast[65] = s_axis_iarg_65_tlast;
            assign dm_tvalid[65] = s_axis_iarg_65_tvalid;
            assign dm_tkeep[65][S_AXIS_IARG_65_DMWIDTH/8-1:0] = s_axis_iarg_65_tkeep;
            assign dm_tstrb[65][S_AXIS_IARG_65_DMWIDTH/8-1:0] = s_axis_iarg_65_tstrb;
            assign dm_tdata[65][S_AXIS_IARG_65_DMWIDTH-1:0] = s_axis_iarg_65_tdata;
            assign s_axis_iarg_65_tready = dm_tready[65];
            assign ap_axis_iarg_65_tlast = ap_tlast[65];
            assign ap_axis_iarg_65_tvalid = ap_tvalid[65];
            assign ap_axis_iarg_65_tkeep = ap_tkeep[65][S_AXIS_IARG_65_WIDTH/8-1:0];
            assign ap_axis_iarg_65_tstrb = ap_tstrb[65][S_AXIS_IARG_65_WIDTH/8-1:0];
            assign ap_axis_iarg_65_tdata = ap_tdata[65][S_AXIS_IARG_65_WIDTH-1:0];
            assign ap_tready[65] = ap_axis_iarg_65_tready;
        end
        if(C_NUM_INPUT_AXISs > 66) begin
            assign axis_clk[66] = s_axis_iarg_66_aclk;
            assign axis_rst[66] = s_axis_iarg_66_aresetn;
            assign dm_tlast[66] = s_axis_iarg_66_tlast;
            assign dm_tvalid[66] = s_axis_iarg_66_tvalid;
            assign dm_tkeep[66][S_AXIS_IARG_66_DMWIDTH/8-1:0] = s_axis_iarg_66_tkeep;
            assign dm_tstrb[66][S_AXIS_IARG_66_DMWIDTH/8-1:0] = s_axis_iarg_66_tstrb;
            assign dm_tdata[66][S_AXIS_IARG_66_DMWIDTH-1:0] = s_axis_iarg_66_tdata;
            assign s_axis_iarg_66_tready = dm_tready[66];
            assign ap_axis_iarg_66_tlast = ap_tlast[66];
            assign ap_axis_iarg_66_tvalid = ap_tvalid[66];
            assign ap_axis_iarg_66_tkeep = ap_tkeep[66][S_AXIS_IARG_66_WIDTH/8-1:0];
            assign ap_axis_iarg_66_tstrb = ap_tstrb[66][S_AXIS_IARG_66_WIDTH/8-1:0];
            assign ap_axis_iarg_66_tdata = ap_tdata[66][S_AXIS_IARG_66_WIDTH-1:0];
            assign ap_tready[66] = ap_axis_iarg_66_tready;
        end
        if(C_NUM_INPUT_AXISs > 67) begin
            assign axis_clk[67] = s_axis_iarg_67_aclk;
            assign axis_rst[67] = s_axis_iarg_67_aresetn;
            assign dm_tlast[67] = s_axis_iarg_67_tlast;
            assign dm_tvalid[67] = s_axis_iarg_67_tvalid;
            assign dm_tkeep[67][S_AXIS_IARG_67_DMWIDTH/8-1:0] = s_axis_iarg_67_tkeep;
            assign dm_tstrb[67][S_AXIS_IARG_67_DMWIDTH/8-1:0] = s_axis_iarg_67_tstrb;
            assign dm_tdata[67][S_AXIS_IARG_67_DMWIDTH-1:0] = s_axis_iarg_67_tdata;
            assign s_axis_iarg_67_tready = dm_tready[67];
            assign ap_axis_iarg_67_tlast = ap_tlast[67];
            assign ap_axis_iarg_67_tvalid = ap_tvalid[67];
            assign ap_axis_iarg_67_tkeep = ap_tkeep[67][S_AXIS_IARG_67_WIDTH/8-1:0];
            assign ap_axis_iarg_67_tstrb = ap_tstrb[67][S_AXIS_IARG_67_WIDTH/8-1:0];
            assign ap_axis_iarg_67_tdata = ap_tdata[67][S_AXIS_IARG_67_WIDTH-1:0];
            assign ap_tready[67] = ap_axis_iarg_67_tready;
        end
        if(C_NUM_INPUT_AXISs > 68) begin
            assign axis_clk[68] = s_axis_iarg_68_aclk;
            assign axis_rst[68] = s_axis_iarg_68_aresetn;
            assign dm_tlast[68] = s_axis_iarg_68_tlast;
            assign dm_tvalid[68] = s_axis_iarg_68_tvalid;
            assign dm_tkeep[68][S_AXIS_IARG_68_DMWIDTH/8-1:0] = s_axis_iarg_68_tkeep;
            assign dm_tstrb[68][S_AXIS_IARG_68_DMWIDTH/8-1:0] = s_axis_iarg_68_tstrb;
            assign dm_tdata[68][S_AXIS_IARG_68_DMWIDTH-1:0] = s_axis_iarg_68_tdata;
            assign s_axis_iarg_68_tready = dm_tready[68];
            assign ap_axis_iarg_68_tlast = ap_tlast[68];
            assign ap_axis_iarg_68_tvalid = ap_tvalid[68];
            assign ap_axis_iarg_68_tkeep = ap_tkeep[68][S_AXIS_IARG_68_WIDTH/8-1:0];
            assign ap_axis_iarg_68_tstrb = ap_tstrb[68][S_AXIS_IARG_68_WIDTH/8-1:0];
            assign ap_axis_iarg_68_tdata = ap_tdata[68][S_AXIS_IARG_68_WIDTH-1:0];
            assign ap_tready[68] = ap_axis_iarg_68_tready;
        end
        if(C_NUM_INPUT_AXISs > 69) begin
            assign axis_clk[69] = s_axis_iarg_69_aclk;
            assign axis_rst[69] = s_axis_iarg_69_aresetn;
            assign dm_tlast[69] = s_axis_iarg_69_tlast;
            assign dm_tvalid[69] = s_axis_iarg_69_tvalid;
            assign dm_tkeep[69][S_AXIS_IARG_69_DMWIDTH/8-1:0] = s_axis_iarg_69_tkeep;
            assign dm_tstrb[69][S_AXIS_IARG_69_DMWIDTH/8-1:0] = s_axis_iarg_69_tstrb;
            assign dm_tdata[69][S_AXIS_IARG_69_DMWIDTH-1:0] = s_axis_iarg_69_tdata;
            assign s_axis_iarg_69_tready = dm_tready[69];
            assign ap_axis_iarg_69_tlast = ap_tlast[69];
            assign ap_axis_iarg_69_tvalid = ap_tvalid[69];
            assign ap_axis_iarg_69_tkeep = ap_tkeep[69][S_AXIS_IARG_69_WIDTH/8-1:0];
            assign ap_axis_iarg_69_tstrb = ap_tstrb[69][S_AXIS_IARG_69_WIDTH/8-1:0];
            assign ap_axis_iarg_69_tdata = ap_tdata[69][S_AXIS_IARG_69_WIDTH-1:0];
            assign ap_tready[69] = ap_axis_iarg_69_tready;
        end
        if(C_NUM_INPUT_AXISs > 70) begin
            assign axis_clk[70] = s_axis_iarg_70_aclk;
            assign axis_rst[70] = s_axis_iarg_70_aresetn;
            assign dm_tlast[70] = s_axis_iarg_70_tlast;
            assign dm_tvalid[70] = s_axis_iarg_70_tvalid;
            assign dm_tkeep[70][S_AXIS_IARG_70_DMWIDTH/8-1:0] = s_axis_iarg_70_tkeep;
            assign dm_tstrb[70][S_AXIS_IARG_70_DMWIDTH/8-1:0] = s_axis_iarg_70_tstrb;
            assign dm_tdata[70][S_AXIS_IARG_70_DMWIDTH-1:0] = s_axis_iarg_70_tdata;
            assign s_axis_iarg_70_tready = dm_tready[70];
            assign ap_axis_iarg_70_tlast = ap_tlast[70];
            assign ap_axis_iarg_70_tvalid = ap_tvalid[70];
            assign ap_axis_iarg_70_tkeep = ap_tkeep[70][S_AXIS_IARG_70_WIDTH/8-1:0];
            assign ap_axis_iarg_70_tstrb = ap_tstrb[70][S_AXIS_IARG_70_WIDTH/8-1:0];
            assign ap_axis_iarg_70_tdata = ap_tdata[70][S_AXIS_IARG_70_WIDTH-1:0];
            assign ap_tready[70] = ap_axis_iarg_70_tready;
        end
        if(C_NUM_INPUT_AXISs > 71) begin
            assign axis_clk[71] = s_axis_iarg_71_aclk;
            assign axis_rst[71] = s_axis_iarg_71_aresetn;
            assign dm_tlast[71] = s_axis_iarg_71_tlast;
            assign dm_tvalid[71] = s_axis_iarg_71_tvalid;
            assign dm_tkeep[71][S_AXIS_IARG_71_DMWIDTH/8-1:0] = s_axis_iarg_71_tkeep;
            assign dm_tstrb[71][S_AXIS_IARG_71_DMWIDTH/8-1:0] = s_axis_iarg_71_tstrb;
            assign dm_tdata[71][S_AXIS_IARG_71_DMWIDTH-1:0] = s_axis_iarg_71_tdata;
            assign s_axis_iarg_71_tready = dm_tready[71];
            assign ap_axis_iarg_71_tlast = ap_tlast[71];
            assign ap_axis_iarg_71_tvalid = ap_tvalid[71];
            assign ap_axis_iarg_71_tkeep = ap_tkeep[71][S_AXIS_IARG_71_WIDTH/8-1:0];
            assign ap_axis_iarg_71_tstrb = ap_tstrb[71][S_AXIS_IARG_71_WIDTH/8-1:0];
            assign ap_axis_iarg_71_tdata = ap_tdata[71][S_AXIS_IARG_71_WIDTH-1:0];
            assign ap_tready[71] = ap_axis_iarg_71_tready;
        end
        if(C_NUM_INPUT_AXISs > 72) begin
            assign axis_clk[72] = s_axis_iarg_72_aclk;
            assign axis_rst[72] = s_axis_iarg_72_aresetn;
            assign dm_tlast[72] = s_axis_iarg_72_tlast;
            assign dm_tvalid[72] = s_axis_iarg_72_tvalid;
            assign dm_tkeep[72][S_AXIS_IARG_72_DMWIDTH/8-1:0] = s_axis_iarg_72_tkeep;
            assign dm_tstrb[72][S_AXIS_IARG_72_DMWIDTH/8-1:0] = s_axis_iarg_72_tstrb;
            assign dm_tdata[72][S_AXIS_IARG_72_DMWIDTH-1:0] = s_axis_iarg_72_tdata;
            assign s_axis_iarg_72_tready = dm_tready[72];
            assign ap_axis_iarg_72_tlast = ap_tlast[72];
            assign ap_axis_iarg_72_tvalid = ap_tvalid[72];
            assign ap_axis_iarg_72_tkeep = ap_tkeep[72][S_AXIS_IARG_72_WIDTH/8-1:0];
            assign ap_axis_iarg_72_tstrb = ap_tstrb[72][S_AXIS_IARG_72_WIDTH/8-1:0];
            assign ap_axis_iarg_72_tdata = ap_tdata[72][S_AXIS_IARG_72_WIDTH-1:0];
            assign ap_tready[72] = ap_axis_iarg_72_tready;
        end
        if(C_NUM_INPUT_AXISs > 73) begin
            assign axis_clk[73] = s_axis_iarg_73_aclk;
            assign axis_rst[73] = s_axis_iarg_73_aresetn;
            assign dm_tlast[73] = s_axis_iarg_73_tlast;
            assign dm_tvalid[73] = s_axis_iarg_73_tvalid;
            assign dm_tkeep[73][S_AXIS_IARG_73_DMWIDTH/8-1:0] = s_axis_iarg_73_tkeep;
            assign dm_tstrb[73][S_AXIS_IARG_73_DMWIDTH/8-1:0] = s_axis_iarg_73_tstrb;
            assign dm_tdata[73][S_AXIS_IARG_73_DMWIDTH-1:0] = s_axis_iarg_73_tdata;
            assign s_axis_iarg_73_tready = dm_tready[73];
            assign ap_axis_iarg_73_tlast = ap_tlast[73];
            assign ap_axis_iarg_73_tvalid = ap_tvalid[73];
            assign ap_axis_iarg_73_tkeep = ap_tkeep[73][S_AXIS_IARG_73_WIDTH/8-1:0];
            assign ap_axis_iarg_73_tstrb = ap_tstrb[73][S_AXIS_IARG_73_WIDTH/8-1:0];
            assign ap_axis_iarg_73_tdata = ap_tdata[73][S_AXIS_IARG_73_WIDTH-1:0];
            assign ap_tready[73] = ap_axis_iarg_73_tready;
        end
        if(C_NUM_INPUT_AXISs > 74) begin
            assign axis_clk[74] = s_axis_iarg_74_aclk;
            assign axis_rst[74] = s_axis_iarg_74_aresetn;
            assign dm_tlast[74] = s_axis_iarg_74_tlast;
            assign dm_tvalid[74] = s_axis_iarg_74_tvalid;
            assign dm_tkeep[74][S_AXIS_IARG_74_DMWIDTH/8-1:0] = s_axis_iarg_74_tkeep;
            assign dm_tstrb[74][S_AXIS_IARG_74_DMWIDTH/8-1:0] = s_axis_iarg_74_tstrb;
            assign dm_tdata[74][S_AXIS_IARG_74_DMWIDTH-1:0] = s_axis_iarg_74_tdata;
            assign s_axis_iarg_74_tready = dm_tready[74];
            assign ap_axis_iarg_74_tlast = ap_tlast[74];
            assign ap_axis_iarg_74_tvalid = ap_tvalid[74];
            assign ap_axis_iarg_74_tkeep = ap_tkeep[74][S_AXIS_IARG_74_WIDTH/8-1:0];
            assign ap_axis_iarg_74_tstrb = ap_tstrb[74][S_AXIS_IARG_74_WIDTH/8-1:0];
            assign ap_axis_iarg_74_tdata = ap_tdata[74][S_AXIS_IARG_74_WIDTH-1:0];
            assign ap_tready[74] = ap_axis_iarg_74_tready;
        end
        if(C_NUM_INPUT_AXISs > 75) begin
            assign axis_clk[75] = s_axis_iarg_75_aclk;
            assign axis_rst[75] = s_axis_iarg_75_aresetn;
            assign dm_tlast[75] = s_axis_iarg_75_tlast;
            assign dm_tvalid[75] = s_axis_iarg_75_tvalid;
            assign dm_tkeep[75][S_AXIS_IARG_75_DMWIDTH/8-1:0] = s_axis_iarg_75_tkeep;
            assign dm_tstrb[75][S_AXIS_IARG_75_DMWIDTH/8-1:0] = s_axis_iarg_75_tstrb;
            assign dm_tdata[75][S_AXIS_IARG_75_DMWIDTH-1:0] = s_axis_iarg_75_tdata;
            assign s_axis_iarg_75_tready = dm_tready[75];
            assign ap_axis_iarg_75_tlast = ap_tlast[75];
            assign ap_axis_iarg_75_tvalid = ap_tvalid[75];
            assign ap_axis_iarg_75_tkeep = ap_tkeep[75][S_AXIS_IARG_75_WIDTH/8-1:0];
            assign ap_axis_iarg_75_tstrb = ap_tstrb[75][S_AXIS_IARG_75_WIDTH/8-1:0];
            assign ap_axis_iarg_75_tdata = ap_tdata[75][S_AXIS_IARG_75_WIDTH-1:0];
            assign ap_tready[75] = ap_axis_iarg_75_tready;
        end
        if(C_NUM_INPUT_AXISs > 76) begin
            assign axis_clk[76] = s_axis_iarg_76_aclk;
            assign axis_rst[76] = s_axis_iarg_76_aresetn;
            assign dm_tlast[76] = s_axis_iarg_76_tlast;
            assign dm_tvalid[76] = s_axis_iarg_76_tvalid;
            assign dm_tkeep[76][S_AXIS_IARG_76_DMWIDTH/8-1:0] = s_axis_iarg_76_tkeep;
            assign dm_tstrb[76][S_AXIS_IARG_76_DMWIDTH/8-1:0] = s_axis_iarg_76_tstrb;
            assign dm_tdata[76][S_AXIS_IARG_76_DMWIDTH-1:0] = s_axis_iarg_76_tdata;
            assign s_axis_iarg_76_tready = dm_tready[76];
            assign ap_axis_iarg_76_tlast = ap_tlast[76];
            assign ap_axis_iarg_76_tvalid = ap_tvalid[76];
            assign ap_axis_iarg_76_tkeep = ap_tkeep[76][S_AXIS_IARG_76_WIDTH/8-1:0];
            assign ap_axis_iarg_76_tstrb = ap_tstrb[76][S_AXIS_IARG_76_WIDTH/8-1:0];
            assign ap_axis_iarg_76_tdata = ap_tdata[76][S_AXIS_IARG_76_WIDTH-1:0];
            assign ap_tready[76] = ap_axis_iarg_76_tready;
        end
        if(C_NUM_INPUT_AXISs > 77) begin
            assign axis_clk[77] = s_axis_iarg_77_aclk;
            assign axis_rst[77] = s_axis_iarg_77_aresetn;
            assign dm_tlast[77] = s_axis_iarg_77_tlast;
            assign dm_tvalid[77] = s_axis_iarg_77_tvalid;
            assign dm_tkeep[77][S_AXIS_IARG_77_DMWIDTH/8-1:0] = s_axis_iarg_77_tkeep;
            assign dm_tstrb[77][S_AXIS_IARG_77_DMWIDTH/8-1:0] = s_axis_iarg_77_tstrb;
            assign dm_tdata[77][S_AXIS_IARG_77_DMWIDTH-1:0] = s_axis_iarg_77_tdata;
            assign s_axis_iarg_77_tready = dm_tready[77];
            assign ap_axis_iarg_77_tlast = ap_tlast[77];
            assign ap_axis_iarg_77_tvalid = ap_tvalid[77];
            assign ap_axis_iarg_77_tkeep = ap_tkeep[77][S_AXIS_IARG_77_WIDTH/8-1:0];
            assign ap_axis_iarg_77_tstrb = ap_tstrb[77][S_AXIS_IARG_77_WIDTH/8-1:0];
            assign ap_axis_iarg_77_tdata = ap_tdata[77][S_AXIS_IARG_77_WIDTH-1:0];
            assign ap_tready[77] = ap_axis_iarg_77_tready;
        end
        if(C_NUM_INPUT_AXISs > 78) begin
            assign axis_clk[78] = s_axis_iarg_78_aclk;
            assign axis_rst[78] = s_axis_iarg_78_aresetn;
            assign dm_tlast[78] = s_axis_iarg_78_tlast;
            assign dm_tvalid[78] = s_axis_iarg_78_tvalid;
            assign dm_tkeep[78][S_AXIS_IARG_78_DMWIDTH/8-1:0] = s_axis_iarg_78_tkeep;
            assign dm_tstrb[78][S_AXIS_IARG_78_DMWIDTH/8-1:0] = s_axis_iarg_78_tstrb;
            assign dm_tdata[78][S_AXIS_IARG_78_DMWIDTH-1:0] = s_axis_iarg_78_tdata;
            assign s_axis_iarg_78_tready = dm_tready[78];
            assign ap_axis_iarg_78_tlast = ap_tlast[78];
            assign ap_axis_iarg_78_tvalid = ap_tvalid[78];
            assign ap_axis_iarg_78_tkeep = ap_tkeep[78][S_AXIS_IARG_78_WIDTH/8-1:0];
            assign ap_axis_iarg_78_tstrb = ap_tstrb[78][S_AXIS_IARG_78_WIDTH/8-1:0];
            assign ap_axis_iarg_78_tdata = ap_tdata[78][S_AXIS_IARG_78_WIDTH-1:0];
            assign ap_tready[78] = ap_axis_iarg_78_tready;
        end
        if(C_NUM_INPUT_AXISs > 79) begin
            assign axis_clk[79] = s_axis_iarg_79_aclk;
            assign axis_rst[79] = s_axis_iarg_79_aresetn;
            assign dm_tlast[79] = s_axis_iarg_79_tlast;
            assign dm_tvalid[79] = s_axis_iarg_79_tvalid;
            assign dm_tkeep[79][S_AXIS_IARG_79_DMWIDTH/8-1:0] = s_axis_iarg_79_tkeep;
            assign dm_tstrb[79][S_AXIS_IARG_79_DMWIDTH/8-1:0] = s_axis_iarg_79_tstrb;
            assign dm_tdata[79][S_AXIS_IARG_79_DMWIDTH-1:0] = s_axis_iarg_79_tdata;
            assign s_axis_iarg_79_tready = dm_tready[79];
            assign ap_axis_iarg_79_tlast = ap_tlast[79];
            assign ap_axis_iarg_79_tvalid = ap_tvalid[79];
            assign ap_axis_iarg_79_tkeep = ap_tkeep[79][S_AXIS_IARG_79_WIDTH/8-1:0];
            assign ap_axis_iarg_79_tstrb = ap_tstrb[79][S_AXIS_IARG_79_WIDTH/8-1:0];
            assign ap_axis_iarg_79_tdata = ap_tdata[79][S_AXIS_IARG_79_WIDTH-1:0];
            assign ap_tready[79] = ap_axis_iarg_79_tready;
        end
        if(C_NUM_INPUT_AXISs > 80) begin
            assign axis_clk[80] = s_axis_iarg_80_aclk;
            assign axis_rst[80] = s_axis_iarg_80_aresetn;
            assign dm_tlast[80] = s_axis_iarg_80_tlast;
            assign dm_tvalid[80] = s_axis_iarg_80_tvalid;
            assign dm_tkeep[80][S_AXIS_IARG_80_DMWIDTH/8-1:0] = s_axis_iarg_80_tkeep;
            assign dm_tstrb[80][S_AXIS_IARG_80_DMWIDTH/8-1:0] = s_axis_iarg_80_tstrb;
            assign dm_tdata[80][S_AXIS_IARG_80_DMWIDTH-1:0] = s_axis_iarg_80_tdata;
            assign s_axis_iarg_80_tready = dm_tready[80];
            assign ap_axis_iarg_80_tlast = ap_tlast[80];
            assign ap_axis_iarg_80_tvalid = ap_tvalid[80];
            assign ap_axis_iarg_80_tkeep = ap_tkeep[80][S_AXIS_IARG_80_WIDTH/8-1:0];
            assign ap_axis_iarg_80_tstrb = ap_tstrb[80][S_AXIS_IARG_80_WIDTH/8-1:0];
            assign ap_axis_iarg_80_tdata = ap_tdata[80][S_AXIS_IARG_80_WIDTH-1:0];
            assign ap_tready[80] = ap_axis_iarg_80_tready;
        end
        if(C_NUM_INPUT_AXISs > 81) begin
            assign axis_clk[81] = s_axis_iarg_81_aclk;
            assign axis_rst[81] = s_axis_iarg_81_aresetn;
            assign dm_tlast[81] = s_axis_iarg_81_tlast;
            assign dm_tvalid[81] = s_axis_iarg_81_tvalid;
            assign dm_tkeep[81][S_AXIS_IARG_81_DMWIDTH/8-1:0] = s_axis_iarg_81_tkeep;
            assign dm_tstrb[81][S_AXIS_IARG_81_DMWIDTH/8-1:0] = s_axis_iarg_81_tstrb;
            assign dm_tdata[81][S_AXIS_IARG_81_DMWIDTH-1:0] = s_axis_iarg_81_tdata;
            assign s_axis_iarg_81_tready = dm_tready[81];
            assign ap_axis_iarg_81_tlast = ap_tlast[81];
            assign ap_axis_iarg_81_tvalid = ap_tvalid[81];
            assign ap_axis_iarg_81_tkeep = ap_tkeep[81][S_AXIS_IARG_81_WIDTH/8-1:0];
            assign ap_axis_iarg_81_tstrb = ap_tstrb[81][S_AXIS_IARG_81_WIDTH/8-1:0];
            assign ap_axis_iarg_81_tdata = ap_tdata[81][S_AXIS_IARG_81_WIDTH-1:0];
            assign ap_tready[81] = ap_axis_iarg_81_tready;
        end
        if(C_NUM_INPUT_AXISs > 82) begin
            assign axis_clk[82] = s_axis_iarg_82_aclk;
            assign axis_rst[82] = s_axis_iarg_82_aresetn;
            assign dm_tlast[82] = s_axis_iarg_82_tlast;
            assign dm_tvalid[82] = s_axis_iarg_82_tvalid;
            assign dm_tkeep[82][S_AXIS_IARG_82_DMWIDTH/8-1:0] = s_axis_iarg_82_tkeep;
            assign dm_tstrb[82][S_AXIS_IARG_82_DMWIDTH/8-1:0] = s_axis_iarg_82_tstrb;
            assign dm_tdata[82][S_AXIS_IARG_82_DMWIDTH-1:0] = s_axis_iarg_82_tdata;
            assign s_axis_iarg_82_tready = dm_tready[82];
            assign ap_axis_iarg_82_tlast = ap_tlast[82];
            assign ap_axis_iarg_82_tvalid = ap_tvalid[82];
            assign ap_axis_iarg_82_tkeep = ap_tkeep[82][S_AXIS_IARG_82_WIDTH/8-1:0];
            assign ap_axis_iarg_82_tstrb = ap_tstrb[82][S_AXIS_IARG_82_WIDTH/8-1:0];
            assign ap_axis_iarg_82_tdata = ap_tdata[82][S_AXIS_IARG_82_WIDTH-1:0];
            assign ap_tready[82] = ap_axis_iarg_82_tready;
        end
        if(C_NUM_INPUT_AXISs > 83) begin
            assign axis_clk[83] = s_axis_iarg_83_aclk;
            assign axis_rst[83] = s_axis_iarg_83_aresetn;
            assign dm_tlast[83] = s_axis_iarg_83_tlast;
            assign dm_tvalid[83] = s_axis_iarg_83_tvalid;
            assign dm_tkeep[83][S_AXIS_IARG_83_DMWIDTH/8-1:0] = s_axis_iarg_83_tkeep;
            assign dm_tstrb[83][S_AXIS_IARG_83_DMWIDTH/8-1:0] = s_axis_iarg_83_tstrb;
            assign dm_tdata[83][S_AXIS_IARG_83_DMWIDTH-1:0] = s_axis_iarg_83_tdata;
            assign s_axis_iarg_83_tready = dm_tready[83];
            assign ap_axis_iarg_83_tlast = ap_tlast[83];
            assign ap_axis_iarg_83_tvalid = ap_tvalid[83];
            assign ap_axis_iarg_83_tkeep = ap_tkeep[83][S_AXIS_IARG_83_WIDTH/8-1:0];
            assign ap_axis_iarg_83_tstrb = ap_tstrb[83][S_AXIS_IARG_83_WIDTH/8-1:0];
            assign ap_axis_iarg_83_tdata = ap_tdata[83][S_AXIS_IARG_83_WIDTH-1:0];
            assign ap_tready[83] = ap_axis_iarg_83_tready;
        end
        if(C_NUM_INPUT_AXISs > 84) begin
            assign axis_clk[84] = s_axis_iarg_84_aclk;
            assign axis_rst[84] = s_axis_iarg_84_aresetn;
            assign dm_tlast[84] = s_axis_iarg_84_tlast;
            assign dm_tvalid[84] = s_axis_iarg_84_tvalid;
            assign dm_tkeep[84][S_AXIS_IARG_84_DMWIDTH/8-1:0] = s_axis_iarg_84_tkeep;
            assign dm_tstrb[84][S_AXIS_IARG_84_DMWIDTH/8-1:0] = s_axis_iarg_84_tstrb;
            assign dm_tdata[84][S_AXIS_IARG_84_DMWIDTH-1:0] = s_axis_iarg_84_tdata;
            assign s_axis_iarg_84_tready = dm_tready[84];
            assign ap_axis_iarg_84_tlast = ap_tlast[84];
            assign ap_axis_iarg_84_tvalid = ap_tvalid[84];
            assign ap_axis_iarg_84_tkeep = ap_tkeep[84][S_AXIS_IARG_84_WIDTH/8-1:0];
            assign ap_axis_iarg_84_tstrb = ap_tstrb[84][S_AXIS_IARG_84_WIDTH/8-1:0];
            assign ap_axis_iarg_84_tdata = ap_tdata[84][S_AXIS_IARG_84_WIDTH-1:0];
            assign ap_tready[84] = ap_axis_iarg_84_tready;
        end
        if(C_NUM_INPUT_AXISs > 85) begin
            assign axis_clk[85] = s_axis_iarg_85_aclk;
            assign axis_rst[85] = s_axis_iarg_85_aresetn;
            assign dm_tlast[85] = s_axis_iarg_85_tlast;
            assign dm_tvalid[85] = s_axis_iarg_85_tvalid;
            assign dm_tkeep[85][S_AXIS_IARG_85_DMWIDTH/8-1:0] = s_axis_iarg_85_tkeep;
            assign dm_tstrb[85][S_AXIS_IARG_85_DMWIDTH/8-1:0] = s_axis_iarg_85_tstrb;
            assign dm_tdata[85][S_AXIS_IARG_85_DMWIDTH-1:0] = s_axis_iarg_85_tdata;
            assign s_axis_iarg_85_tready = dm_tready[85];
            assign ap_axis_iarg_85_tlast = ap_tlast[85];
            assign ap_axis_iarg_85_tvalid = ap_tvalid[85];
            assign ap_axis_iarg_85_tkeep = ap_tkeep[85][S_AXIS_IARG_85_WIDTH/8-1:0];
            assign ap_axis_iarg_85_tstrb = ap_tstrb[85][S_AXIS_IARG_85_WIDTH/8-1:0];
            assign ap_axis_iarg_85_tdata = ap_tdata[85][S_AXIS_IARG_85_WIDTH-1:0];
            assign ap_tready[85] = ap_axis_iarg_85_tready;
        end
        if(C_NUM_INPUT_AXISs > 86) begin
            assign axis_clk[86] = s_axis_iarg_86_aclk;
            assign axis_rst[86] = s_axis_iarg_86_aresetn;
            assign dm_tlast[86] = s_axis_iarg_86_tlast;
            assign dm_tvalid[86] = s_axis_iarg_86_tvalid;
            assign dm_tkeep[86][S_AXIS_IARG_86_DMWIDTH/8-1:0] = s_axis_iarg_86_tkeep;
            assign dm_tstrb[86][S_AXIS_IARG_86_DMWIDTH/8-1:0] = s_axis_iarg_86_tstrb;
            assign dm_tdata[86][S_AXIS_IARG_86_DMWIDTH-1:0] = s_axis_iarg_86_tdata;
            assign s_axis_iarg_86_tready = dm_tready[86];
            assign ap_axis_iarg_86_tlast = ap_tlast[86];
            assign ap_axis_iarg_86_tvalid = ap_tvalid[86];
            assign ap_axis_iarg_86_tkeep = ap_tkeep[86][S_AXIS_IARG_86_WIDTH/8-1:0];
            assign ap_axis_iarg_86_tstrb = ap_tstrb[86][S_AXIS_IARG_86_WIDTH/8-1:0];
            assign ap_axis_iarg_86_tdata = ap_tdata[86][S_AXIS_IARG_86_WIDTH-1:0];
            assign ap_tready[86] = ap_axis_iarg_86_tready;
        end
        if(C_NUM_INPUT_AXISs > 87) begin
            assign axis_clk[87] = s_axis_iarg_87_aclk;
            assign axis_rst[87] = s_axis_iarg_87_aresetn;
            assign dm_tlast[87] = s_axis_iarg_87_tlast;
            assign dm_tvalid[87] = s_axis_iarg_87_tvalid;
            assign dm_tkeep[87][S_AXIS_IARG_87_DMWIDTH/8-1:0] = s_axis_iarg_87_tkeep;
            assign dm_tstrb[87][S_AXIS_IARG_87_DMWIDTH/8-1:0] = s_axis_iarg_87_tstrb;
            assign dm_tdata[87][S_AXIS_IARG_87_DMWIDTH-1:0] = s_axis_iarg_87_tdata;
            assign s_axis_iarg_87_tready = dm_tready[87];
            assign ap_axis_iarg_87_tlast = ap_tlast[87];
            assign ap_axis_iarg_87_tvalid = ap_tvalid[87];
            assign ap_axis_iarg_87_tkeep = ap_tkeep[87][S_AXIS_IARG_87_WIDTH/8-1:0];
            assign ap_axis_iarg_87_tstrb = ap_tstrb[87][S_AXIS_IARG_87_WIDTH/8-1:0];
            assign ap_axis_iarg_87_tdata = ap_tdata[87][S_AXIS_IARG_87_WIDTH-1:0];
            assign ap_tready[87] = ap_axis_iarg_87_tready;
        end
        if(C_NUM_INPUT_AXISs > 88) begin
            assign axis_clk[88] = s_axis_iarg_88_aclk;
            assign axis_rst[88] = s_axis_iarg_88_aresetn;
            assign dm_tlast[88] = s_axis_iarg_88_tlast;
            assign dm_tvalid[88] = s_axis_iarg_88_tvalid;
            assign dm_tkeep[88][S_AXIS_IARG_88_DMWIDTH/8-1:0] = s_axis_iarg_88_tkeep;
            assign dm_tstrb[88][S_AXIS_IARG_88_DMWIDTH/8-1:0] = s_axis_iarg_88_tstrb;
            assign dm_tdata[88][S_AXIS_IARG_88_DMWIDTH-1:0] = s_axis_iarg_88_tdata;
            assign s_axis_iarg_88_tready = dm_tready[88];
            assign ap_axis_iarg_88_tlast = ap_tlast[88];
            assign ap_axis_iarg_88_tvalid = ap_tvalid[88];
            assign ap_axis_iarg_88_tkeep = ap_tkeep[88][S_AXIS_IARG_88_WIDTH/8-1:0];
            assign ap_axis_iarg_88_tstrb = ap_tstrb[88][S_AXIS_IARG_88_WIDTH/8-1:0];
            assign ap_axis_iarg_88_tdata = ap_tdata[88][S_AXIS_IARG_88_WIDTH-1:0];
            assign ap_tready[88] = ap_axis_iarg_88_tready;
        end
        if(C_NUM_INPUT_AXISs > 89) begin
            assign axis_clk[89] = s_axis_iarg_89_aclk;
            assign axis_rst[89] = s_axis_iarg_89_aresetn;
            assign dm_tlast[89] = s_axis_iarg_89_tlast;
            assign dm_tvalid[89] = s_axis_iarg_89_tvalid;
            assign dm_tkeep[89][S_AXIS_IARG_89_DMWIDTH/8-1:0] = s_axis_iarg_89_tkeep;
            assign dm_tstrb[89][S_AXIS_IARG_89_DMWIDTH/8-1:0] = s_axis_iarg_89_tstrb;
            assign dm_tdata[89][S_AXIS_IARG_89_DMWIDTH-1:0] = s_axis_iarg_89_tdata;
            assign s_axis_iarg_89_tready = dm_tready[89];
            assign ap_axis_iarg_89_tlast = ap_tlast[89];
            assign ap_axis_iarg_89_tvalid = ap_tvalid[89];
            assign ap_axis_iarg_89_tkeep = ap_tkeep[89][S_AXIS_IARG_89_WIDTH/8-1:0];
            assign ap_axis_iarg_89_tstrb = ap_tstrb[89][S_AXIS_IARG_89_WIDTH/8-1:0];
            assign ap_axis_iarg_89_tdata = ap_tdata[89][S_AXIS_IARG_89_WIDTH-1:0];
            assign ap_tready[89] = ap_axis_iarg_89_tready;
        end
        if(C_NUM_INPUT_AXISs > 90) begin
            assign axis_clk[90] = s_axis_iarg_90_aclk;
            assign axis_rst[90] = s_axis_iarg_90_aresetn;
            assign dm_tlast[90] = s_axis_iarg_90_tlast;
            assign dm_tvalid[90] = s_axis_iarg_90_tvalid;
            assign dm_tkeep[90][S_AXIS_IARG_90_DMWIDTH/8-1:0] = s_axis_iarg_90_tkeep;
            assign dm_tstrb[90][S_AXIS_IARG_90_DMWIDTH/8-1:0] = s_axis_iarg_90_tstrb;
            assign dm_tdata[90][S_AXIS_IARG_90_DMWIDTH-1:0] = s_axis_iarg_90_tdata;
            assign s_axis_iarg_90_tready = dm_tready[90];
            assign ap_axis_iarg_90_tlast = ap_tlast[90];
            assign ap_axis_iarg_90_tvalid = ap_tvalid[90];
            assign ap_axis_iarg_90_tkeep = ap_tkeep[90][S_AXIS_IARG_90_WIDTH/8-1:0];
            assign ap_axis_iarg_90_tstrb = ap_tstrb[90][S_AXIS_IARG_90_WIDTH/8-1:0];
            assign ap_axis_iarg_90_tdata = ap_tdata[90][S_AXIS_IARG_90_WIDTH-1:0];
            assign ap_tready[90] = ap_axis_iarg_90_tready;
        end
        if(C_NUM_INPUT_AXISs > 91) begin
            assign axis_clk[91] = s_axis_iarg_91_aclk;
            assign axis_rst[91] = s_axis_iarg_91_aresetn;
            assign dm_tlast[91] = s_axis_iarg_91_tlast;
            assign dm_tvalid[91] = s_axis_iarg_91_tvalid;
            assign dm_tkeep[91][S_AXIS_IARG_91_DMWIDTH/8-1:0] = s_axis_iarg_91_tkeep;
            assign dm_tstrb[91][S_AXIS_IARG_91_DMWIDTH/8-1:0] = s_axis_iarg_91_tstrb;
            assign dm_tdata[91][S_AXIS_IARG_91_DMWIDTH-1:0] = s_axis_iarg_91_tdata;
            assign s_axis_iarg_91_tready = dm_tready[91];
            assign ap_axis_iarg_91_tlast = ap_tlast[91];
            assign ap_axis_iarg_91_tvalid = ap_tvalid[91];
            assign ap_axis_iarg_91_tkeep = ap_tkeep[91][S_AXIS_IARG_91_WIDTH/8-1:0];
            assign ap_axis_iarg_91_tstrb = ap_tstrb[91][S_AXIS_IARG_91_WIDTH/8-1:0];
            assign ap_axis_iarg_91_tdata = ap_tdata[91][S_AXIS_IARG_91_WIDTH-1:0];
            assign ap_tready[91] = ap_axis_iarg_91_tready;
        end
        if(C_NUM_INPUT_AXISs > 92) begin
            assign axis_clk[92] = s_axis_iarg_92_aclk;
            assign axis_rst[92] = s_axis_iarg_92_aresetn;
            assign dm_tlast[92] = s_axis_iarg_92_tlast;
            assign dm_tvalid[92] = s_axis_iarg_92_tvalid;
            assign dm_tkeep[92][S_AXIS_IARG_92_DMWIDTH/8-1:0] = s_axis_iarg_92_tkeep;
            assign dm_tstrb[92][S_AXIS_IARG_92_DMWIDTH/8-1:0] = s_axis_iarg_92_tstrb;
            assign dm_tdata[92][S_AXIS_IARG_92_DMWIDTH-1:0] = s_axis_iarg_92_tdata;
            assign s_axis_iarg_92_tready = dm_tready[92];
            assign ap_axis_iarg_92_tlast = ap_tlast[92];
            assign ap_axis_iarg_92_tvalid = ap_tvalid[92];
            assign ap_axis_iarg_92_tkeep = ap_tkeep[92][S_AXIS_IARG_92_WIDTH/8-1:0];
            assign ap_axis_iarg_92_tstrb = ap_tstrb[92][S_AXIS_IARG_92_WIDTH/8-1:0];
            assign ap_axis_iarg_92_tdata = ap_tdata[92][S_AXIS_IARG_92_WIDTH-1:0];
            assign ap_tready[92] = ap_axis_iarg_92_tready;
        end
        if(C_NUM_INPUT_AXISs > 93) begin
            assign axis_clk[93] = s_axis_iarg_93_aclk;
            assign axis_rst[93] = s_axis_iarg_93_aresetn;
            assign dm_tlast[93] = s_axis_iarg_93_tlast;
            assign dm_tvalid[93] = s_axis_iarg_93_tvalid;
            assign dm_tkeep[93][S_AXIS_IARG_93_DMWIDTH/8-1:0] = s_axis_iarg_93_tkeep;
            assign dm_tstrb[93][S_AXIS_IARG_93_DMWIDTH/8-1:0] = s_axis_iarg_93_tstrb;
            assign dm_tdata[93][S_AXIS_IARG_93_DMWIDTH-1:0] = s_axis_iarg_93_tdata;
            assign s_axis_iarg_93_tready = dm_tready[93];
            assign ap_axis_iarg_93_tlast = ap_tlast[93];
            assign ap_axis_iarg_93_tvalid = ap_tvalid[93];
            assign ap_axis_iarg_93_tkeep = ap_tkeep[93][S_AXIS_IARG_93_WIDTH/8-1:0];
            assign ap_axis_iarg_93_tstrb = ap_tstrb[93][S_AXIS_IARG_93_WIDTH/8-1:0];
            assign ap_axis_iarg_93_tdata = ap_tdata[93][S_AXIS_IARG_93_WIDTH-1:0];
            assign ap_tready[93] = ap_axis_iarg_93_tready;
        end
        if(C_NUM_INPUT_AXISs > 94) begin
            assign axis_clk[94] = s_axis_iarg_94_aclk;
            assign axis_rst[94] = s_axis_iarg_94_aresetn;
            assign dm_tlast[94] = s_axis_iarg_94_tlast;
            assign dm_tvalid[94] = s_axis_iarg_94_tvalid;
            assign dm_tkeep[94][S_AXIS_IARG_94_DMWIDTH/8-1:0] = s_axis_iarg_94_tkeep;
            assign dm_tstrb[94][S_AXIS_IARG_94_DMWIDTH/8-1:0] = s_axis_iarg_94_tstrb;
            assign dm_tdata[94][S_AXIS_IARG_94_DMWIDTH-1:0] = s_axis_iarg_94_tdata;
            assign s_axis_iarg_94_tready = dm_tready[94];
            assign ap_axis_iarg_94_tlast = ap_tlast[94];
            assign ap_axis_iarg_94_tvalid = ap_tvalid[94];
            assign ap_axis_iarg_94_tkeep = ap_tkeep[94][S_AXIS_IARG_94_WIDTH/8-1:0];
            assign ap_axis_iarg_94_tstrb = ap_tstrb[94][S_AXIS_IARG_94_WIDTH/8-1:0];
            assign ap_axis_iarg_94_tdata = ap_tdata[94][S_AXIS_IARG_94_WIDTH-1:0];
            assign ap_tready[94] = ap_axis_iarg_94_tready;
        end
        if(C_NUM_INPUT_AXISs > 95) begin
            assign axis_clk[95] = s_axis_iarg_95_aclk;
            assign axis_rst[95] = s_axis_iarg_95_aresetn;
            assign dm_tlast[95] = s_axis_iarg_95_tlast;
            assign dm_tvalid[95] = s_axis_iarg_95_tvalid;
            assign dm_tkeep[95][S_AXIS_IARG_95_DMWIDTH/8-1:0] = s_axis_iarg_95_tkeep;
            assign dm_tstrb[95][S_AXIS_IARG_95_DMWIDTH/8-1:0] = s_axis_iarg_95_tstrb;
            assign dm_tdata[95][S_AXIS_IARG_95_DMWIDTH-1:0] = s_axis_iarg_95_tdata;
            assign s_axis_iarg_95_tready = dm_tready[95];
            assign ap_axis_iarg_95_tlast = ap_tlast[95];
            assign ap_axis_iarg_95_tvalid = ap_tvalid[95];
            assign ap_axis_iarg_95_tkeep = ap_tkeep[95][S_AXIS_IARG_95_WIDTH/8-1:0];
            assign ap_axis_iarg_95_tstrb = ap_tstrb[95][S_AXIS_IARG_95_WIDTH/8-1:0];
            assign ap_axis_iarg_95_tdata = ap_tdata[95][S_AXIS_IARG_95_WIDTH-1:0];
            assign ap_tready[95] = ap_axis_iarg_95_tready;
        end
        if(C_NUM_INPUT_AXISs > 96) begin
            assign axis_clk[96] = s_axis_iarg_96_aclk;
            assign axis_rst[96] = s_axis_iarg_96_aresetn;
            assign dm_tlast[96] = s_axis_iarg_96_tlast;
            assign dm_tvalid[96] = s_axis_iarg_96_tvalid;
            assign dm_tkeep[96][S_AXIS_IARG_96_DMWIDTH/8-1:0] = s_axis_iarg_96_tkeep;
            assign dm_tstrb[96][S_AXIS_IARG_96_DMWIDTH/8-1:0] = s_axis_iarg_96_tstrb;
            assign dm_tdata[96][S_AXIS_IARG_96_DMWIDTH-1:0] = s_axis_iarg_96_tdata;
            assign s_axis_iarg_96_tready = dm_tready[96];
            assign ap_axis_iarg_96_tlast = ap_tlast[96];
            assign ap_axis_iarg_96_tvalid = ap_tvalid[96];
            assign ap_axis_iarg_96_tkeep = ap_tkeep[96][S_AXIS_IARG_96_WIDTH/8-1:0];
            assign ap_axis_iarg_96_tstrb = ap_tstrb[96][S_AXIS_IARG_96_WIDTH/8-1:0];
            assign ap_axis_iarg_96_tdata = ap_tdata[96][S_AXIS_IARG_96_WIDTH-1:0];
            assign ap_tready[96] = ap_axis_iarg_96_tready;
        end
        if(C_NUM_INPUT_AXISs > 97) begin
            assign axis_clk[97] = s_axis_iarg_97_aclk;
            assign axis_rst[97] = s_axis_iarg_97_aresetn;
            assign dm_tlast[97] = s_axis_iarg_97_tlast;
            assign dm_tvalid[97] = s_axis_iarg_97_tvalid;
            assign dm_tkeep[97][S_AXIS_IARG_97_DMWIDTH/8-1:0] = s_axis_iarg_97_tkeep;
            assign dm_tstrb[97][S_AXIS_IARG_97_DMWIDTH/8-1:0] = s_axis_iarg_97_tstrb;
            assign dm_tdata[97][S_AXIS_IARG_97_DMWIDTH-1:0] = s_axis_iarg_97_tdata;
            assign s_axis_iarg_97_tready = dm_tready[97];
            assign ap_axis_iarg_97_tlast = ap_tlast[97];
            assign ap_axis_iarg_97_tvalid = ap_tvalid[97];
            assign ap_axis_iarg_97_tkeep = ap_tkeep[97][S_AXIS_IARG_97_WIDTH/8-1:0];
            assign ap_axis_iarg_97_tstrb = ap_tstrb[97][S_AXIS_IARG_97_WIDTH/8-1:0];
            assign ap_axis_iarg_97_tdata = ap_tdata[97][S_AXIS_IARG_97_WIDTH-1:0];
            assign ap_tready[97] = ap_axis_iarg_97_tready;
        end
        if(C_NUM_INPUT_AXISs > 98) begin
            assign axis_clk[98] = s_axis_iarg_98_aclk;
            assign axis_rst[98] = s_axis_iarg_98_aresetn;
            assign dm_tlast[98] = s_axis_iarg_98_tlast;
            assign dm_tvalid[98] = s_axis_iarg_98_tvalid;
            assign dm_tkeep[98][S_AXIS_IARG_98_DMWIDTH/8-1:0] = s_axis_iarg_98_tkeep;
            assign dm_tstrb[98][S_AXIS_IARG_98_DMWIDTH/8-1:0] = s_axis_iarg_98_tstrb;
            assign dm_tdata[98][S_AXIS_IARG_98_DMWIDTH-1:0] = s_axis_iarg_98_tdata;
            assign s_axis_iarg_98_tready = dm_tready[98];
            assign ap_axis_iarg_98_tlast = ap_tlast[98];
            assign ap_axis_iarg_98_tvalid = ap_tvalid[98];
            assign ap_axis_iarg_98_tkeep = ap_tkeep[98][S_AXIS_IARG_98_WIDTH/8-1:0];
            assign ap_axis_iarg_98_tstrb = ap_tstrb[98][S_AXIS_IARG_98_WIDTH/8-1:0];
            assign ap_axis_iarg_98_tdata = ap_tdata[98][S_AXIS_IARG_98_WIDTH-1:0];
            assign ap_tready[98] = ap_axis_iarg_98_tready;
        end
        if(C_NUM_INPUT_AXISs > 99) begin
            assign axis_clk[99] = s_axis_iarg_99_aclk;
            assign axis_rst[99] = s_axis_iarg_99_aresetn;
            assign dm_tlast[99] = s_axis_iarg_99_tlast;
            assign dm_tvalid[99] = s_axis_iarg_99_tvalid;
            assign dm_tkeep[99][S_AXIS_IARG_99_DMWIDTH/8-1:0] = s_axis_iarg_99_tkeep;
            assign dm_tstrb[99][S_AXIS_IARG_99_DMWIDTH/8-1:0] = s_axis_iarg_99_tstrb;
            assign dm_tdata[99][S_AXIS_IARG_99_DMWIDTH-1:0] = s_axis_iarg_99_tdata;
            assign s_axis_iarg_99_tready = dm_tready[99];
            assign ap_axis_iarg_99_tlast = ap_tlast[99];
            assign ap_axis_iarg_99_tvalid = ap_tvalid[99];
            assign ap_axis_iarg_99_tkeep = ap_tkeep[99][S_AXIS_IARG_99_WIDTH/8-1:0];
            assign ap_axis_iarg_99_tstrb = ap_tstrb[99][S_AXIS_IARG_99_WIDTH/8-1:0];
            assign ap_axis_iarg_99_tdata = ap_tdata[99][S_AXIS_IARG_99_WIDTH-1:0];
            assign ap_tready[99] = ap_axis_iarg_99_tready;
        end
        if(C_NUM_INPUT_AXISs > 100) begin
            assign axis_clk[100] = s_axis_iarg_100_aclk;
            assign axis_rst[100] = s_axis_iarg_100_aresetn;
            assign dm_tlast[100] = s_axis_iarg_100_tlast;
            assign dm_tvalid[100] = s_axis_iarg_100_tvalid;
            assign dm_tkeep[100][S_AXIS_IARG_100_DMWIDTH/8-1:0] = s_axis_iarg_100_tkeep;
            assign dm_tstrb[100][S_AXIS_IARG_100_DMWIDTH/8-1:0] = s_axis_iarg_100_tstrb;
            assign dm_tdata[100][S_AXIS_IARG_100_DMWIDTH-1:0] = s_axis_iarg_100_tdata;
            assign s_axis_iarg_100_tready = dm_tready[100];
            assign ap_axis_iarg_100_tlast = ap_tlast[100];
            assign ap_axis_iarg_100_tvalid = ap_tvalid[100];
            assign ap_axis_iarg_100_tkeep = ap_tkeep[100][S_AXIS_IARG_100_WIDTH/8-1:0];
            assign ap_axis_iarg_100_tstrb = ap_tstrb[100][S_AXIS_IARG_100_WIDTH/8-1:0];
            assign ap_axis_iarg_100_tdata = ap_tdata[100][S_AXIS_IARG_100_WIDTH-1:0];
            assign ap_tready[100] = ap_axis_iarg_100_tready;
        end
        if(C_NUM_INPUT_AXISs > 101) begin
            assign axis_clk[101] = s_axis_iarg_101_aclk;
            assign axis_rst[101] = s_axis_iarg_101_aresetn;
            assign dm_tlast[101] = s_axis_iarg_101_tlast;
            assign dm_tvalid[101] = s_axis_iarg_101_tvalid;
            assign dm_tkeep[101][S_AXIS_IARG_101_DMWIDTH/8-1:0] = s_axis_iarg_101_tkeep;
            assign dm_tstrb[101][S_AXIS_IARG_101_DMWIDTH/8-1:0] = s_axis_iarg_101_tstrb;
            assign dm_tdata[101][S_AXIS_IARG_101_DMWIDTH-1:0] = s_axis_iarg_101_tdata;
            assign s_axis_iarg_101_tready = dm_tready[101];
            assign ap_axis_iarg_101_tlast = ap_tlast[101];
            assign ap_axis_iarg_101_tvalid = ap_tvalid[101];
            assign ap_axis_iarg_101_tkeep = ap_tkeep[101][S_AXIS_IARG_101_WIDTH/8-1:0];
            assign ap_axis_iarg_101_tstrb = ap_tstrb[101][S_AXIS_IARG_101_WIDTH/8-1:0];
            assign ap_axis_iarg_101_tdata = ap_tdata[101][S_AXIS_IARG_101_WIDTH-1:0];
            assign ap_tready[101] = ap_axis_iarg_101_tready;
        end
        if(C_NUM_INPUT_AXISs > 102) begin
            assign axis_clk[102] = s_axis_iarg_102_aclk;
            assign axis_rst[102] = s_axis_iarg_102_aresetn;
            assign dm_tlast[102] = s_axis_iarg_102_tlast;
            assign dm_tvalid[102] = s_axis_iarg_102_tvalid;
            assign dm_tkeep[102][S_AXIS_IARG_102_DMWIDTH/8-1:0] = s_axis_iarg_102_tkeep;
            assign dm_tstrb[102][S_AXIS_IARG_102_DMWIDTH/8-1:0] = s_axis_iarg_102_tstrb;
            assign dm_tdata[102][S_AXIS_IARG_102_DMWIDTH-1:0] = s_axis_iarg_102_tdata;
            assign s_axis_iarg_102_tready = dm_tready[102];
            assign ap_axis_iarg_102_tlast = ap_tlast[102];
            assign ap_axis_iarg_102_tvalid = ap_tvalid[102];
            assign ap_axis_iarg_102_tkeep = ap_tkeep[102][S_AXIS_IARG_102_WIDTH/8-1:0];
            assign ap_axis_iarg_102_tstrb = ap_tstrb[102][S_AXIS_IARG_102_WIDTH/8-1:0];
            assign ap_axis_iarg_102_tdata = ap_tdata[102][S_AXIS_IARG_102_WIDTH-1:0];
            assign ap_tready[102] = ap_axis_iarg_102_tready;
        end
        if(C_NUM_INPUT_AXISs > 103) begin
            assign axis_clk[103] = s_axis_iarg_103_aclk;
            assign axis_rst[103] = s_axis_iarg_103_aresetn;
            assign dm_tlast[103] = s_axis_iarg_103_tlast;
            assign dm_tvalid[103] = s_axis_iarg_103_tvalid;
            assign dm_tkeep[103][S_AXIS_IARG_103_DMWIDTH/8-1:0] = s_axis_iarg_103_tkeep;
            assign dm_tstrb[103][S_AXIS_IARG_103_DMWIDTH/8-1:0] = s_axis_iarg_103_tstrb;
            assign dm_tdata[103][S_AXIS_IARG_103_DMWIDTH-1:0] = s_axis_iarg_103_tdata;
            assign s_axis_iarg_103_tready = dm_tready[103];
            assign ap_axis_iarg_103_tlast = ap_tlast[103];
            assign ap_axis_iarg_103_tvalid = ap_tvalid[103];
            assign ap_axis_iarg_103_tkeep = ap_tkeep[103][S_AXIS_IARG_103_WIDTH/8-1:0];
            assign ap_axis_iarg_103_tstrb = ap_tstrb[103][S_AXIS_IARG_103_WIDTH/8-1:0];
            assign ap_axis_iarg_103_tdata = ap_tdata[103][S_AXIS_IARG_103_WIDTH-1:0];
            assign ap_tready[103] = ap_axis_iarg_103_tready;
        end
        if(C_NUM_INPUT_AXISs > 104) begin
            assign axis_clk[104] = s_axis_iarg_104_aclk;
            assign axis_rst[104] = s_axis_iarg_104_aresetn;
            assign dm_tlast[104] = s_axis_iarg_104_tlast;
            assign dm_tvalid[104] = s_axis_iarg_104_tvalid;
            assign dm_tkeep[104][S_AXIS_IARG_104_DMWIDTH/8-1:0] = s_axis_iarg_104_tkeep;
            assign dm_tstrb[104][S_AXIS_IARG_104_DMWIDTH/8-1:0] = s_axis_iarg_104_tstrb;
            assign dm_tdata[104][S_AXIS_IARG_104_DMWIDTH-1:0] = s_axis_iarg_104_tdata;
            assign s_axis_iarg_104_tready = dm_tready[104];
            assign ap_axis_iarg_104_tlast = ap_tlast[104];
            assign ap_axis_iarg_104_tvalid = ap_tvalid[104];
            assign ap_axis_iarg_104_tkeep = ap_tkeep[104][S_AXIS_IARG_104_WIDTH/8-1:0];
            assign ap_axis_iarg_104_tstrb = ap_tstrb[104][S_AXIS_IARG_104_WIDTH/8-1:0];
            assign ap_axis_iarg_104_tdata = ap_tdata[104][S_AXIS_IARG_104_WIDTH-1:0];
            assign ap_tready[104] = ap_axis_iarg_104_tready;
        end
        if(C_NUM_INPUT_AXISs > 105) begin
            assign axis_clk[105] = s_axis_iarg_105_aclk;
            assign axis_rst[105] = s_axis_iarg_105_aresetn;
            assign dm_tlast[105] = s_axis_iarg_105_tlast;
            assign dm_tvalid[105] = s_axis_iarg_105_tvalid;
            assign dm_tkeep[105][S_AXIS_IARG_105_DMWIDTH/8-1:0] = s_axis_iarg_105_tkeep;
            assign dm_tstrb[105][S_AXIS_IARG_105_DMWIDTH/8-1:0] = s_axis_iarg_105_tstrb;
            assign dm_tdata[105][S_AXIS_IARG_105_DMWIDTH-1:0] = s_axis_iarg_105_tdata;
            assign s_axis_iarg_105_tready = dm_tready[105];
            assign ap_axis_iarg_105_tlast = ap_tlast[105];
            assign ap_axis_iarg_105_tvalid = ap_tvalid[105];
            assign ap_axis_iarg_105_tkeep = ap_tkeep[105][S_AXIS_IARG_105_WIDTH/8-1:0];
            assign ap_axis_iarg_105_tstrb = ap_tstrb[105][S_AXIS_IARG_105_WIDTH/8-1:0];
            assign ap_axis_iarg_105_tdata = ap_tdata[105][S_AXIS_IARG_105_WIDTH-1:0];
            assign ap_tready[105] = ap_axis_iarg_105_tready;
        end
        if(C_NUM_INPUT_AXISs > 106) begin
            assign axis_clk[106] = s_axis_iarg_106_aclk;
            assign axis_rst[106] = s_axis_iarg_106_aresetn;
            assign dm_tlast[106] = s_axis_iarg_106_tlast;
            assign dm_tvalid[106] = s_axis_iarg_106_tvalid;
            assign dm_tkeep[106][S_AXIS_IARG_106_DMWIDTH/8-1:0] = s_axis_iarg_106_tkeep;
            assign dm_tstrb[106][S_AXIS_IARG_106_DMWIDTH/8-1:0] = s_axis_iarg_106_tstrb;
            assign dm_tdata[106][S_AXIS_IARG_106_DMWIDTH-1:0] = s_axis_iarg_106_tdata;
            assign s_axis_iarg_106_tready = dm_tready[106];
            assign ap_axis_iarg_106_tlast = ap_tlast[106];
            assign ap_axis_iarg_106_tvalid = ap_tvalid[106];
            assign ap_axis_iarg_106_tkeep = ap_tkeep[106][S_AXIS_IARG_106_WIDTH/8-1:0];
            assign ap_axis_iarg_106_tstrb = ap_tstrb[106][S_AXIS_IARG_106_WIDTH/8-1:0];
            assign ap_axis_iarg_106_tdata = ap_tdata[106][S_AXIS_IARG_106_WIDTH-1:0];
            assign ap_tready[106] = ap_axis_iarg_106_tready;
        end
        if(C_NUM_INPUT_AXISs > 107) begin
            assign axis_clk[107] = s_axis_iarg_107_aclk;
            assign axis_rst[107] = s_axis_iarg_107_aresetn;
            assign dm_tlast[107] = s_axis_iarg_107_tlast;
            assign dm_tvalid[107] = s_axis_iarg_107_tvalid;
            assign dm_tkeep[107][S_AXIS_IARG_107_DMWIDTH/8-1:0] = s_axis_iarg_107_tkeep;
            assign dm_tstrb[107][S_AXIS_IARG_107_DMWIDTH/8-1:0] = s_axis_iarg_107_tstrb;
            assign dm_tdata[107][S_AXIS_IARG_107_DMWIDTH-1:0] = s_axis_iarg_107_tdata;
            assign s_axis_iarg_107_tready = dm_tready[107];
            assign ap_axis_iarg_107_tlast = ap_tlast[107];
            assign ap_axis_iarg_107_tvalid = ap_tvalid[107];
            assign ap_axis_iarg_107_tkeep = ap_tkeep[107][S_AXIS_IARG_107_WIDTH/8-1:0];
            assign ap_axis_iarg_107_tstrb = ap_tstrb[107][S_AXIS_IARG_107_WIDTH/8-1:0];
            assign ap_axis_iarg_107_tdata = ap_tdata[107][S_AXIS_IARG_107_WIDTH-1:0];
            assign ap_tready[107] = ap_axis_iarg_107_tready;
        end
        if(C_NUM_INPUT_AXISs > 108) begin
            assign axis_clk[108] = s_axis_iarg_108_aclk;
            assign axis_rst[108] = s_axis_iarg_108_aresetn;
            assign dm_tlast[108] = s_axis_iarg_108_tlast;
            assign dm_tvalid[108] = s_axis_iarg_108_tvalid;
            assign dm_tkeep[108][S_AXIS_IARG_108_DMWIDTH/8-1:0] = s_axis_iarg_108_tkeep;
            assign dm_tstrb[108][S_AXIS_IARG_108_DMWIDTH/8-1:0] = s_axis_iarg_108_tstrb;
            assign dm_tdata[108][S_AXIS_IARG_108_DMWIDTH-1:0] = s_axis_iarg_108_tdata;
            assign s_axis_iarg_108_tready = dm_tready[108];
            assign ap_axis_iarg_108_tlast = ap_tlast[108];
            assign ap_axis_iarg_108_tvalid = ap_tvalid[108];
            assign ap_axis_iarg_108_tkeep = ap_tkeep[108][S_AXIS_IARG_108_WIDTH/8-1:0];
            assign ap_axis_iarg_108_tstrb = ap_tstrb[108][S_AXIS_IARG_108_WIDTH/8-1:0];
            assign ap_axis_iarg_108_tdata = ap_tdata[108][S_AXIS_IARG_108_WIDTH-1:0];
            assign ap_tready[108] = ap_axis_iarg_108_tready;
        end
        if(C_NUM_INPUT_AXISs > 109) begin
            assign axis_clk[109] = s_axis_iarg_109_aclk;
            assign axis_rst[109] = s_axis_iarg_109_aresetn;
            assign dm_tlast[109] = s_axis_iarg_109_tlast;
            assign dm_tvalid[109] = s_axis_iarg_109_tvalid;
            assign dm_tkeep[109][S_AXIS_IARG_109_DMWIDTH/8-1:0] = s_axis_iarg_109_tkeep;
            assign dm_tstrb[109][S_AXIS_IARG_109_DMWIDTH/8-1:0] = s_axis_iarg_109_tstrb;
            assign dm_tdata[109][S_AXIS_IARG_109_DMWIDTH-1:0] = s_axis_iarg_109_tdata;
            assign s_axis_iarg_109_tready = dm_tready[109];
            assign ap_axis_iarg_109_tlast = ap_tlast[109];
            assign ap_axis_iarg_109_tvalid = ap_tvalid[109];
            assign ap_axis_iarg_109_tkeep = ap_tkeep[109][S_AXIS_IARG_109_WIDTH/8-1:0];
            assign ap_axis_iarg_109_tstrb = ap_tstrb[109][S_AXIS_IARG_109_WIDTH/8-1:0];
            assign ap_axis_iarg_109_tdata = ap_tdata[109][S_AXIS_IARG_109_WIDTH-1:0];
            assign ap_tready[109] = ap_axis_iarg_109_tready;
        end
        if(C_NUM_INPUT_AXISs > 110) begin
            assign axis_clk[110] = s_axis_iarg_110_aclk;
            assign axis_rst[110] = s_axis_iarg_110_aresetn;
            assign dm_tlast[110] = s_axis_iarg_110_tlast;
            assign dm_tvalid[110] = s_axis_iarg_110_tvalid;
            assign dm_tkeep[110][S_AXIS_IARG_110_DMWIDTH/8-1:0] = s_axis_iarg_110_tkeep;
            assign dm_tstrb[110][S_AXIS_IARG_110_DMWIDTH/8-1:0] = s_axis_iarg_110_tstrb;
            assign dm_tdata[110][S_AXIS_IARG_110_DMWIDTH-1:0] = s_axis_iarg_110_tdata;
            assign s_axis_iarg_110_tready = dm_tready[110];
            assign ap_axis_iarg_110_tlast = ap_tlast[110];
            assign ap_axis_iarg_110_tvalid = ap_tvalid[110];
            assign ap_axis_iarg_110_tkeep = ap_tkeep[110][S_AXIS_IARG_110_WIDTH/8-1:0];
            assign ap_axis_iarg_110_tstrb = ap_tstrb[110][S_AXIS_IARG_110_WIDTH/8-1:0];
            assign ap_axis_iarg_110_tdata = ap_tdata[110][S_AXIS_IARG_110_WIDTH-1:0];
            assign ap_tready[110] = ap_axis_iarg_110_tready;
        end
        if(C_NUM_INPUT_AXISs > 111) begin
            assign axis_clk[111] = s_axis_iarg_111_aclk;
            assign axis_rst[111] = s_axis_iarg_111_aresetn;
            assign dm_tlast[111] = s_axis_iarg_111_tlast;
            assign dm_tvalid[111] = s_axis_iarg_111_tvalid;
            assign dm_tkeep[111][S_AXIS_IARG_111_DMWIDTH/8-1:0] = s_axis_iarg_111_tkeep;
            assign dm_tstrb[111][S_AXIS_IARG_111_DMWIDTH/8-1:0] = s_axis_iarg_111_tstrb;
            assign dm_tdata[111][S_AXIS_IARG_111_DMWIDTH-1:0] = s_axis_iarg_111_tdata;
            assign s_axis_iarg_111_tready = dm_tready[111];
            assign ap_axis_iarg_111_tlast = ap_tlast[111];
            assign ap_axis_iarg_111_tvalid = ap_tvalid[111];
            assign ap_axis_iarg_111_tkeep = ap_tkeep[111][S_AXIS_IARG_111_WIDTH/8-1:0];
            assign ap_axis_iarg_111_tstrb = ap_tstrb[111][S_AXIS_IARG_111_WIDTH/8-1:0];
            assign ap_axis_iarg_111_tdata = ap_tdata[111][S_AXIS_IARG_111_WIDTH-1:0];
            assign ap_tready[111] = ap_axis_iarg_111_tready;
        end
        if(C_NUM_INPUT_AXISs > 112) begin
            assign axis_clk[112] = s_axis_iarg_112_aclk;
            assign axis_rst[112] = s_axis_iarg_112_aresetn;
            assign dm_tlast[112] = s_axis_iarg_112_tlast;
            assign dm_tvalid[112] = s_axis_iarg_112_tvalid;
            assign dm_tkeep[112][S_AXIS_IARG_112_DMWIDTH/8-1:0] = s_axis_iarg_112_tkeep;
            assign dm_tstrb[112][S_AXIS_IARG_112_DMWIDTH/8-1:0] = s_axis_iarg_112_tstrb;
            assign dm_tdata[112][S_AXIS_IARG_112_DMWIDTH-1:0] = s_axis_iarg_112_tdata;
            assign s_axis_iarg_112_tready = dm_tready[112];
            assign ap_axis_iarg_112_tlast = ap_tlast[112];
            assign ap_axis_iarg_112_tvalid = ap_tvalid[112];
            assign ap_axis_iarg_112_tkeep = ap_tkeep[112][S_AXIS_IARG_112_WIDTH/8-1:0];
            assign ap_axis_iarg_112_tstrb = ap_tstrb[112][S_AXIS_IARG_112_WIDTH/8-1:0];
            assign ap_axis_iarg_112_tdata = ap_tdata[112][S_AXIS_IARG_112_WIDTH-1:0];
            assign ap_tready[112] = ap_axis_iarg_112_tready;
        end
        if(C_NUM_INPUT_AXISs > 113) begin
            assign axis_clk[113] = s_axis_iarg_113_aclk;
            assign axis_rst[113] = s_axis_iarg_113_aresetn;
            assign dm_tlast[113] = s_axis_iarg_113_tlast;
            assign dm_tvalid[113] = s_axis_iarg_113_tvalid;
            assign dm_tkeep[113][S_AXIS_IARG_113_DMWIDTH/8-1:0] = s_axis_iarg_113_tkeep;
            assign dm_tstrb[113][S_AXIS_IARG_113_DMWIDTH/8-1:0] = s_axis_iarg_113_tstrb;
            assign dm_tdata[113][S_AXIS_IARG_113_DMWIDTH-1:0] = s_axis_iarg_113_tdata;
            assign s_axis_iarg_113_tready = dm_tready[113];
            assign ap_axis_iarg_113_tlast = ap_tlast[113];
            assign ap_axis_iarg_113_tvalid = ap_tvalid[113];
            assign ap_axis_iarg_113_tkeep = ap_tkeep[113][S_AXIS_IARG_113_WIDTH/8-1:0];
            assign ap_axis_iarg_113_tstrb = ap_tstrb[113][S_AXIS_IARG_113_WIDTH/8-1:0];
            assign ap_axis_iarg_113_tdata = ap_tdata[113][S_AXIS_IARG_113_WIDTH-1:0];
            assign ap_tready[113] = ap_axis_iarg_113_tready;
        end
        if(C_NUM_INPUT_AXISs > 114) begin
            assign axis_clk[114] = s_axis_iarg_114_aclk;
            assign axis_rst[114] = s_axis_iarg_114_aresetn;
            assign dm_tlast[114] = s_axis_iarg_114_tlast;
            assign dm_tvalid[114] = s_axis_iarg_114_tvalid;
            assign dm_tkeep[114][S_AXIS_IARG_114_DMWIDTH/8-1:0] = s_axis_iarg_114_tkeep;
            assign dm_tstrb[114][S_AXIS_IARG_114_DMWIDTH/8-1:0] = s_axis_iarg_114_tstrb;
            assign dm_tdata[114][S_AXIS_IARG_114_DMWIDTH-1:0] = s_axis_iarg_114_tdata;
            assign s_axis_iarg_114_tready = dm_tready[114];
            assign ap_axis_iarg_114_tlast = ap_tlast[114];
            assign ap_axis_iarg_114_tvalid = ap_tvalid[114];
            assign ap_axis_iarg_114_tkeep = ap_tkeep[114][S_AXIS_IARG_114_WIDTH/8-1:0];
            assign ap_axis_iarg_114_tstrb = ap_tstrb[114][S_AXIS_IARG_114_WIDTH/8-1:0];
            assign ap_axis_iarg_114_tdata = ap_tdata[114][S_AXIS_IARG_114_WIDTH-1:0];
            assign ap_tready[114] = ap_axis_iarg_114_tready;
        end
        if(C_NUM_INPUT_AXISs > 115) begin
            assign axis_clk[115] = s_axis_iarg_115_aclk;
            assign axis_rst[115] = s_axis_iarg_115_aresetn;
            assign dm_tlast[115] = s_axis_iarg_115_tlast;
            assign dm_tvalid[115] = s_axis_iarg_115_tvalid;
            assign dm_tkeep[115][S_AXIS_IARG_115_DMWIDTH/8-1:0] = s_axis_iarg_115_tkeep;
            assign dm_tstrb[115][S_AXIS_IARG_115_DMWIDTH/8-1:0] = s_axis_iarg_115_tstrb;
            assign dm_tdata[115][S_AXIS_IARG_115_DMWIDTH-1:0] = s_axis_iarg_115_tdata;
            assign s_axis_iarg_115_tready = dm_tready[115];
            assign ap_axis_iarg_115_tlast = ap_tlast[115];
            assign ap_axis_iarg_115_tvalid = ap_tvalid[115];
            assign ap_axis_iarg_115_tkeep = ap_tkeep[115][S_AXIS_IARG_115_WIDTH/8-1:0];
            assign ap_axis_iarg_115_tstrb = ap_tstrb[115][S_AXIS_IARG_115_WIDTH/8-1:0];
            assign ap_axis_iarg_115_tdata = ap_tdata[115][S_AXIS_IARG_115_WIDTH-1:0];
            assign ap_tready[115] = ap_axis_iarg_115_tready;
        end
        if(C_NUM_INPUT_AXISs > 116) begin
            assign axis_clk[116] = s_axis_iarg_116_aclk;
            assign axis_rst[116] = s_axis_iarg_116_aresetn;
            assign dm_tlast[116] = s_axis_iarg_116_tlast;
            assign dm_tvalid[116] = s_axis_iarg_116_tvalid;
            assign dm_tkeep[116][S_AXIS_IARG_116_DMWIDTH/8-1:0] = s_axis_iarg_116_tkeep;
            assign dm_tstrb[116][S_AXIS_IARG_116_DMWIDTH/8-1:0] = s_axis_iarg_116_tstrb;
            assign dm_tdata[116][S_AXIS_IARG_116_DMWIDTH-1:0] = s_axis_iarg_116_tdata;
            assign s_axis_iarg_116_tready = dm_tready[116];
            assign ap_axis_iarg_116_tlast = ap_tlast[116];
            assign ap_axis_iarg_116_tvalid = ap_tvalid[116];
            assign ap_axis_iarg_116_tkeep = ap_tkeep[116][S_AXIS_IARG_116_WIDTH/8-1:0];
            assign ap_axis_iarg_116_tstrb = ap_tstrb[116][S_AXIS_IARG_116_WIDTH/8-1:0];
            assign ap_axis_iarg_116_tdata = ap_tdata[116][S_AXIS_IARG_116_WIDTH-1:0];
            assign ap_tready[116] = ap_axis_iarg_116_tready;
        end
        if(C_NUM_INPUT_AXISs > 117) begin
            assign axis_clk[117] = s_axis_iarg_117_aclk;
            assign axis_rst[117] = s_axis_iarg_117_aresetn;
            assign dm_tlast[117] = s_axis_iarg_117_tlast;
            assign dm_tvalid[117] = s_axis_iarg_117_tvalid;
            assign dm_tkeep[117][S_AXIS_IARG_117_DMWIDTH/8-1:0] = s_axis_iarg_117_tkeep;
            assign dm_tstrb[117][S_AXIS_IARG_117_DMWIDTH/8-1:0] = s_axis_iarg_117_tstrb;
            assign dm_tdata[117][S_AXIS_IARG_117_DMWIDTH-1:0] = s_axis_iarg_117_tdata;
            assign s_axis_iarg_117_tready = dm_tready[117];
            assign ap_axis_iarg_117_tlast = ap_tlast[117];
            assign ap_axis_iarg_117_tvalid = ap_tvalid[117];
            assign ap_axis_iarg_117_tkeep = ap_tkeep[117][S_AXIS_IARG_117_WIDTH/8-1:0];
            assign ap_axis_iarg_117_tstrb = ap_tstrb[117][S_AXIS_IARG_117_WIDTH/8-1:0];
            assign ap_axis_iarg_117_tdata = ap_tdata[117][S_AXIS_IARG_117_WIDTH-1:0];
            assign ap_tready[117] = ap_axis_iarg_117_tready;
        end
        if(C_NUM_INPUT_AXISs > 118) begin
            assign axis_clk[118] = s_axis_iarg_118_aclk;
            assign axis_rst[118] = s_axis_iarg_118_aresetn;
            assign dm_tlast[118] = s_axis_iarg_118_tlast;
            assign dm_tvalid[118] = s_axis_iarg_118_tvalid;
            assign dm_tkeep[118][S_AXIS_IARG_118_DMWIDTH/8-1:0] = s_axis_iarg_118_tkeep;
            assign dm_tstrb[118][S_AXIS_IARG_118_DMWIDTH/8-1:0] = s_axis_iarg_118_tstrb;
            assign dm_tdata[118][S_AXIS_IARG_118_DMWIDTH-1:0] = s_axis_iarg_118_tdata;
            assign s_axis_iarg_118_tready = dm_tready[118];
            assign ap_axis_iarg_118_tlast = ap_tlast[118];
            assign ap_axis_iarg_118_tvalid = ap_tvalid[118];
            assign ap_axis_iarg_118_tkeep = ap_tkeep[118][S_AXIS_IARG_118_WIDTH/8-1:0];
            assign ap_axis_iarg_118_tstrb = ap_tstrb[118][S_AXIS_IARG_118_WIDTH/8-1:0];
            assign ap_axis_iarg_118_tdata = ap_tdata[118][S_AXIS_IARG_118_WIDTH-1:0];
            assign ap_tready[118] = ap_axis_iarg_118_tready;
        end
        if(C_NUM_INPUT_AXISs > 119) begin
            assign axis_clk[119] = s_axis_iarg_119_aclk;
            assign axis_rst[119] = s_axis_iarg_119_aresetn;
            assign dm_tlast[119] = s_axis_iarg_119_tlast;
            assign dm_tvalid[119] = s_axis_iarg_119_tvalid;
            assign dm_tkeep[119][S_AXIS_IARG_119_DMWIDTH/8-1:0] = s_axis_iarg_119_tkeep;
            assign dm_tstrb[119][S_AXIS_IARG_119_DMWIDTH/8-1:0] = s_axis_iarg_119_tstrb;
            assign dm_tdata[119][S_AXIS_IARG_119_DMWIDTH-1:0] = s_axis_iarg_119_tdata;
            assign s_axis_iarg_119_tready = dm_tready[119];
            assign ap_axis_iarg_119_tlast = ap_tlast[119];
            assign ap_axis_iarg_119_tvalid = ap_tvalid[119];
            assign ap_axis_iarg_119_tkeep = ap_tkeep[119][S_AXIS_IARG_119_WIDTH/8-1:0];
            assign ap_axis_iarg_119_tstrb = ap_tstrb[119][S_AXIS_IARG_119_WIDTH/8-1:0];
            assign ap_axis_iarg_119_tdata = ap_tdata[119][S_AXIS_IARG_119_WIDTH-1:0];
            assign ap_tready[119] = ap_axis_iarg_119_tready;
        end
        if(C_NUM_INPUT_AXISs > 120) begin
            assign axis_clk[120] = s_axis_iarg_120_aclk;
            assign axis_rst[120] = s_axis_iarg_120_aresetn;
            assign dm_tlast[120] = s_axis_iarg_120_tlast;
            assign dm_tvalid[120] = s_axis_iarg_120_tvalid;
            assign dm_tkeep[120][S_AXIS_IARG_120_DMWIDTH/8-1:0] = s_axis_iarg_120_tkeep;
            assign dm_tstrb[120][S_AXIS_IARG_120_DMWIDTH/8-1:0] = s_axis_iarg_120_tstrb;
            assign dm_tdata[120][S_AXIS_IARG_120_DMWIDTH-1:0] = s_axis_iarg_120_tdata;
            assign s_axis_iarg_120_tready = dm_tready[120];
            assign ap_axis_iarg_120_tlast = ap_tlast[120];
            assign ap_axis_iarg_120_tvalid = ap_tvalid[120];
            assign ap_axis_iarg_120_tkeep = ap_tkeep[120][S_AXIS_IARG_120_WIDTH/8-1:0];
            assign ap_axis_iarg_120_tstrb = ap_tstrb[120][S_AXIS_IARG_120_WIDTH/8-1:0];
            assign ap_axis_iarg_120_tdata = ap_tdata[120][S_AXIS_IARG_120_WIDTH-1:0];
            assign ap_tready[120] = ap_axis_iarg_120_tready;
        end
        if(C_NUM_INPUT_AXISs > 121) begin
            assign axis_clk[121] = s_axis_iarg_121_aclk;
            assign axis_rst[121] = s_axis_iarg_121_aresetn;
            assign dm_tlast[121] = s_axis_iarg_121_tlast;
            assign dm_tvalid[121] = s_axis_iarg_121_tvalid;
            assign dm_tkeep[121][S_AXIS_IARG_121_DMWIDTH/8-1:0] = s_axis_iarg_121_tkeep;
            assign dm_tstrb[121][S_AXIS_IARG_121_DMWIDTH/8-1:0] = s_axis_iarg_121_tstrb;
            assign dm_tdata[121][S_AXIS_IARG_121_DMWIDTH-1:0] = s_axis_iarg_121_tdata;
            assign s_axis_iarg_121_tready = dm_tready[121];
            assign ap_axis_iarg_121_tlast = ap_tlast[121];
            assign ap_axis_iarg_121_tvalid = ap_tvalid[121];
            assign ap_axis_iarg_121_tkeep = ap_tkeep[121][S_AXIS_IARG_121_WIDTH/8-1:0];
            assign ap_axis_iarg_121_tstrb = ap_tstrb[121][S_AXIS_IARG_121_WIDTH/8-1:0];
            assign ap_axis_iarg_121_tdata = ap_tdata[121][S_AXIS_IARG_121_WIDTH-1:0];
            assign ap_tready[121] = ap_axis_iarg_121_tready;
        end
        if(C_NUM_INPUT_AXISs > 122) begin
            assign axis_clk[122] = s_axis_iarg_122_aclk;
            assign axis_rst[122] = s_axis_iarg_122_aresetn;
            assign dm_tlast[122] = s_axis_iarg_122_tlast;
            assign dm_tvalid[122] = s_axis_iarg_122_tvalid;
            assign dm_tkeep[122][S_AXIS_IARG_122_DMWIDTH/8-1:0] = s_axis_iarg_122_tkeep;
            assign dm_tstrb[122][S_AXIS_IARG_122_DMWIDTH/8-1:0] = s_axis_iarg_122_tstrb;
            assign dm_tdata[122][S_AXIS_IARG_122_DMWIDTH-1:0] = s_axis_iarg_122_tdata;
            assign s_axis_iarg_122_tready = dm_tready[122];
            assign ap_axis_iarg_122_tlast = ap_tlast[122];
            assign ap_axis_iarg_122_tvalid = ap_tvalid[122];
            assign ap_axis_iarg_122_tkeep = ap_tkeep[122][S_AXIS_IARG_122_WIDTH/8-1:0];
            assign ap_axis_iarg_122_tstrb = ap_tstrb[122][S_AXIS_IARG_122_WIDTH/8-1:0];
            assign ap_axis_iarg_122_tdata = ap_tdata[122][S_AXIS_IARG_122_WIDTH-1:0];
            assign ap_tready[122] = ap_axis_iarg_122_tready;
        end
        if(C_NUM_INPUT_AXISs > 123) begin
            assign axis_clk[123] = s_axis_iarg_123_aclk;
            assign axis_rst[123] = s_axis_iarg_123_aresetn;
            assign dm_tlast[123] = s_axis_iarg_123_tlast;
            assign dm_tvalid[123] = s_axis_iarg_123_tvalid;
            assign dm_tkeep[123][S_AXIS_IARG_123_DMWIDTH/8-1:0] = s_axis_iarg_123_tkeep;
            assign dm_tstrb[123][S_AXIS_IARG_123_DMWIDTH/8-1:0] = s_axis_iarg_123_tstrb;
            assign dm_tdata[123][S_AXIS_IARG_123_DMWIDTH-1:0] = s_axis_iarg_123_tdata;
            assign s_axis_iarg_123_tready = dm_tready[123];
            assign ap_axis_iarg_123_tlast = ap_tlast[123];
            assign ap_axis_iarg_123_tvalid = ap_tvalid[123];
            assign ap_axis_iarg_123_tkeep = ap_tkeep[123][S_AXIS_IARG_123_WIDTH/8-1:0];
            assign ap_axis_iarg_123_tstrb = ap_tstrb[123][S_AXIS_IARG_123_WIDTH/8-1:0];
            assign ap_axis_iarg_123_tdata = ap_tdata[123][S_AXIS_IARG_123_WIDTH-1:0];
            assign ap_tready[123] = ap_axis_iarg_123_tready;
        end
        if(C_NUM_INPUT_AXISs > 124) begin
            assign axis_clk[124] = s_axis_iarg_124_aclk;
            assign axis_rst[124] = s_axis_iarg_124_aresetn;
            assign dm_tlast[124] = s_axis_iarg_124_tlast;
            assign dm_tvalid[124] = s_axis_iarg_124_tvalid;
            assign dm_tkeep[124][S_AXIS_IARG_124_DMWIDTH/8-1:0] = s_axis_iarg_124_tkeep;
            assign dm_tstrb[124][S_AXIS_IARG_124_DMWIDTH/8-1:0] = s_axis_iarg_124_tstrb;
            assign dm_tdata[124][S_AXIS_IARG_124_DMWIDTH-1:0] = s_axis_iarg_124_tdata;
            assign s_axis_iarg_124_tready = dm_tready[124];
            assign ap_axis_iarg_124_tlast = ap_tlast[124];
            assign ap_axis_iarg_124_tvalid = ap_tvalid[124];
            assign ap_axis_iarg_124_tkeep = ap_tkeep[124][S_AXIS_IARG_124_WIDTH/8-1:0];
            assign ap_axis_iarg_124_tstrb = ap_tstrb[124][S_AXIS_IARG_124_WIDTH/8-1:0];
            assign ap_axis_iarg_124_tdata = ap_tdata[124][S_AXIS_IARG_124_WIDTH-1:0];
            assign ap_tready[124] = ap_axis_iarg_124_tready;
        end
        if(C_NUM_INPUT_AXISs > 125) begin
            assign axis_clk[125] = s_axis_iarg_125_aclk;
            assign axis_rst[125] = s_axis_iarg_125_aresetn;
            assign dm_tlast[125] = s_axis_iarg_125_tlast;
            assign dm_tvalid[125] = s_axis_iarg_125_tvalid;
            assign dm_tkeep[125][S_AXIS_IARG_125_DMWIDTH/8-1:0] = s_axis_iarg_125_tkeep;
            assign dm_tstrb[125][S_AXIS_IARG_125_DMWIDTH/8-1:0] = s_axis_iarg_125_tstrb;
            assign dm_tdata[125][S_AXIS_IARG_125_DMWIDTH-1:0] = s_axis_iarg_125_tdata;
            assign s_axis_iarg_125_tready = dm_tready[125];
            assign ap_axis_iarg_125_tlast = ap_tlast[125];
            assign ap_axis_iarg_125_tvalid = ap_tvalid[125];
            assign ap_axis_iarg_125_tkeep = ap_tkeep[125][S_AXIS_IARG_125_WIDTH/8-1:0];
            assign ap_axis_iarg_125_tstrb = ap_tstrb[125][S_AXIS_IARG_125_WIDTH/8-1:0];
            assign ap_axis_iarg_125_tdata = ap_tdata[125][S_AXIS_IARG_125_WIDTH-1:0];
            assign ap_tready[125] = ap_axis_iarg_125_tready;
        end
        if(C_NUM_INPUT_AXISs > 126) begin
            assign axis_clk[126] = s_axis_iarg_126_aclk;
            assign axis_rst[126] = s_axis_iarg_126_aresetn;
            assign dm_tlast[126] = s_axis_iarg_126_tlast;
            assign dm_tvalid[126] = s_axis_iarg_126_tvalid;
            assign dm_tkeep[126][S_AXIS_IARG_126_DMWIDTH/8-1:0] = s_axis_iarg_126_tkeep;
            assign dm_tstrb[126][S_AXIS_IARG_126_DMWIDTH/8-1:0] = s_axis_iarg_126_tstrb;
            assign dm_tdata[126][S_AXIS_IARG_126_DMWIDTH-1:0] = s_axis_iarg_126_tdata;
            assign s_axis_iarg_126_tready = dm_tready[126];
            assign ap_axis_iarg_126_tlast = ap_tlast[126];
            assign ap_axis_iarg_126_tvalid = ap_tvalid[126];
            assign ap_axis_iarg_126_tkeep = ap_tkeep[126][S_AXIS_IARG_126_WIDTH/8-1:0];
            assign ap_axis_iarg_126_tstrb = ap_tstrb[126][S_AXIS_IARG_126_WIDTH/8-1:0];
            assign ap_axis_iarg_126_tdata = ap_tdata[126][S_AXIS_IARG_126_WIDTH-1:0];
            assign ap_tready[126] = ap_axis_iarg_126_tready;
        end
        if(C_NUM_INPUT_AXISs > 127) begin
            assign axis_clk[127] = s_axis_iarg_127_aclk;
            assign axis_rst[127] = s_axis_iarg_127_aresetn;
            assign dm_tlast[127] = s_axis_iarg_127_tlast;
            assign dm_tvalid[127] = s_axis_iarg_127_tvalid;
            assign dm_tkeep[127][S_AXIS_IARG_127_DMWIDTH/8-1:0] = s_axis_iarg_127_tkeep;
            assign dm_tstrb[127][S_AXIS_IARG_127_DMWIDTH/8-1:0] = s_axis_iarg_127_tstrb;
            assign dm_tdata[127][S_AXIS_IARG_127_DMWIDTH-1:0] = s_axis_iarg_127_tdata;
            assign s_axis_iarg_127_tready = dm_tready[127];
            assign ap_axis_iarg_127_tlast = ap_tlast[127];
            assign ap_axis_iarg_127_tvalid = ap_tvalid[127];
            assign ap_axis_iarg_127_tkeep = ap_tkeep[127][S_AXIS_IARG_127_WIDTH/8-1:0];
            assign ap_axis_iarg_127_tstrb = ap_tstrb[127][S_AXIS_IARG_127_WIDTH/8-1:0];
            assign ap_axis_iarg_127_tdata = ap_tdata[127][S_AXIS_IARG_127_WIDTH-1:0];
            assign ap_tready[127] = ap_axis_iarg_127_tready;
        end
    endgenerate
    
    //instantiate the axis2axis modules
    genvar idx;
    generate
        for(idx=0; idx<C_NUM_INPUT_AXISs; idx=idx+1) begin: IN_AXIS_GEN
            //check if data width converter is needed
            if(C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx] != C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]) begin
                 axis_dwidth_converter_v1_1_9_axis_dwidth_converter #(
                    .C_S_AXIS_TDATA_WIDTH(C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_M_AXIS_TDATA_WIDTH(C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_AXIS_TID_WIDTH(1),
                    .C_AXIS_TDEST_WIDTH(1),
                    .C_S_AXIS_TUSER_WIDTH(1),
                    .C_M_AXIS_TUSER_WIDTH(1),
                    .C_AXIS_SIGNAL_SET(32'h1F)  //Enabled: TLAST, TKEEP, TSTRB, TDATA, TREADY
                ) data_width_conv_i (
                    .aclk(axis_clk[idx]),
                    .aresetn(axis_rst[idx]),
                    .aclken(1'b1),
                    .s_axis_tvalid(dm_tvalid[idx]),
                    .s_axis_tready(dm_tready[idx]),
                    .s_axis_tdata(dm_tdata[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .s_axis_tstrb(dm_tstrb[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tkeep(dm_tkeep[idx][C_DMWIDTH_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0]),
                    .s_axis_tlast(dm_tlast[idx]),
//                    .s_axis_tid(),
//                    .s_axis_tdest(),
//                    .s_axis_tuser(),
                    .m_axis_tvalid(dwconv_tvalid[idx]),
                    .m_axis_tready(dwconv_tready[idx]),
                    .m_axis_tdata(dwconv_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
//                    .m_axis_tstrb(),
//                    .m_axis_tkeep(),
                    .m_axis_tlast(dwconv_tlast[idx])
//                    .m_axis_tid(),
//                    .m_axis_tdest(),
//                    .m_axis_tuser()
                );
            end
            else begin
                //if no buffering, wire the input signals straight through
                assign dwconv_tlast[idx] = dm_tlast[idx];
                assign dwconv_tvalid[idx] = dm_tvalid[idx];
                assign dm_tready[idx] = dwconv_tready[idx];   //output
                assign dwconv_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = dm_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            end
            
            if(C_DEPTH_BIT_ARRAY[32*(idx+1)-1:32*idx] > 0) begin
                //use fifo
                axis_fifo #(
                    .C_DATA_WIDTH(C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_DATA_DEPTH(C_DEPTH_BIT_ARRAY[32*(idx+1)-1:32*idx]),
                    .C_IS_ASYNC(C_IS_ASYNC_BIT_ARRAY[32*(idx+1)-1:32*idx])
                ) axis_fifo_i (
                    .aresetn(axis_rst[idx]),
                    .inclk(axis_clk[idx]),
                    .in_tdata(dwconv_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .in_tlast(dwconv_tlast[idx]),  
                    .in_tvalid(dwconv_tvalid[idx]),
                    .in_tready(dwconv_tready[idx]),
                    .outclk(acc_clk), 
                    .out_tdata(buf_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                    .out_tready(buf_tready[idx]),
                    .out_tvalid(buf_tvalid[idx]),
                    .out_tlast(buf_tlast[idx])
                );
            end
            else begin
                //if not, wire the input signals straight through
                assign buf_tlast[idx] = dwconv_tlast[idx];
                assign buf_tvalid[idx] = dwconv_tvalid[idx];
                assign dwconv_tready[idx] = buf_tready[idx];   //output
                assign buf_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = dwconv_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            end
            
            inaxis #( 
                .DATA_WIDTH(C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx])
            ) inaxis_i (
                .ACC_CLK(acc_clk),
                .ARESETN(acc_aresetn),
                .CTRL_ALLOW(in_axis_allow),
                .CTRL_READY(in_axis_ready[idx]),
                .CTRL_FINISHED(in_axis_finished[idx]),
                .DM_TLAST(buf_tlast[idx]),
                .DM_TVALID(buf_tvalid[idx]),
                .DM_TDATA(buf_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .DM_TREADY(buf_tready[idx]),
                .AP_TLAST(ap_tlast[idx]),
                .AP_TVALID(ap_tvalid[idx]),
                .AP_TDATA(ap_tdata[idx][C_INAXIS_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0]),
                .AP_TREADY(ap_tready[idx])
            );
        end
    endgenerate
endmodule
