// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689
`timescale 1ns / 1ps

module top #(
    //adapter parameters
    parameter C_HAS_CTRL = 1,
    parameter C_ACC_RESET_POLARITY = 0,
    parameter C_QUEUE_DEPTH = 16,
    
    //scalar parameters
    parameter C_N_INPUT_SCALARS = 0,
    parameter C_N_OUTPUT_SCALARS = 0,
    parameter C_FIFO_DEPTH = 16,
    parameter C_HAS_RETURN = 0,
    parameter [31:0] C_INPUT_SCALAR_0_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_1_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_2_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_3_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_4_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_5_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_6_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_7_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_8_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_9_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_10_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_11_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_12_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_13_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_14_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_15_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_16_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_17_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_18_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_19_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_20_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_21_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_22_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_23_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_24_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_25_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_26_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_27_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_28_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_29_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_30_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_31_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_32_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_33_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_34_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_35_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_36_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_37_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_38_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_39_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_40_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_41_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_42_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_43_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_44_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_45_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_46_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_47_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_48_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_49_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_50_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_51_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_52_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_53_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_54_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_55_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_56_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_57_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_58_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_59_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_60_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_61_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_62_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_63_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_64_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_65_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_66_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_67_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_68_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_69_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_70_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_71_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_72_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_73_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_74_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_75_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_76_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_77_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_78_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_79_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_80_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_81_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_82_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_83_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_84_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_85_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_86_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_87_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_88_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_89_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_90_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_91_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_92_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_93_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_94_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_95_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_96_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_97_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_98_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_99_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_100_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_101_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_102_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_103_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_104_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_105_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_106_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_107_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_108_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_109_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_110_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_111_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_112_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_113_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_114_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_115_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_116_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_117_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_118_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_119_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_120_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_121_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_122_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_123_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_124_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_125_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_126_WIDTH = 1,
    parameter [31:0] C_INPUT_SCALAR_127_WIDTH = 1,
    parameter [31:0] S_AXIS_SCALAR_0_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_1_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_2_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_3_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_4_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_5_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_6_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_7_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_8_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_9_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_10_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_11_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_12_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_13_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_14_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_15_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_16_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_17_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_18_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_19_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_20_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_21_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_22_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_23_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_24_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_25_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_26_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_27_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_28_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_29_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_30_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_31_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_32_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_33_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_34_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_35_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_36_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_37_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_38_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_39_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_40_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_41_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_42_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_43_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_44_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_45_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_46_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_47_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_48_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_49_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_50_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_51_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_52_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_53_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_54_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_55_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_56_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_57_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_58_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_59_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_60_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_61_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_62_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_63_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_64_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_65_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_66_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_67_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_68_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_69_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_70_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_71_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_72_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_73_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_74_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_75_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_76_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_77_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_78_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_79_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_80_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_81_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_82_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_83_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_84_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_85_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_86_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_87_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_88_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_89_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_90_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_91_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_92_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_93_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_94_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_95_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_96_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_97_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_98_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_99_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_100_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_101_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_102_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_103_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_104_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_105_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_106_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_107_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_108_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_109_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_110_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_111_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_112_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_113_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_114_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_115_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_116_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_117_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_118_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_119_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_120_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_121_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_122_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_123_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_124_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_125_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_126_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_127_IS_DIRECT = 0,
    parameter [31:0] S_AXIS_SCALAR_0_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_1_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_2_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_3_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_4_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_5_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_6_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_7_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_8_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_9_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_10_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_11_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_12_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_13_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_14_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_15_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_16_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_17_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_18_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_19_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_20_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_21_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_22_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_23_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_24_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_25_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_26_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_27_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_28_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_29_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_30_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_31_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_32_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_33_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_34_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_35_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_36_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_37_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_38_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_39_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_40_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_41_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_42_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_43_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_44_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_45_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_46_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_47_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_48_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_49_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_50_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_51_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_52_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_53_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_54_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_55_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_56_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_57_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_58_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_59_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_60_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_61_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_62_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_63_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_64_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_65_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_66_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_67_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_68_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_69_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_70_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_71_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_72_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_73_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_74_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_75_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_76_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_77_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_78_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_79_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_80_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_81_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_82_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_83_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_84_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_85_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_86_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_87_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_88_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_89_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_90_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_91_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_92_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_93_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_94_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_95_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_96_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_97_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_98_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_99_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_100_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_101_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_102_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_103_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_104_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_105_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_106_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_107_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_108_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_109_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_110_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_111_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_112_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_113_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_114_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_115_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_116_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_117_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_118_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_119_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_120_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_121_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_122_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_123_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_124_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_125_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_126_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_127_DIRECT_DMWIDTH = 32,
    parameter [31:0] S_AXIS_SCALAR_0_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_1_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_2_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_3_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_4_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_5_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_6_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_7_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_8_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_9_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_10_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_11_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_12_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_13_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_14_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_15_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_16_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_17_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_18_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_19_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_20_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_21_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_22_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_23_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_24_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_25_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_26_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_27_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_28_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_29_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_30_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_31_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_32_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_33_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_34_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_35_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_36_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_37_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_38_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_39_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_40_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_41_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_42_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_43_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_44_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_45_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_46_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_47_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_48_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_49_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_50_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_51_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_52_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_53_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_54_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_55_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_56_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_57_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_58_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_59_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_60_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_61_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_62_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_63_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_64_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_65_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_66_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_67_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_68_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_69_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_70_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_71_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_72_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_73_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_74_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_75_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_76_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_77_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_78_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_79_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_80_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_81_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_82_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_83_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_84_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_85_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_86_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_87_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_88_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_89_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_90_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_91_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_92_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_93_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_94_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_95_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_96_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_97_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_98_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_99_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_100_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_101_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_102_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_103_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_104_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_105_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_106_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_107_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_108_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_109_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_110_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_111_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_112_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_113_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_114_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_115_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_116_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_117_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_118_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_119_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_120_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_121_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_122_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_123_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_124_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_125_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_126_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_127_DIRECT_IS_ASYNC = 1,
    parameter [31:0] S_AXIS_SCALAR_0_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_1_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_2_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_3_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_4_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_5_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_6_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_7_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_8_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_9_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_10_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_11_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_12_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_13_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_14_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_15_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_16_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_17_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_18_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_19_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_20_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_21_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_22_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_23_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_24_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_25_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_26_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_27_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_28_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_29_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_30_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_31_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_32_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_33_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_34_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_35_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_36_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_37_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_38_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_39_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_40_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_41_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_42_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_43_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_44_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_45_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_46_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_47_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_48_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_49_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_50_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_51_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_52_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_53_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_54_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_55_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_56_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_57_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_58_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_59_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_60_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_61_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_62_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_63_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_64_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_65_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_66_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_67_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_68_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_69_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_70_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_71_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_72_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_73_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_74_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_75_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_76_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_77_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_78_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_79_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_80_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_81_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_82_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_83_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_84_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_85_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_86_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_87_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_88_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_89_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_90_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_91_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_92_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_93_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_94_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_95_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_96_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_97_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_98_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_99_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_100_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_101_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_102_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_103_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_104_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_105_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_106_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_107_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_108_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_109_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_110_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_111_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_112_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_113_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_114_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_115_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_116_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_117_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_118_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_119_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_120_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_121_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_122_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_123_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_124_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_125_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_126_DIRECT_DEPTH = 16,
    parameter [31:0] S_AXIS_SCALAR_127_DIRECT_DEPTH = 16,
    parameter [31:0]  C_OUTPUT_SCALAR_0_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_1_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_2_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_3_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_4_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_5_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_6_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_7_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_8_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_9_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_10_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_11_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_12_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_13_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_14_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_15_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_16_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_17_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_18_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_19_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_20_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_21_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_22_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_23_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_24_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_25_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_26_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_27_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_28_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_29_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_30_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_31_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_32_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_33_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_34_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_35_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_36_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_37_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_38_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_39_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_40_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_41_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_42_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_43_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_44_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_45_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_46_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_47_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_48_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_49_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_50_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_51_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_52_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_53_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_54_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_55_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_56_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_57_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_58_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_59_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_60_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_61_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_62_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_63_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_64_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_65_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_66_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_67_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_68_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_69_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_70_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_71_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_72_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_73_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_74_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_75_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_76_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_77_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_78_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_79_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_80_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_81_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_82_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_83_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_84_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_85_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_86_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_87_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_88_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_89_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_90_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_91_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_92_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_93_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_94_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_95_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_96_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_97_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_98_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_99_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_100_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_101_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_102_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_103_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_104_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_105_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_106_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_107_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_108_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_109_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_110_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_111_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_112_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_113_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_114_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_115_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_116_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_117_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_118_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_119_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_120_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_121_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_122_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_123_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_124_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_125_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_126_WIDTH = 1,
    parameter [31:0]  C_OUTPUT_SCALAR_127_WIDTH = 1,
    parameter [31:0]  M_AXIS_SCALAR_0_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_1_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_2_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_3_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_4_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_5_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_6_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_7_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_8_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_9_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_10_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_11_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_12_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_13_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_14_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_15_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_16_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_17_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_18_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_19_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_20_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_21_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_22_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_23_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_24_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_25_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_26_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_27_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_28_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_29_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_30_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_31_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_32_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_33_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_34_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_35_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_36_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_37_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_38_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_39_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_40_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_41_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_42_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_43_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_44_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_45_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_46_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_47_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_48_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_49_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_50_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_51_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_52_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_53_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_54_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_55_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_56_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_57_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_58_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_59_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_60_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_61_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_62_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_63_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_64_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_65_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_66_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_67_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_68_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_69_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_70_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_71_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_72_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_73_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_74_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_75_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_76_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_77_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_78_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_79_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_80_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_81_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_82_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_83_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_84_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_85_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_86_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_87_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_88_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_89_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_90_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_91_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_92_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_93_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_94_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_95_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_96_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_97_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_98_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_99_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_100_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_101_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_102_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_103_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_104_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_105_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_106_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_107_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_108_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_109_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_110_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_111_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_112_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_113_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_114_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_115_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_116_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_117_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_118_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_119_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_120_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_121_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_122_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_123_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_124_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_125_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_126_IS_DIRECT = 0,
    parameter [31:0]  M_AXIS_SCALAR_127_IS_DIRECT = 0,
    parameter [31:0] M_AXIS_SCALAR_0_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_1_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_2_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_3_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_4_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_5_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_6_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_7_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_8_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_9_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_10_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_11_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_12_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_13_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_14_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_15_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_16_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_17_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_18_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_19_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_20_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_21_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_22_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_23_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_24_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_25_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_26_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_27_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_28_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_29_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_30_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_31_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_32_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_33_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_34_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_35_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_36_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_37_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_38_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_39_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_40_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_41_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_42_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_43_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_44_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_45_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_46_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_47_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_48_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_49_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_50_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_51_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_52_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_53_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_54_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_55_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_56_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_57_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_58_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_59_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_60_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_61_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_62_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_63_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_64_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_65_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_66_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_67_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_68_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_69_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_70_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_71_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_72_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_73_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_74_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_75_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_76_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_77_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_78_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_79_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_80_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_81_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_82_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_83_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_84_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_85_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_86_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_87_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_88_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_89_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_90_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_91_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_92_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_93_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_94_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_95_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_96_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_97_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_98_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_99_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_100_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_101_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_102_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_103_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_104_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_105_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_106_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_107_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_108_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_109_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_110_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_111_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_112_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_113_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_114_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_115_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_116_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_117_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_118_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_119_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_120_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_121_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_122_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_123_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_124_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_125_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_126_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_127_DIRECT_DMWIDTH = 32,
    parameter [31:0] M_AXIS_SCALAR_0_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_1_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_2_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_3_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_4_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_5_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_6_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_7_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_8_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_9_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_10_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_11_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_12_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_13_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_14_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_15_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_16_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_17_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_18_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_19_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_20_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_21_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_22_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_23_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_24_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_25_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_26_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_27_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_28_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_29_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_30_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_31_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_32_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_33_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_34_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_35_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_36_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_37_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_38_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_39_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_40_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_41_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_42_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_43_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_44_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_45_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_46_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_47_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_48_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_49_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_50_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_51_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_52_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_53_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_54_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_55_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_56_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_57_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_58_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_59_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_60_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_61_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_62_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_63_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_64_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_65_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_66_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_67_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_68_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_69_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_70_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_71_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_72_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_73_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_74_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_75_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_76_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_77_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_78_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_79_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_80_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_81_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_82_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_83_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_84_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_85_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_86_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_87_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_88_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_89_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_90_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_91_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_92_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_93_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_94_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_95_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_96_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_97_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_98_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_99_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_100_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_101_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_102_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_103_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_104_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_105_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_106_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_107_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_108_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_109_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_110_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_111_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_112_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_113_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_114_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_115_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_116_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_117_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_118_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_119_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_120_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_121_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_122_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_123_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_124_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_125_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_126_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_127_DIRECT_IS_ASYNC = 1,
    parameter [31:0] M_AXIS_SCALAR_0_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_1_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_2_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_3_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_4_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_5_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_6_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_7_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_8_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_9_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_10_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_11_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_12_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_13_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_14_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_15_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_16_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_17_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_18_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_19_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_20_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_21_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_22_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_23_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_24_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_25_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_26_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_27_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_28_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_29_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_30_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_31_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_32_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_33_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_34_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_35_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_36_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_37_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_38_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_39_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_40_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_41_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_42_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_43_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_44_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_45_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_46_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_47_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_48_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_49_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_50_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_51_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_52_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_53_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_54_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_55_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_56_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_57_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_58_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_59_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_60_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_61_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_62_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_63_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_64_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_65_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_66_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_67_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_68_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_69_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_70_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_71_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_72_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_73_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_74_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_75_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_76_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_77_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_78_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_79_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_80_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_81_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_82_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_83_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_84_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_85_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_86_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_87_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_88_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_89_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_90_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_91_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_92_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_93_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_94_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_95_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_96_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_97_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_98_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_99_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_100_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_101_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_102_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_103_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_104_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_105_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_106_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_107_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_108_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_109_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_110_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_111_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_112_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_113_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_114_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_115_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_116_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_117_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_118_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_119_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_120_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_121_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_122_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_123_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_124_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_125_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_126_DIRECT_DEPTH = 16,
    parameter [31:0] M_AXIS_SCALAR_127_DIRECT_DEPTH = 16,
    
    //fifo arg parameters
    parameter C_NUM_INPUT_FIFOs = 0,                //number of input fifo interfaces on the accelerator
    parameter C_NUM_OUTPUT_FIFOs = 0,               //number of output fifo interfaces on the accelerator
    parameter [31:0] S_AXIS_FIFO_0_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_1_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_2_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_3_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_4_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_5_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_6_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_7_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_8_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_9_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_10_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_11_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_12_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_13_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_14_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_15_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_16_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_17_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_18_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_19_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_20_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_21_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_22_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_23_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_24_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_25_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_26_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_27_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_28_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_29_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_30_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_31_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_32_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_33_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_34_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_35_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_36_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_37_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_38_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_39_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_40_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_41_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_42_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_43_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_44_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_45_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_46_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_47_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_48_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_49_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_50_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_51_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_52_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_53_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_54_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_55_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_56_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_57_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_58_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_59_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_60_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_61_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_62_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_63_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_64_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_65_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_66_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_67_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_68_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_69_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_70_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_71_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_72_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_73_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_74_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_75_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_76_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_77_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_78_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_79_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_80_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_81_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_82_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_83_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_84_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_85_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_86_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_87_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_88_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_89_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_90_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_91_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_92_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_93_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_94_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_95_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_96_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_97_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_98_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_99_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_100_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_101_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_102_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_103_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_104_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_105_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_106_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_107_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_108_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_109_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_110_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_111_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_112_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_113_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_114_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_115_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_116_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_117_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_118_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_119_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_120_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_121_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_122_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_123_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_124_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_125_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_126_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_127_WIDTH = 8,     //width of input fifo interface on the accelerator
    parameter [31:0] S_AXIS_FIFO_0_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_1_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_2_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_3_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_4_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_5_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_6_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_7_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_8_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_9_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_10_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_11_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_12_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_13_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_14_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_15_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_16_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_17_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_18_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_19_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_20_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_21_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_22_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_23_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_24_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_25_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_26_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_27_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_28_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_29_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_30_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_31_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_32_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_33_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_34_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_35_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_36_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_37_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_38_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_39_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_40_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_41_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_42_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_43_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_44_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_45_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_46_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_47_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_48_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_49_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_50_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_51_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_52_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_53_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_54_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_55_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_56_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_57_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_58_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_59_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_60_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_61_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_62_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_63_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_64_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_65_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_66_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_67_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_68_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_69_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_70_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_71_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_72_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_73_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_74_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_75_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_76_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_77_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_78_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_79_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_80_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_81_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_82_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_83_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_84_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_85_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_86_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_87_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_88_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_89_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_90_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_91_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_92_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_93_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_94_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_95_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_96_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_97_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_98_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_99_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_100_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_101_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_102_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_103_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_104_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_105_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_106_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_107_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_108_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_109_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_110_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_111_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_112_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_113_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_114_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_115_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_116_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_117_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_118_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_119_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_120_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_121_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_122_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_123_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_124_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_125_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_126_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_127_DEPTH = 16,      //depth of FIFO in adapter for input fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_FIFO_0_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_1_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_2_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_3_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_4_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_5_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_6_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_7_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_8_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_9_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_10_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_11_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_12_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_13_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_14_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_15_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_16_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_17_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_18_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_19_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_20_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_21_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_22_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_23_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_24_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_25_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_26_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_27_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_28_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_29_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_30_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_31_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_32_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_33_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_34_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_35_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_36_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_37_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_38_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_39_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_40_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_41_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_42_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_43_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_44_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_45_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_46_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_47_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_48_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_49_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_50_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_51_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_52_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_53_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_54_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_55_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_56_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_57_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_58_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_59_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_60_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_61_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_62_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_63_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_64_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_65_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_66_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_67_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_68_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_69_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_70_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_71_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_72_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_73_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_74_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_75_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_76_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_77_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_78_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_79_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_80_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_81_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_82_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_83_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_84_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_85_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_86_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_87_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_88_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_89_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_90_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_91_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_92_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_93_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_94_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_95_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_96_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_97_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_98_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_99_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_100_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_101_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_102_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_103_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_104_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_105_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_106_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_107_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_108_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_109_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_110_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_111_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_112_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_113_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_114_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_115_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_116_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_117_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_118_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_119_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_120_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_121_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_122_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_123_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_124_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_125_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_126_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_127_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input fifo interface
    parameter [31:0] S_AXIS_FIFO_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_FIFO_0_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_1_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_2_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_3_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_4_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_5_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_6_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_7_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_8_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_9_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_10_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_11_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_12_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_13_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_14_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_15_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_16_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_17_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_18_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_19_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_20_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_21_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_22_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_23_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_24_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_25_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_26_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_27_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_28_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_29_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_30_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_31_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_32_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_33_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_34_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_35_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_36_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_37_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_38_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_39_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_40_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_41_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_42_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_43_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_44_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_45_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_46_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_47_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_48_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_49_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_50_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_51_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_52_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_53_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_54_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_55_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_56_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_57_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_58_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_59_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_60_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_61_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_62_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_63_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_64_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_65_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_66_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_67_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_68_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_69_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_70_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_71_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_72_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_73_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_74_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_75_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_76_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_77_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_78_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_79_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_80_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_81_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_82_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_83_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_84_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_85_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_86_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_87_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_88_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_89_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_90_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_91_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_92_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_93_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_94_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_95_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_96_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_97_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_98_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_99_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_100_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_101_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_102_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_103_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_104_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_105_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_106_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_107_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_108_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_109_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_110_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_111_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_112_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_113_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_114_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_115_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_116_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_117_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_118_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_119_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_120_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_121_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_122_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_123_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_124_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_125_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_126_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] S_AXIS_FIFO_127_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_0_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_1_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_2_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_3_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_4_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_5_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_6_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_7_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_8_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_9_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_10_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_11_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_12_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_13_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_14_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_15_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_16_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_17_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_18_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_19_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_20_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_21_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_22_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_23_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_24_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_25_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_26_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_27_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_28_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_29_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_30_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_31_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_32_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_33_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_34_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_35_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_36_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_37_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_38_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_39_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_40_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_41_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_42_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_43_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_44_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_45_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_46_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_47_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_48_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_49_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_50_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_51_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_52_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_53_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_54_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_55_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_56_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_57_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_58_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_59_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_60_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_61_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_62_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_63_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_64_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_65_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_66_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_67_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_68_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_69_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_70_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_71_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_72_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_73_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_74_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_75_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_76_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_77_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_78_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_79_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_80_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_81_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_82_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_83_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_84_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_85_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_86_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_87_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_88_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_89_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_90_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_91_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_92_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_93_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_94_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_95_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_96_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_97_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_98_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_99_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_100_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_101_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_102_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_103_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_104_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_105_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_106_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_107_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_108_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_109_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_110_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_111_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_112_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_113_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_114_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_115_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_116_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_117_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_118_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_119_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_120_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_121_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_122_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_123_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_124_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_125_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_126_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_127_WIDTH = 8,    //width of output fifo interface on the accelerator
    parameter [31:0] M_AXIS_FIFO_0_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_1_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_2_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_3_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_4_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_5_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_6_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_7_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_8_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_9_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_10_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_11_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_12_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_13_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_14_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_15_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_16_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_17_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_18_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_19_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_20_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_21_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_22_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_23_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_24_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_25_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_26_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_27_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_28_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_29_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_30_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_31_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_32_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_33_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_34_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_35_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_36_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_37_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_38_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_39_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_40_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_41_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_42_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_43_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_44_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_45_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_46_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_47_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_48_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_49_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_50_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_51_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_52_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_53_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_54_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_55_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_56_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_57_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_58_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_59_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_60_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_61_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_62_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_63_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_64_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_65_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_66_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_67_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_68_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_69_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_70_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_71_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_72_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_73_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_74_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_75_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_76_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_77_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_78_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_79_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_80_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_81_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_82_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_83_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_84_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_85_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_86_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_87_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_88_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_89_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_90_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_91_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_92_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_93_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_94_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_95_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_96_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_97_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_98_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_99_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_100_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_101_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_102_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_103_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_104_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_105_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_106_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_107_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_108_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_109_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_110_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_111_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_112_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_113_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_114_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_115_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_116_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_117_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_118_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_119_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_120_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_121_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_122_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_123_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_124_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_125_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_126_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_127_DEPTH = 16,     //depth of FIFO in adapter for output fifo interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_FIFO_0_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_1_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_2_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_3_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_4_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_5_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_6_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_7_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_8_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_9_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_10_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_11_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_12_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_13_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_14_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_15_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_16_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_17_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_18_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_19_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_20_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_21_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_22_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_23_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_24_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_25_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_26_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_27_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_28_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_29_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_30_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_31_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_32_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_33_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_34_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_35_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_36_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_37_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_38_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_39_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_40_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_41_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_42_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_43_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_44_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_45_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_46_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_47_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_48_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_49_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_50_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_51_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_52_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_53_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_54_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_55_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_56_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_57_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_58_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_59_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_60_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_61_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_62_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_63_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_64_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_65_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_66_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_67_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_68_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_69_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_70_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_71_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_72_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_73_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_74_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_75_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_76_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_77_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_78_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_79_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_80_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_81_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_82_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_83_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_84_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_85_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_86_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_87_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_88_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_89_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_90_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_91_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_92_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_93_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_94_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_95_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_96_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_97_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_98_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_99_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_100_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_101_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_102_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_103_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_104_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_105_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_106_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_107_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_108_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_109_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_110_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_111_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_112_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_113_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_114_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_115_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_116_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_117_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_118_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_119_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_120_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_121_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_122_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_123_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_124_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_125_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_126_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_127_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output fifo interface
    parameter [31:0] M_AXIS_FIFO_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_FIFO_0_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_1_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_2_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_3_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_4_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_5_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_6_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_7_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_8_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_9_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_10_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_11_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_12_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_13_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_14_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_15_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_16_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_17_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_18_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_19_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_20_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_21_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_22_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_23_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_24_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_25_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_26_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_27_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_28_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_29_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_30_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_31_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_32_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_33_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_34_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_35_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_36_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_37_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_38_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_39_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_40_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_41_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_42_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_43_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_44_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_45_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_46_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_47_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_48_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_49_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_50_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_51_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_52_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_53_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_54_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_55_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_56_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_57_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_58_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_59_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_60_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_61_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_62_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_63_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_64_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_65_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_66_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_67_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_68_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_69_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_70_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_71_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_72_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_73_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_74_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_75_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_76_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_77_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_78_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_79_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_80_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_81_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_82_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_83_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_84_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_85_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_86_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_87_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_88_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_89_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_90_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_91_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_92_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_93_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_94_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_95_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_96_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_97_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_98_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_99_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_100_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_101_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_102_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_103_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_104_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_105_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_106_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_107_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_108_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_109_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_110_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_111_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_112_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_113_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_114_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_115_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_116_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_117_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_118_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_119_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_120_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_121_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_122_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_123_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_124_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_125_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_126_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    parameter [31:0] M_AXIS_FIFO_127_BYTE_WIDTH = 8,     //width of input fifo interface on the accelerator, padded
    
    //bram arg parameters
    parameter C_NUM_INPUT_BRAMs = 0, 
    parameter C_NUM_OUTPUT_BRAMs = 0, 
    parameter S_AXIS_BRAM_0_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_1_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_2_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_3_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_4_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_5_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_6_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_7_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_8_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_9_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_10_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_11_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_12_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_13_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_14_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_15_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_16_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_17_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_18_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_19_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_20_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_21_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_22_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_23_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_24_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_25_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_26_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_27_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_28_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_29_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_30_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_31_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_32_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_33_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_34_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_35_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_36_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_37_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_38_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_39_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_40_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_41_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_42_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_43_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_44_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_45_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_46_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_47_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_48_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_49_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_50_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_51_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_52_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_53_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_54_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_55_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_56_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_57_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_58_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_59_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_60_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_61_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_62_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_63_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_64_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_65_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_66_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_67_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_68_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_69_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_70_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_71_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_72_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_73_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_74_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_75_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_76_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_77_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_78_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_79_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_80_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_81_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_82_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_83_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_84_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_85_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_86_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_87_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_88_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_89_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_90_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_91_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_92_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_93_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_94_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_95_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_96_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_97_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_98_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_99_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_100_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_101_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_102_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_103_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_104_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_105_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_106_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_107_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_108_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_109_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_110_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_111_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_112_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_113_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_114_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_115_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_116_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_117_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_118_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_119_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_120_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_121_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_122_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_123_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_124_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_125_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_126_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter S_AXIS_BRAM_127_PORTS = 1,            //number of bram ports (dual-ported, partitioned)
    parameter [31:0] S_AXIS_BRAM_0_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_1_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_2_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_3_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_4_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_5_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_6_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_7_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_8_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_9_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_10_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_11_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_12_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_13_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_14_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_15_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_16_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_17_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_18_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_19_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_20_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_21_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_22_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_23_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_24_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_25_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_26_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_27_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_28_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_29_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_30_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_31_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_32_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_33_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_34_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_35_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_36_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_37_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_38_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_39_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_40_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_41_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_42_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_43_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_44_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_45_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_46_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_47_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_48_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_49_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_50_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_51_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_52_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_53_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_54_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_55_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_56_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_57_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_58_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_59_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_60_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_61_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_62_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_63_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_64_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_65_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_66_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_67_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_68_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_69_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_70_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_71_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_72_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_73_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_74_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_75_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_76_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_77_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_78_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_79_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_80_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_81_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_82_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_83_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_84_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_85_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_86_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_87_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_88_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_89_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_90_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_91_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_92_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_93_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_94_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_95_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_96_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_97_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_98_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_99_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_100_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_101_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_102_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_103_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_104_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_105_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_106_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_107_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_108_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_109_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_110_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_111_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_112_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_113_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_114_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_115_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_116_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_117_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_118_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_119_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_120_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_121_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_122_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_123_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_124_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_125_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_126_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_127_WIDTH = 8,     //width of input bram interface on the accelerator
    parameter [31:0] S_AXIS_BRAM_0_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_1_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_2_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_3_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_4_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_5_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_6_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_7_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_8_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_9_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_10_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_11_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_12_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_13_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_14_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_15_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_16_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_17_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_18_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_19_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_20_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_21_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_22_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_23_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_24_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_25_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_26_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_27_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_28_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_29_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_30_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_31_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_32_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_33_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_34_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_35_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_36_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_37_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_38_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_39_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_40_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_41_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_42_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_43_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_44_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_45_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_46_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_47_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_48_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_49_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_50_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_51_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_52_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_53_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_54_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_55_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_56_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_57_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_58_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_59_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_60_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_61_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_62_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_63_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_64_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_65_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_66_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_67_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_68_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_69_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_70_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_71_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_72_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_73_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_74_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_75_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_76_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_77_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_78_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_79_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_80_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_81_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_82_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_83_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_84_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_85_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_86_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_87_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_88_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_89_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_90_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_91_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_92_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_93_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_94_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_95_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_96_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_97_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_98_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_99_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_100_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_101_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_102_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_103_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_104_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_105_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_106_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_107_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_108_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_109_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_110_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_111_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_112_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_113_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_114_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_115_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_116_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_117_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_118_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_119_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_120_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_121_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_122_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_123_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_124_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_125_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_126_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_127_DEPTH = 2,     //depth of BRAM in adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_0_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_1_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_2_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_3_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_4_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_5_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_6_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_7_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_8_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_9_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_10_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_11_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_12_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_13_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_14_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_15_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_16_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_17_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_18_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_19_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_20_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_21_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_22_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_23_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_24_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_25_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_26_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_27_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_28_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_29_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_30_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_31_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_32_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_33_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_34_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_35_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_36_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_37_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_38_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_39_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_40_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_41_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_42_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_43_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_44_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_45_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_46_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_47_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_48_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_49_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_50_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_51_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_52_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_53_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_54_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_55_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_56_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_57_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_58_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_59_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_60_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_61_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_62_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_63_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_64_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_65_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_66_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_67_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_68_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_69_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_70_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_71_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_72_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_73_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_74_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_75_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_76_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_77_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_78_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_79_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_80_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_81_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_82_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_83_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_84_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_85_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_86_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_87_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_88_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_89_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_90_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_91_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_92_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_93_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_94_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_95_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_96_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_97_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_98_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_99_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_100_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_101_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_102_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_103_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_104_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_105_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_106_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_107_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_108_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_109_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_110_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_111_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_112_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_113_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_114_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_115_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_116_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_117_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_118_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_119_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_120_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_121_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_122_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_123_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_124_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_125_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_126_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] S_AXIS_BRAM_127_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input bram interface
    parameter [31:0] M_AXIS_BRAMIO_0_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_1_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_2_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_3_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_4_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_5_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_6_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_7_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_8_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_9_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_10_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_11_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_12_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_13_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_14_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_15_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_16_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_17_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_18_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_19_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_20_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_21_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_22_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_23_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_24_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_25_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_26_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_27_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_28_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_29_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_30_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_31_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_32_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_33_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_34_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_35_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_36_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_37_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_38_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_39_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_40_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_41_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_42_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_43_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_44_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_45_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_46_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_47_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_48_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_49_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_50_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_51_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_52_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_53_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_54_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_55_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_56_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_57_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_58_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_59_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_60_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_61_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_62_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_63_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_64_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_65_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_66_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_67_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_68_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_69_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_70_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_71_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_72_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_73_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_74_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_75_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_76_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_77_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_78_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_79_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_80_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_81_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_82_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_83_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_84_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_85_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_86_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_87_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_88_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_89_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_90_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_91_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_92_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_93_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_94_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_95_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_96_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_97_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_98_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_99_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_100_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_101_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_102_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_103_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_104_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_105_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_106_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_107_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_108_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_109_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_110_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_111_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_112_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_113_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_114_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_115_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_116_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_117_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_118_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_119_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_120_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_121_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_122_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_123_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_124_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_125_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_126_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] M_AXIS_BRAMIO_127_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for inout (output) bram interface
    parameter [31:0] S_AXIS_BRAM_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_BRAM_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAMIO_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [0:0] S_AXIS_BRAM_0_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_1_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_2_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_3_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_4_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_5_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_6_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_7_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_8_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_9_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_10_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_11_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_12_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_13_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_14_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_15_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_16_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_17_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_18_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_19_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_20_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_21_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_22_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_23_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_24_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_25_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_26_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_27_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_28_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_29_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_30_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_31_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_32_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_33_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_34_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_35_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_36_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_37_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_38_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_39_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_40_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_41_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_42_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_43_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_44_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_45_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_46_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_47_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_48_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_49_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_50_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_51_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_52_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_53_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_54_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_55_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_56_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_57_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_58_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_59_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_60_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_61_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_62_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_63_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_64_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_65_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_66_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_67_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_68_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_69_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_70_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_71_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_72_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_73_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_74_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_75_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_76_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_77_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_78_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_79_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_80_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_81_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_82_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_83_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_84_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_85_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_86_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_87_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_88_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_89_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_90_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_91_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_92_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_93_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_94_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_95_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_96_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_97_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_98_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_99_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_100_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_101_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_102_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_103_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_104_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_105_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_106_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_107_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_108_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_109_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_110_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_111_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_112_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_113_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_114_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_115_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_116_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_117_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_118_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_119_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_120_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_121_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_122_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_123_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_124_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_125_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_126_IS_INOUT = 0,         //enables the input bram also for output
    parameter [0:0] S_AXIS_BRAM_127_IS_INOUT = 0,         //enables the input bram also for output
    parameter [31:0] S_AXIS_BRAM_0_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_1_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_2_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_3_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_4_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_5_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_6_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_7_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_8_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_9_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_10_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_11_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_12_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_13_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_14_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_15_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_16_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_17_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_18_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_19_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_20_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_21_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_22_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_23_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_24_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_25_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_26_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_27_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_28_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_29_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_30_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_31_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_32_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_33_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_34_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_35_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_36_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_37_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_38_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_39_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_40_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_41_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_42_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_43_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_44_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_45_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_46_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_47_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_48_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_49_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_50_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_51_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_52_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_53_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_54_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_55_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_56_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_57_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_58_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_59_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_60_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_61_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_62_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_63_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_64_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_65_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_66_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_67_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_68_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_69_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_70_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_71_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_72_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_73_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_74_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_75_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_76_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_77_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_78_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_79_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_80_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_81_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_82_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_83_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_84_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_85_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_86_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_87_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_88_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_89_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_90_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_91_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_92_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_93_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_94_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_95_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_96_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_97_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_98_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_99_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_100_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_101_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_102_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_103_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_104_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_105_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_106_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_107_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_108_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_109_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_110_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_111_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_112_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_113_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_114_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_115_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_116_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_117_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_118_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_119_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_120_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_121_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_122_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_123_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_124_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_125_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_126_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter [31:0] S_AXIS_BRAM_127_MB_DEPTH = 1,  //depth, number of copies of BRAM args
    parameter M_AXIS_BRAM_0_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_1_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_2_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_3_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_4_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_5_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_6_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_7_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_8_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_9_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_10_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_11_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_12_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_13_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_14_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_15_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_16_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_17_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_18_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_19_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_20_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_21_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_22_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_23_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_24_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_25_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_26_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_27_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_28_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_29_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_30_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_31_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_32_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_33_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_34_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_35_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_36_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_37_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_38_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_39_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_40_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_41_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_42_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_43_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_44_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_45_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_46_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_47_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_48_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_49_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_50_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_51_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_52_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_53_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_54_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_55_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_56_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_57_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_58_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_59_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_60_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_61_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_62_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_63_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_64_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_65_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_66_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_67_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_68_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_69_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_70_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_71_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_72_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_73_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_74_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_75_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_76_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_77_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_78_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_79_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_80_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_81_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_82_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_83_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_84_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_85_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_86_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_87_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_88_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_89_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_90_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_91_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_92_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_93_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_94_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_95_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_96_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_97_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_98_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_99_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_100_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_101_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_102_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_103_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_104_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_105_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_106_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_107_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_108_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_109_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_110_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_111_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_112_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_113_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_114_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_115_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_116_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_117_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_118_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_119_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_120_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_121_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_122_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_123_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_124_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_125_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_126_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter M_AXIS_BRAM_127_PORTS = 1,           //number of bram ports (dual-ported, partitioned)
    parameter [31:0] M_AXIS_BRAM_0_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_1_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_2_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_3_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_4_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_5_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_6_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_7_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_8_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_9_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_10_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_11_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_12_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_13_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_14_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_15_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_16_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_17_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_18_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_19_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_20_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_21_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_22_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_23_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_24_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_25_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_26_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_27_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_28_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_29_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_30_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_31_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_32_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_33_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_34_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_35_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_36_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_37_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_38_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_39_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_40_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_41_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_42_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_43_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_44_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_45_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_46_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_47_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_48_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_49_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_50_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_51_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_52_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_53_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_54_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_55_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_56_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_57_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_58_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_59_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_60_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_61_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_62_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_63_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_64_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_65_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_66_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_67_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_68_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_69_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_70_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_71_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_72_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_73_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_74_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_75_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_76_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_77_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_78_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_79_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_80_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_81_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_82_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_83_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_84_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_85_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_86_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_87_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_88_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_89_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_90_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_91_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_92_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_93_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_94_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_95_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_96_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_97_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_98_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_99_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_100_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_101_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_102_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_103_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_104_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_105_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_106_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_107_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_108_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_109_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_110_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_111_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_112_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_113_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_114_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_115_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_116_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_117_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_118_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_119_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_120_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_121_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_122_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_123_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_124_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_125_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_126_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_127_WIDTH = 8,    //width of output bram interface on the accelerator
    parameter [31:0] M_AXIS_BRAM_0_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_1_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_2_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_3_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_4_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_5_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_6_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_7_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_8_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_9_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_10_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_11_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_12_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_13_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_14_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_15_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_16_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_17_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_18_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_19_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_20_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_21_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_22_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_23_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_24_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_25_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_26_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_27_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_28_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_29_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_30_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_31_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_32_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_33_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_34_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_35_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_36_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_37_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_38_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_39_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_40_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_41_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_42_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_43_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_44_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_45_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_46_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_47_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_48_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_49_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_50_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_51_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_52_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_53_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_54_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_55_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_56_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_57_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_58_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_59_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_60_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_61_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_62_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_63_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_64_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_65_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_66_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_67_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_68_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_69_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_70_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_71_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_72_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_73_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_74_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_75_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_76_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_77_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_78_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_79_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_80_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_81_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_82_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_83_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_84_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_85_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_86_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_87_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_88_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_89_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_90_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_91_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_92_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_93_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_94_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_95_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_96_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_97_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_98_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_99_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_100_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_101_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_102_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_103_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_104_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_105_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_106_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_107_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_108_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_109_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_110_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_111_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_112_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_113_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_114_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_115_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_116_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_117_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_118_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_119_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_120_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_121_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_122_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_123_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_124_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_125_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_126_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_127_DEPTH = 2,    //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_0_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_1_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_2_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_3_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_4_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_5_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_6_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_7_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_8_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_9_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_10_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_11_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_12_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_13_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_14_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_15_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_16_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_17_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_18_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_19_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_20_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_21_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_22_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_23_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_24_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_25_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_26_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_27_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_28_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_29_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_30_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_31_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_32_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_33_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_34_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_35_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_36_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_37_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_38_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_39_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_40_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_41_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_42_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_43_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_44_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_45_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_46_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_47_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_48_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_49_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_50_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_51_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_52_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_53_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_54_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_55_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_56_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_57_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_58_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_59_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_60_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_61_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_62_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_63_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_64_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_65_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_66_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_67_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_68_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_69_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_70_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_71_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_72_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_73_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_74_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_75_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_76_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_77_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_78_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_79_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_80_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_81_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_82_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_83_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_84_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_85_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_86_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_87_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_88_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_89_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_90_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_91_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_92_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_93_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_94_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_95_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_96_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_97_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_98_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_99_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_100_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_101_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_102_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_103_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_104_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_105_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_106_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_107_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_108_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_109_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_110_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_111_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_112_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_113_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_114_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_115_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_116_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_117_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_118_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_119_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_120_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_121_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_122_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_123_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_124_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_125_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_126_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_127_DMWIDTH = 8,  //width of AXIS interface from adapter to DM for output bram interface
    parameter [31:0] M_AXIS_BRAM_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_BRAM_0_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_1_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_2_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_3_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_4_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_5_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_6_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_7_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_8_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_9_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_10_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_11_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_12_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_13_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_14_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_15_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_16_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_17_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_18_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_19_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_20_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_21_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_22_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_23_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_24_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_25_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_26_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_27_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_28_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_29_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_30_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_31_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_32_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_33_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_34_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_35_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_36_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_37_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_38_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_39_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_40_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_41_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_42_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_43_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_44_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_45_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_46_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_47_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_48_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_49_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_50_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_51_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_52_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_53_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_54_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_55_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_56_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_57_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_58_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_59_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_60_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_61_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_62_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_63_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_64_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_65_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_66_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_67_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_68_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_69_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_70_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_71_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_72_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_73_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_74_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_75_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_76_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_77_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_78_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_79_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_80_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_81_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_82_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_83_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_84_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_85_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_86_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_87_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_88_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_89_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_90_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_91_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_92_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_93_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_94_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_95_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_96_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_97_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_98_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_99_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_100_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_101_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_102_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_103_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_104_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_105_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_106_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_107_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_108_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_109_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_110_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_111_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_112_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_113_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_114_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_115_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_116_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_117_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_118_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_119_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_120_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_121_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_122_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_123_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_124_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_125_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_126_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    parameter [31:0] M_AXIS_BRAM_127_MB_DEPTH = 1, //depth of BRAM in adapter for output bram interface
    
    parameter S_AXIS_BRAM_0_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_1_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_2_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_3_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_4_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_5_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_6_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_7_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_8_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_9_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_10_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_11_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_12_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_13_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_14_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_15_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_16_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_17_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_18_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_19_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_20_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_21_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_22_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_23_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_24_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_25_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_26_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_27_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_28_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_29_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_30_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_31_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_32_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_33_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_34_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_35_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_36_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_37_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_38_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_39_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_40_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_41_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_42_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_43_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_44_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_45_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_46_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_47_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_48_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_49_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_50_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_51_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_52_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_53_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_54_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_55_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_56_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_57_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_58_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_59_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_60_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_61_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_62_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_63_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_64_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_65_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_66_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_67_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_68_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_69_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_70_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_71_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_72_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_73_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_74_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_75_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_76_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_77_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_78_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_79_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_80_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_81_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_82_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_83_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_84_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_85_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_86_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_87_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_88_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_89_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_90_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_91_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_92_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_93_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_94_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_95_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_96_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_97_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_98_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_99_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_100_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_101_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_102_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_103_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_104_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_105_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_106_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_107_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_108_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_109_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_110_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_111_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_112_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_113_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_114_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_115_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_116_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_117_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_118_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_119_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_120_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_121_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_122_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_123_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_124_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_125_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_126_ADDR_WIDTH = 1,
    parameter S_AXIS_BRAM_127_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_0_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_1_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_2_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_3_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_4_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_5_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_6_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_7_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_8_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_9_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_10_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_11_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_12_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_13_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_14_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_15_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_16_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_17_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_18_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_19_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_20_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_21_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_22_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_23_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_24_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_25_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_26_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_27_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_28_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_29_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_30_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_31_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_32_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_33_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_34_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_35_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_36_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_37_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_38_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_39_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_40_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_41_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_42_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_43_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_44_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_45_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_46_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_47_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_48_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_49_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_50_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_51_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_52_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_53_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_54_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_55_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_56_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_57_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_58_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_59_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_60_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_61_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_62_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_63_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_64_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_65_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_66_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_67_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_68_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_69_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_70_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_71_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_72_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_73_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_74_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_75_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_76_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_77_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_78_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_79_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_80_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_81_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_82_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_83_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_84_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_85_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_86_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_87_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_88_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_89_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_90_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_91_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_92_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_93_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_94_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_95_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_96_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_97_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_98_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_99_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_100_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_101_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_102_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_103_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_104_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_105_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_106_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_107_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_108_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_109_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_110_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_111_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_112_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_113_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_114_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_115_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_116_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_117_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_118_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_119_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_120_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_121_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_122_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_123_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_124_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_125_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_126_ADDR_WIDTH = 1,
    parameter M_AXIS_BRAM_127_ADDR_WIDTH = 1,
    //axis arg parameters
    parameter C_NUM_INPUT_AXISs = 0,                //number of input fifo interfaces on the accelerator
    parameter C_NUM_OUTPUT_AXISs = 0,               //number of output fifo interfaces on the accelerator
    parameter [31:0] S_AXIS_IARG_0_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_1_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_2_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_3_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_4_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_5_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_6_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_7_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_8_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_9_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_10_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_11_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_12_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_13_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_14_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_15_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_16_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_17_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_18_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_19_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_20_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_21_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_22_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_23_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_24_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_25_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_26_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_27_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_28_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_29_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_30_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_31_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_32_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_33_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_34_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_35_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_36_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_37_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_38_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_39_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_40_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_41_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_42_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_43_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_44_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_45_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_46_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_47_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_48_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_49_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_50_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_51_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_52_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_53_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_54_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_55_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_56_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_57_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_58_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_59_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_60_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_61_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_62_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_63_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_64_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_65_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_66_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_67_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_68_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_69_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_70_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_71_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_72_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_73_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_74_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_75_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_76_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_77_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_78_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_79_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_80_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_81_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_82_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_83_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_84_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_85_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_86_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_87_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_88_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_89_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_90_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_91_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_92_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_93_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_94_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_95_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_96_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_97_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_98_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_99_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_100_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_101_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_102_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_103_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_104_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_105_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_106_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_107_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_108_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_109_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_110_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_111_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_112_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_113_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_114_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_115_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_116_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_117_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_118_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_119_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_120_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_121_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_122_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_123_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_124_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_125_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_126_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_127_WIDTH = 8,     //width of input AXIS interface on the accelerator
    parameter [31:0] S_AXIS_IARG_0_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_1_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_2_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_3_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_4_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_5_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_6_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_7_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_8_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_9_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_10_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_11_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_12_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_13_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_14_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_15_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_16_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_17_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_18_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_19_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_20_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_21_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_22_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_23_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_24_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_25_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_26_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_27_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_28_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_29_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_30_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_31_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_32_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_33_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_34_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_35_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_36_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_37_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_38_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_39_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_40_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_41_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_42_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_43_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_44_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_45_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_46_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_47_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_48_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_49_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_50_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_51_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_52_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_53_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_54_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_55_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_56_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_57_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_58_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_59_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_60_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_61_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_62_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_63_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_64_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_65_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_66_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_67_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_68_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_69_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_70_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_71_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_72_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_73_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_74_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_75_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_76_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_77_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_78_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_79_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_80_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_81_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_82_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_83_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_84_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_85_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_86_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_87_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_88_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_89_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_90_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_91_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_92_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_93_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_94_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_95_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_96_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_97_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_98_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_99_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_100_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_101_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_102_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_103_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_104_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_105_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_106_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_107_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_108_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_109_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_110_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_111_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_112_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_113_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_114_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_115_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_116_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_117_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_118_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_119_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_120_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_121_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_122_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_123_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_124_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_125_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_126_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_127_DEPTH = 16,      //depth of AXIS in adapter for input AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] S_AXIS_IARG_0_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_1_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_2_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_3_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_4_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_5_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_6_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_7_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_8_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_9_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_10_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_11_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_12_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_13_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_14_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_15_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_16_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_17_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_18_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_19_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_20_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_21_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_22_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_23_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_24_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_25_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_26_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_27_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_28_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_29_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_30_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_31_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_32_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_33_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_34_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_35_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_36_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_37_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_38_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_39_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_40_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_41_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_42_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_43_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_44_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_45_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_46_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_47_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_48_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_49_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_50_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_51_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_52_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_53_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_54_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_55_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_56_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_57_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_58_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_59_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_60_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_61_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_62_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_63_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_64_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_65_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_66_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_67_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_68_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_69_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_70_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_71_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_72_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_73_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_74_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_75_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_76_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_77_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_78_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_79_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_80_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_81_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_82_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_83_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_84_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_85_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_86_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_87_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_88_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_89_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_90_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_91_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_92_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_93_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_94_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_95_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_96_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_97_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_98_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_99_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_100_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_101_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_102_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_103_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_104_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_105_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_106_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_107_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_108_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_109_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_110_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_111_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_112_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_113_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_114_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_115_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_116_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_117_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_118_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_119_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_120_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_121_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_122_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_123_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_124_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_125_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_126_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_127_DMWIDTH = 8,   //width of AXIS interface from DM to adapter for input AXIS interface
    parameter [31:0] S_AXIS_IARG_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] S_AXIS_IARG_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_0_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_1_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_2_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_3_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_4_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_5_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_6_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_7_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_8_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_9_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_10_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_11_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_12_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_13_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_14_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_15_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_16_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_17_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_18_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_19_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_20_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_21_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_22_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_23_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_24_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_25_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_26_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_27_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_28_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_29_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_30_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_31_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_32_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_33_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_34_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_35_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_36_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_37_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_38_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_39_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_40_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_41_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_42_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_43_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_44_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_45_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_46_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_47_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_48_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_49_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_50_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_51_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_52_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_53_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_54_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_55_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_56_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_57_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_58_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_59_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_60_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_61_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_62_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_63_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_64_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_65_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_66_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_67_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_68_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_69_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_70_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_71_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_72_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_73_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_74_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_75_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_76_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_77_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_78_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_79_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_80_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_81_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_82_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_83_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_84_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_85_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_86_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_87_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_88_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_89_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_90_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_91_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_92_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_93_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_94_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_95_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_96_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_97_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_98_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_99_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_100_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_101_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_102_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_103_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_104_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_105_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_106_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_107_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_108_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_109_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_110_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_111_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_112_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_113_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_114_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_115_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_116_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_117_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_118_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_119_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_120_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_121_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_122_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_123_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_124_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_125_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_126_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_127_WIDTH = 8,    //width of output AXIS interface on the accelerator
    parameter [31:0] M_AXIS_OARG_0_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_1_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_2_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_3_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_4_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_5_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_6_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_7_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_8_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_9_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_10_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_11_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_12_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_13_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_14_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_15_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_16_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_17_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_18_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_19_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_20_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_21_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_22_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_23_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_24_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_25_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_26_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_27_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_28_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_29_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_30_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_31_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_32_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_33_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_34_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_35_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_36_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_37_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_38_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_39_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_40_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_41_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_42_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_43_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_44_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_45_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_46_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_47_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_48_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_49_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_50_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_51_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_52_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_53_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_54_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_55_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_56_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_57_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_58_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_59_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_60_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_61_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_62_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_63_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_64_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_65_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_66_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_67_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_68_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_69_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_70_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_71_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_72_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_73_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_74_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_75_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_76_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_77_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_78_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_79_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_80_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_81_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_82_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_83_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_84_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_85_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_86_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_87_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_88_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_89_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_90_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_91_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_92_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_93_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_94_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_95_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_96_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_97_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_98_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_99_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_100_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_101_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_102_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_103_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_104_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_105_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_106_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_107_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_108_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_109_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_110_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_111_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_112_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_113_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_114_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_115_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_116_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_117_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_118_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_119_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_120_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_121_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_122_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_123_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_124_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_125_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_126_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_127_DEPTH = 16,     //depth of AXIS in adapter for output AXIS interface (minimum value 1, required for clock conversion)
    parameter [31:0] M_AXIS_OARG_0_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_1_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_2_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_3_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_4_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_5_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_6_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_7_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_8_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_9_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_10_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_11_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_12_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_13_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_14_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_15_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_16_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_17_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_18_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_19_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_20_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_21_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_22_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_23_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_24_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_25_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_26_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_27_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_28_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_29_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_30_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_31_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_32_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_33_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_34_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_35_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_36_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_37_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_38_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_39_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_40_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_41_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_42_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_43_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_44_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_45_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_46_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_47_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_48_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_49_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_50_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_51_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_52_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_53_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_54_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_55_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_56_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_57_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_58_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_59_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_60_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_61_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_62_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_63_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_64_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_65_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_66_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_67_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_68_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_69_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_70_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_71_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_72_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_73_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_74_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_75_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_76_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_77_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_78_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_79_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_80_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_81_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_82_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_83_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_84_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_85_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_86_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_87_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_88_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_89_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_90_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_91_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_92_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_93_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_94_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_95_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_96_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_97_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_98_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_99_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_100_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_101_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_102_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_103_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_104_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_105_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_106_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_107_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_108_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_109_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_110_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_111_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_112_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_113_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_114_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_115_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_116_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_117_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_118_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_119_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_120_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_121_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_122_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_123_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_124_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_125_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_126_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_127_DMWIDTH = 8,  //width of AXIS interface from DM to adapter for output AXIS interface
    parameter [31:0] M_AXIS_OARG_0_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_1_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_2_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_3_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_4_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_5_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_6_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_7_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_8_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_9_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_10_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_11_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_12_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_13_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_14_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_15_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_16_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_17_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_18_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_19_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_20_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_21_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_22_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_23_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_24_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_25_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_26_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_27_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_28_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_29_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_30_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_31_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_32_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_33_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_34_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_35_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_36_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_37_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_38_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_39_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_40_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_41_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_42_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_43_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_44_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_45_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_46_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_47_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_48_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_49_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_50_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_51_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_52_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_53_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_54_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_55_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_56_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_57_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_58_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_59_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_60_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_61_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_62_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_63_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_64_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_65_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_66_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_67_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_68_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_69_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_70_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_71_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_72_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_73_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_74_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_75_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_76_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_77_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_78_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_79_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_80_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_81_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_82_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_83_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_84_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_85_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_86_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_87_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_88_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_89_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_90_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_91_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_92_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_93_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_94_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_95_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_96_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_97_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_98_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_99_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_100_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_101_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_102_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_103_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_104_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_105_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_106_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_107_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_108_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_109_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_110_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_111_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_112_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_113_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_114_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_115_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_116_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_117_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_118_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_119_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_120_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_121_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_122_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_123_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_124_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_125_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_126_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_127_IS_ASYNC = 0,  //should fifo buffer be asynchronous (0) or synchronours (1)
    parameter [31:0] M_AXIS_OARG_0_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_1_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_2_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_3_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_4_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_5_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_6_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_7_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_8_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_9_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_10_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_11_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_12_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_13_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_14_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_15_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_16_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_17_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_18_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_19_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_20_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_21_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_22_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_23_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_24_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_25_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_26_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_27_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_28_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_29_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_30_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_31_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_32_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_33_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_34_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_35_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_36_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_37_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_38_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_39_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_40_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_41_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_42_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_43_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_44_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_45_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_46_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_47_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_48_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_49_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_50_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_51_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_52_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_53_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_54_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_55_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_56_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_57_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_58_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_59_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_60_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_61_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_62_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_63_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_64_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_65_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_66_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_67_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_68_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_69_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_70_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_71_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_72_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_73_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_74_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_75_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_76_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_77_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_78_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_79_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_80_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_81_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_82_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_83_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_84_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_85_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_86_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_87_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_88_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_89_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_90_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_91_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_92_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_93_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_94_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_95_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_96_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_97_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_98_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_99_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_100_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_101_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_102_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_103_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_104_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_105_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_106_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_107_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_108_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_109_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_110_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_111_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_112_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_113_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_114_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_115_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_116_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_117_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_118_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_119_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_120_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_121_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_122_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_123_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_124_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_125_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_126_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    parameter [31:0] M_AXIS_OARG_127_GEN_TLAST = 0,  //generate TLAST signal for output AXIS interface
    //aximm arg parameters
    parameter C_NUM_AXIMMs = 0,                //number of aximm interfaces on the accelerator
    parameter M_AXIMM_ADDR_WIDTH = 32,
    parameter M_AXIMM_0_DATA_WIDTH = 32,
    parameter M_AXIMM_1_DATA_WIDTH = 32,
    parameter M_AXIMM_2_DATA_WIDTH = 32,
    parameter M_AXIMM_3_DATA_WIDTH = 32,
    parameter M_AXIMM_4_DATA_WIDTH = 32,
    parameter M_AXIMM_5_DATA_WIDTH = 32,
    parameter M_AXIMM_6_DATA_WIDTH = 32,
    parameter M_AXIMM_7_DATA_WIDTH = 32,
    parameter M_AXIMM_8_DATA_WIDTH = 32,
    parameter M_AXIMM_9_DATA_WIDTH = 32,
    parameter M_AXIMM_10_DATA_WIDTH = 32,
    parameter M_AXIMM_11_DATA_WIDTH = 32,
    parameter M_AXIMM_12_DATA_WIDTH = 32,
    parameter M_AXIMM_13_DATA_WIDTH = 32,
    parameter M_AXIMM_14_DATA_WIDTH = 32,
    parameter M_AXIMM_15_DATA_WIDTH = 32,
    parameter M_AXIMM_16_DATA_WIDTH = 32,
    parameter M_AXIMM_17_DATA_WIDTH = 32,
    parameter M_AXIMM_18_DATA_WIDTH = 32,
    parameter M_AXIMM_19_DATA_WIDTH = 32,
    parameter M_AXIMM_20_DATA_WIDTH = 32,
    parameter M_AXIMM_21_DATA_WIDTH = 32,
    parameter M_AXIMM_22_DATA_WIDTH = 32,
    parameter M_AXIMM_23_DATA_WIDTH = 32,
    parameter M_AXIMM_24_DATA_WIDTH = 32,
    parameter M_AXIMM_25_DATA_WIDTH = 32,
    parameter M_AXIMM_26_DATA_WIDTH = 32,
    parameter M_AXIMM_27_DATA_WIDTH = 32,
    parameter M_AXIMM_28_DATA_WIDTH = 32,
    parameter M_AXIMM_29_DATA_WIDTH = 32,
    parameter M_AXIMM_30_DATA_WIDTH = 32,
    parameter M_AXIMM_31_DATA_WIDTH = 32,
    parameter M_AXIMM_32_DATA_WIDTH = 32,
    parameter M_AXIMM_33_DATA_WIDTH = 32,
    parameter M_AXIMM_34_DATA_WIDTH = 32,
    parameter M_AXIMM_35_DATA_WIDTH = 32,
    parameter M_AXIMM_36_DATA_WIDTH = 32,
    parameter M_AXIMM_37_DATA_WIDTH = 32,
    parameter M_AXIMM_38_DATA_WIDTH = 32,
    parameter M_AXIMM_39_DATA_WIDTH = 32,
    parameter M_AXIMM_40_DATA_WIDTH = 32,
    parameter M_AXIMM_41_DATA_WIDTH = 32,
    parameter M_AXIMM_42_DATA_WIDTH = 32,
    parameter M_AXIMM_43_DATA_WIDTH = 32,
    parameter M_AXIMM_44_DATA_WIDTH = 32,
    parameter M_AXIMM_45_DATA_WIDTH = 32,
    parameter M_AXIMM_46_DATA_WIDTH = 32,
    parameter M_AXIMM_47_DATA_WIDTH = 32,
    parameter M_AXIMM_48_DATA_WIDTH = 32,
    parameter M_AXIMM_49_DATA_WIDTH = 32,
    parameter M_AXIMM_50_DATA_WIDTH = 32,
    parameter M_AXIMM_51_DATA_WIDTH = 32,
    parameter M_AXIMM_52_DATA_WIDTH = 32,
    parameter M_AXIMM_53_DATA_WIDTH = 32,
    parameter M_AXIMM_54_DATA_WIDTH = 32,
    parameter M_AXIMM_55_DATA_WIDTH = 32,
    parameter M_AXIMM_56_DATA_WIDTH = 32,
    parameter M_AXIMM_57_DATA_WIDTH = 32,
    parameter M_AXIMM_58_DATA_WIDTH = 32,
    parameter M_AXIMM_59_DATA_WIDTH = 32,
    parameter M_AXIMM_60_DATA_WIDTH = 32,
    parameter M_AXIMM_61_DATA_WIDTH = 32,
    parameter M_AXIMM_62_DATA_WIDTH = 32,
    parameter M_AXIMM_63_DATA_WIDTH = 32,
    parameter M_AXIMM_64_DATA_WIDTH = 32,
    parameter M_AXIMM_65_DATA_WIDTH = 32,
    parameter M_AXIMM_66_DATA_WIDTH = 32,
    parameter M_AXIMM_67_DATA_WIDTH = 32,
    parameter M_AXIMM_68_DATA_WIDTH = 32,
    parameter M_AXIMM_69_DATA_WIDTH = 32,
    parameter M_AXIMM_70_DATA_WIDTH = 32,
    parameter M_AXIMM_71_DATA_WIDTH = 32,
    parameter M_AXIMM_72_DATA_WIDTH = 32,
    parameter M_AXIMM_73_DATA_WIDTH = 32,
    parameter M_AXIMM_74_DATA_WIDTH = 32,
    parameter M_AXIMM_75_DATA_WIDTH = 32,
    parameter M_AXIMM_76_DATA_WIDTH = 32,
    parameter M_AXIMM_77_DATA_WIDTH = 32,
    parameter M_AXIMM_78_DATA_WIDTH = 32,
    parameter M_AXIMM_79_DATA_WIDTH = 32,
    parameter M_AXIMM_80_DATA_WIDTH = 32,
    parameter M_AXIMM_81_DATA_WIDTH = 32,
    parameter M_AXIMM_82_DATA_WIDTH = 32,
    parameter M_AXIMM_83_DATA_WIDTH = 32,
    parameter M_AXIMM_84_DATA_WIDTH = 32,
    parameter M_AXIMM_85_DATA_WIDTH = 32,
    parameter M_AXIMM_86_DATA_WIDTH = 32,
    parameter M_AXIMM_87_DATA_WIDTH = 32,
    parameter M_AXIMM_88_DATA_WIDTH = 32,
    parameter M_AXIMM_89_DATA_WIDTH = 32,
    parameter M_AXIMM_90_DATA_WIDTH = 32,
    parameter M_AXIMM_91_DATA_WIDTH = 32,
    parameter M_AXIMM_92_DATA_WIDTH = 32,
    parameter M_AXIMM_93_DATA_WIDTH = 32,
    parameter M_AXIMM_94_DATA_WIDTH = 32,
    parameter M_AXIMM_95_DATA_WIDTH = 32,
    parameter M_AXIMM_96_DATA_WIDTH = 32,
    parameter M_AXIMM_97_DATA_WIDTH = 32,
    parameter M_AXIMM_98_DATA_WIDTH = 32,
    parameter M_AXIMM_99_DATA_WIDTH = 32,
    parameter M_AXIMM_100_DATA_WIDTH = 32,
    parameter M_AXIMM_101_DATA_WIDTH = 32,
    parameter M_AXIMM_102_DATA_WIDTH = 32,
    parameter M_AXIMM_103_DATA_WIDTH = 32,
    parameter M_AXIMM_104_DATA_WIDTH = 32,
    parameter M_AXIMM_105_DATA_WIDTH = 32,
    parameter M_AXIMM_106_DATA_WIDTH = 32,
    parameter M_AXIMM_107_DATA_WIDTH = 32,
    parameter M_AXIMM_108_DATA_WIDTH = 32,
    parameter M_AXIMM_109_DATA_WIDTH = 32,
    parameter M_AXIMM_110_DATA_WIDTH = 32,
    parameter M_AXIMM_111_DATA_WIDTH = 32,
    parameter M_AXIMM_112_DATA_WIDTH = 32,
    parameter M_AXIMM_113_DATA_WIDTH = 32,
    parameter M_AXIMM_114_DATA_WIDTH = 32,
    parameter M_AXIMM_115_DATA_WIDTH = 32,
    parameter M_AXIMM_116_DATA_WIDTH = 32,
    parameter M_AXIMM_117_DATA_WIDTH = 32,
    parameter M_AXIMM_118_DATA_WIDTH = 32,
    parameter M_AXIMM_119_DATA_WIDTH = 32,
    parameter M_AXIMM_120_DATA_WIDTH = 32,
    parameter M_AXIMM_121_DATA_WIDTH = 32,
    parameter M_AXIMM_122_DATA_WIDTH = 32,
    parameter M_AXIMM_123_DATA_WIDTH = 32,
    parameter M_AXIMM_124_DATA_WIDTH = 32,
    parameter M_AXIMM_125_DATA_WIDTH = 32,
    parameter M_AXIMM_126_DATA_WIDTH = 32,
    parameter M_AXIMM_127_DATA_WIDTH = 32,
    parameter [0:0] M_AXIMM_0_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_WID_WIDTH = 0
 ) (
    //axi lite interface
    input s_axi_aclk,
    input s_axi_aresetn,
    input [31 : 0] S_AXI_AWADDR,
    input [2 : 0] S_AXI_AWPROT,
    input S_AXI_AWVALID,
    output S_AXI_AWREADY,
    input [31 : 0] S_AXI_WDATA,
    input [3 : 0] S_AXI_WSTRB,
    input S_AXI_WVALID,
    output S_AXI_WREADY,
    output [1 : 0] S_AXI_BRESP,
    output S_AXI_BVALID,
    input S_AXI_BREADY,
    input [31 : 0] S_AXI_ARADDR,
    input [2 : 0] S_AXI_ARPROT,
    input S_AXI_ARVALID,
    output S_AXI_ARREADY,
    output [31 : 0] S_AXI_RDATA,
    output [1 : 0] S_AXI_RRESP,
    output S_AXI_RVALID,
    input S_AXI_RREADY,
    //acc clock
    input acc_aclk,
    input acc_aresetn,
    //acc interface
    output ap_resetn,
    output ap_clk,
    output ap_start,
    input ap_idle,
    input ap_done,
    input ap_ready,
    output ap_continue,
    //-----------------------------------------------------
    //input scalar ports
    output [C_INPUT_SCALAR_0_WIDTH-1:0] ap_iscalar_0_dout,
    output [C_INPUT_SCALAR_1_WIDTH-1:0] ap_iscalar_1_dout,
    output [C_INPUT_SCALAR_2_WIDTH-1:0] ap_iscalar_2_dout,
    output [C_INPUT_SCALAR_3_WIDTH-1:0] ap_iscalar_3_dout,
    output [C_INPUT_SCALAR_4_WIDTH-1:0] ap_iscalar_4_dout,
    output [C_INPUT_SCALAR_5_WIDTH-1:0] ap_iscalar_5_dout,
    output [C_INPUT_SCALAR_6_WIDTH-1:0] ap_iscalar_6_dout,
    output [C_INPUT_SCALAR_7_WIDTH-1:0] ap_iscalar_7_dout,
    output [C_INPUT_SCALAR_8_WIDTH-1:0] ap_iscalar_8_dout,
    output [C_INPUT_SCALAR_9_WIDTH-1:0] ap_iscalar_9_dout,
    output [C_INPUT_SCALAR_10_WIDTH-1:0] ap_iscalar_10_dout,
    output [C_INPUT_SCALAR_11_WIDTH-1:0] ap_iscalar_11_dout,
    output [C_INPUT_SCALAR_12_WIDTH-1:0] ap_iscalar_12_dout,
    output [C_INPUT_SCALAR_13_WIDTH-1:0] ap_iscalar_13_dout,
    output [C_INPUT_SCALAR_14_WIDTH-1:0] ap_iscalar_14_dout,
    output [C_INPUT_SCALAR_15_WIDTH-1:0] ap_iscalar_15_dout,
    output [C_INPUT_SCALAR_16_WIDTH-1:0] ap_iscalar_16_dout,
    output [C_INPUT_SCALAR_17_WIDTH-1:0] ap_iscalar_17_dout,
    output [C_INPUT_SCALAR_18_WIDTH-1:0] ap_iscalar_18_dout,
    output [C_INPUT_SCALAR_19_WIDTH-1:0] ap_iscalar_19_dout,
    output [C_INPUT_SCALAR_20_WIDTH-1:0] ap_iscalar_20_dout,
    output [C_INPUT_SCALAR_21_WIDTH-1:0] ap_iscalar_21_dout,
    output [C_INPUT_SCALAR_22_WIDTH-1:0] ap_iscalar_22_dout,
    output [C_INPUT_SCALAR_23_WIDTH-1:0] ap_iscalar_23_dout,
    output [C_INPUT_SCALAR_24_WIDTH-1:0] ap_iscalar_24_dout,
    output [C_INPUT_SCALAR_25_WIDTH-1:0] ap_iscalar_25_dout,
    output [C_INPUT_SCALAR_26_WIDTH-1:0] ap_iscalar_26_dout,
    output [C_INPUT_SCALAR_27_WIDTH-1:0] ap_iscalar_27_dout,
    output [C_INPUT_SCALAR_28_WIDTH-1:0] ap_iscalar_28_dout,
    output [C_INPUT_SCALAR_29_WIDTH-1:0] ap_iscalar_29_dout,
    output [C_INPUT_SCALAR_30_WIDTH-1:0] ap_iscalar_30_dout,
    output [C_INPUT_SCALAR_31_WIDTH-1:0] ap_iscalar_31_dout,
    output [C_INPUT_SCALAR_32_WIDTH-1:0] ap_iscalar_32_dout,
    output [C_INPUT_SCALAR_33_WIDTH-1:0] ap_iscalar_33_dout,
    output [C_INPUT_SCALAR_34_WIDTH-1:0] ap_iscalar_34_dout,
    output [C_INPUT_SCALAR_35_WIDTH-1:0] ap_iscalar_35_dout,
    output [C_INPUT_SCALAR_36_WIDTH-1:0] ap_iscalar_36_dout,
    output [C_INPUT_SCALAR_37_WIDTH-1:0] ap_iscalar_37_dout,
    output [C_INPUT_SCALAR_38_WIDTH-1:0] ap_iscalar_38_dout,
    output [C_INPUT_SCALAR_39_WIDTH-1:0] ap_iscalar_39_dout,
    output [C_INPUT_SCALAR_40_WIDTH-1:0] ap_iscalar_40_dout,
    output [C_INPUT_SCALAR_41_WIDTH-1:0] ap_iscalar_41_dout,
    output [C_INPUT_SCALAR_42_WIDTH-1:0] ap_iscalar_42_dout,
    output [C_INPUT_SCALAR_43_WIDTH-1:0] ap_iscalar_43_dout,
    output [C_INPUT_SCALAR_44_WIDTH-1:0] ap_iscalar_44_dout,
    output [C_INPUT_SCALAR_45_WIDTH-1:0] ap_iscalar_45_dout,
    output [C_INPUT_SCALAR_46_WIDTH-1:0] ap_iscalar_46_dout,
    output [C_INPUT_SCALAR_47_WIDTH-1:0] ap_iscalar_47_dout,
    output [C_INPUT_SCALAR_48_WIDTH-1:0] ap_iscalar_48_dout,
    output [C_INPUT_SCALAR_49_WIDTH-1:0] ap_iscalar_49_dout,
    output [C_INPUT_SCALAR_50_WIDTH-1:0] ap_iscalar_50_dout,
    output [C_INPUT_SCALAR_51_WIDTH-1:0] ap_iscalar_51_dout,
    output [C_INPUT_SCALAR_52_WIDTH-1:0] ap_iscalar_52_dout,
    output [C_INPUT_SCALAR_53_WIDTH-1:0] ap_iscalar_53_dout,
    output [C_INPUT_SCALAR_54_WIDTH-1:0] ap_iscalar_54_dout,
    output [C_INPUT_SCALAR_55_WIDTH-1:0] ap_iscalar_55_dout,
    output [C_INPUT_SCALAR_56_WIDTH-1:0] ap_iscalar_56_dout,
    output [C_INPUT_SCALAR_57_WIDTH-1:0] ap_iscalar_57_dout,
    output [C_INPUT_SCALAR_58_WIDTH-1:0] ap_iscalar_58_dout,
    output [C_INPUT_SCALAR_59_WIDTH-1:0] ap_iscalar_59_dout,
    output [C_INPUT_SCALAR_60_WIDTH-1:0] ap_iscalar_60_dout,
    output [C_INPUT_SCALAR_61_WIDTH-1:0] ap_iscalar_61_dout,
    output [C_INPUT_SCALAR_62_WIDTH-1:0] ap_iscalar_62_dout,
    output [C_INPUT_SCALAR_63_WIDTH-1:0] ap_iscalar_63_dout,
    output [C_INPUT_SCALAR_64_WIDTH-1:0] ap_iscalar_64_dout,
    output [C_INPUT_SCALAR_65_WIDTH-1:0] ap_iscalar_65_dout,
    output [C_INPUT_SCALAR_66_WIDTH-1:0] ap_iscalar_66_dout,
    output [C_INPUT_SCALAR_67_WIDTH-1:0] ap_iscalar_67_dout,
    output [C_INPUT_SCALAR_68_WIDTH-1:0] ap_iscalar_68_dout,
    output [C_INPUT_SCALAR_69_WIDTH-1:0] ap_iscalar_69_dout,
    output [C_INPUT_SCALAR_70_WIDTH-1:0] ap_iscalar_70_dout,
    output [C_INPUT_SCALAR_71_WIDTH-1:0] ap_iscalar_71_dout,
    output [C_INPUT_SCALAR_72_WIDTH-1:0] ap_iscalar_72_dout,
    output [C_INPUT_SCALAR_73_WIDTH-1:0] ap_iscalar_73_dout,
    output [C_INPUT_SCALAR_74_WIDTH-1:0] ap_iscalar_74_dout,
    output [C_INPUT_SCALAR_75_WIDTH-1:0] ap_iscalar_75_dout,
    output [C_INPUT_SCALAR_76_WIDTH-1:0] ap_iscalar_76_dout,
    output [C_INPUT_SCALAR_77_WIDTH-1:0] ap_iscalar_77_dout,
    output [C_INPUT_SCALAR_78_WIDTH-1:0] ap_iscalar_78_dout,
    output [C_INPUT_SCALAR_79_WIDTH-1:0] ap_iscalar_79_dout,
    output [C_INPUT_SCALAR_80_WIDTH-1:0] ap_iscalar_80_dout,
    output [C_INPUT_SCALAR_81_WIDTH-1:0] ap_iscalar_81_dout,
    output [C_INPUT_SCALAR_82_WIDTH-1:0] ap_iscalar_82_dout,
    output [C_INPUT_SCALAR_83_WIDTH-1:0] ap_iscalar_83_dout,
    output [C_INPUT_SCALAR_84_WIDTH-1:0] ap_iscalar_84_dout,
    output [C_INPUT_SCALAR_85_WIDTH-1:0] ap_iscalar_85_dout,
    output [C_INPUT_SCALAR_86_WIDTH-1:0] ap_iscalar_86_dout,
    output [C_INPUT_SCALAR_87_WIDTH-1:0] ap_iscalar_87_dout,
    output [C_INPUT_SCALAR_88_WIDTH-1:0] ap_iscalar_88_dout,
    output [C_INPUT_SCALAR_89_WIDTH-1:0] ap_iscalar_89_dout,
    output [C_INPUT_SCALAR_90_WIDTH-1:0] ap_iscalar_90_dout,
    output [C_INPUT_SCALAR_91_WIDTH-1:0] ap_iscalar_91_dout,
    output [C_INPUT_SCALAR_92_WIDTH-1:0] ap_iscalar_92_dout,
    output [C_INPUT_SCALAR_93_WIDTH-1:0] ap_iscalar_93_dout,
    output [C_INPUT_SCALAR_94_WIDTH-1:0] ap_iscalar_94_dout,
    output [C_INPUT_SCALAR_95_WIDTH-1:0] ap_iscalar_95_dout,
    output [C_INPUT_SCALAR_96_WIDTH-1:0] ap_iscalar_96_dout,
    output [C_INPUT_SCALAR_97_WIDTH-1:0] ap_iscalar_97_dout,
    output [C_INPUT_SCALAR_98_WIDTH-1:0] ap_iscalar_98_dout,
    output [C_INPUT_SCALAR_99_WIDTH-1:0] ap_iscalar_99_dout,
    output [C_INPUT_SCALAR_100_WIDTH-1:0] ap_iscalar_100_dout,
    output [C_INPUT_SCALAR_101_WIDTH-1:0] ap_iscalar_101_dout,
    output [C_INPUT_SCALAR_102_WIDTH-1:0] ap_iscalar_102_dout,
    output [C_INPUT_SCALAR_103_WIDTH-1:0] ap_iscalar_103_dout,
    output [C_INPUT_SCALAR_104_WIDTH-1:0] ap_iscalar_104_dout,
    output [C_INPUT_SCALAR_105_WIDTH-1:0] ap_iscalar_105_dout,
    output [C_INPUT_SCALAR_106_WIDTH-1:0] ap_iscalar_106_dout,
    output [C_INPUT_SCALAR_107_WIDTH-1:0] ap_iscalar_107_dout,
    output [C_INPUT_SCALAR_108_WIDTH-1:0] ap_iscalar_108_dout,
    output [C_INPUT_SCALAR_109_WIDTH-1:0] ap_iscalar_109_dout,
    output [C_INPUT_SCALAR_110_WIDTH-1:0] ap_iscalar_110_dout,
    output [C_INPUT_SCALAR_111_WIDTH-1:0] ap_iscalar_111_dout,
    output [C_INPUT_SCALAR_112_WIDTH-1:0] ap_iscalar_112_dout,
    output [C_INPUT_SCALAR_113_WIDTH-1:0] ap_iscalar_113_dout,
    output [C_INPUT_SCALAR_114_WIDTH-1:0] ap_iscalar_114_dout,
    output [C_INPUT_SCALAR_115_WIDTH-1:0] ap_iscalar_115_dout,
    output [C_INPUT_SCALAR_116_WIDTH-1:0] ap_iscalar_116_dout,
    output [C_INPUT_SCALAR_117_WIDTH-1:0] ap_iscalar_117_dout,
    output [C_INPUT_SCALAR_118_WIDTH-1:0] ap_iscalar_118_dout,
    output [C_INPUT_SCALAR_119_WIDTH-1:0] ap_iscalar_119_dout,
    output [C_INPUT_SCALAR_120_WIDTH-1:0] ap_iscalar_120_dout,
    output [C_INPUT_SCALAR_121_WIDTH-1:0] ap_iscalar_121_dout,
    output [C_INPUT_SCALAR_122_WIDTH-1:0] ap_iscalar_122_dout,
    output [C_INPUT_SCALAR_123_WIDTH-1:0] ap_iscalar_123_dout,
    output [C_INPUT_SCALAR_124_WIDTH-1:0] ap_iscalar_124_dout,
    output [C_INPUT_SCALAR_125_WIDTH-1:0] ap_iscalar_125_dout,
    output [C_INPUT_SCALAR_126_WIDTH-1:0] ap_iscalar_126_dout,
    output [C_INPUT_SCALAR_127_WIDTH-1:0] ap_iscalar_127_dout,
    //input scalar direct AXIS interfaces
    //input AXI-Stream to Scalar interface 0
    input s_axis_scalar_0_aclk,
    input s_axis_scalar_0_aresetn,
    input s_axis_scalar_0_tlast,
    input s_axis_scalar_0_tvalid,
    input [S_AXIS_SCALAR_0_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_0_tkeep,
    input [S_AXIS_SCALAR_0_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_0_tstrb,
    input [S_AXIS_SCALAR_0_DIRECT_DMWIDTH-1:0] s_axis_scalar_0_tdata,
    output s_axis_scalar_0_tready,
    //input AXI-Stream to Scalar interface 1
    input s_axis_scalar_1_aclk,
    input s_axis_scalar_1_aresetn,
    input s_axis_scalar_1_tlast,
    input s_axis_scalar_1_tvalid,
    input [S_AXIS_SCALAR_1_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_1_tkeep,
    input [S_AXIS_SCALAR_1_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_1_tstrb,
    input [S_AXIS_SCALAR_1_DIRECT_DMWIDTH-1:0] s_axis_scalar_1_tdata,
    output s_axis_scalar_1_tready,
    //input AXI-Stream to Scalar interface 2
    input s_axis_scalar_2_aclk,
    input s_axis_scalar_2_aresetn,
    input s_axis_scalar_2_tlast,
    input s_axis_scalar_2_tvalid,
    input [S_AXIS_SCALAR_2_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_2_tkeep,
    input [S_AXIS_SCALAR_2_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_2_tstrb,
    input [S_AXIS_SCALAR_2_DIRECT_DMWIDTH-1:0] s_axis_scalar_2_tdata,
    output s_axis_scalar_2_tready,
    //input AXI-Stream to Scalar interface 3
    input s_axis_scalar_3_aclk,
    input s_axis_scalar_3_aresetn,
    input s_axis_scalar_3_tlast,
    input s_axis_scalar_3_tvalid,
    input [S_AXIS_SCALAR_3_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_3_tkeep,
    input [S_AXIS_SCALAR_3_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_3_tstrb,
    input [S_AXIS_SCALAR_3_DIRECT_DMWIDTH-1:0] s_axis_scalar_3_tdata,
    output s_axis_scalar_3_tready,
    //input AXI-Stream to Scalar interface 4
    input s_axis_scalar_4_aclk,
    input s_axis_scalar_4_aresetn,
    input s_axis_scalar_4_tlast,
    input s_axis_scalar_4_tvalid,
    input [S_AXIS_SCALAR_4_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_4_tkeep,
    input [S_AXIS_SCALAR_4_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_4_tstrb,
    input [S_AXIS_SCALAR_4_DIRECT_DMWIDTH-1:0] s_axis_scalar_4_tdata,
    output s_axis_scalar_4_tready,
    //input AXI-Stream to Scalar interface 5
    input s_axis_scalar_5_aclk,
    input s_axis_scalar_5_aresetn,
    input s_axis_scalar_5_tlast,
    input s_axis_scalar_5_tvalid,
    input [S_AXIS_SCALAR_5_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_5_tkeep,
    input [S_AXIS_SCALAR_5_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_5_tstrb,
    input [S_AXIS_SCALAR_5_DIRECT_DMWIDTH-1:0] s_axis_scalar_5_tdata,
    output s_axis_scalar_5_tready,
    //input AXI-Stream to Scalar interface 6
    input s_axis_scalar_6_aclk,
    input s_axis_scalar_6_aresetn,
    input s_axis_scalar_6_tlast,
    input s_axis_scalar_6_tvalid,
    input [S_AXIS_SCALAR_6_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_6_tkeep,
    input [S_AXIS_SCALAR_6_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_6_tstrb,
    input [S_AXIS_SCALAR_6_DIRECT_DMWIDTH-1:0] s_axis_scalar_6_tdata,
    output s_axis_scalar_6_tready,
    //input AXI-Stream to Scalar interface 7
    input s_axis_scalar_7_aclk,
    input s_axis_scalar_7_aresetn,
    input s_axis_scalar_7_tlast,
    input s_axis_scalar_7_tvalid,
    input [S_AXIS_SCALAR_7_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_7_tkeep,
    input [S_AXIS_SCALAR_7_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_7_tstrb,
    input [S_AXIS_SCALAR_7_DIRECT_DMWIDTH-1:0] s_axis_scalar_7_tdata,
    output s_axis_scalar_7_tready,
    //input AXI-Stream to Scalar interface 8
    input s_axis_scalar_8_aclk,
    input s_axis_scalar_8_aresetn,
    input s_axis_scalar_8_tlast,
    input s_axis_scalar_8_tvalid,
    input [S_AXIS_SCALAR_8_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_8_tkeep,
    input [S_AXIS_SCALAR_8_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_8_tstrb,
    input [S_AXIS_SCALAR_8_DIRECT_DMWIDTH-1:0] s_axis_scalar_8_tdata,
    output s_axis_scalar_8_tready,
    //input AXI-Stream to Scalar interface 9
    input s_axis_scalar_9_aclk,
    input s_axis_scalar_9_aresetn,
    input s_axis_scalar_9_tlast,
    input s_axis_scalar_9_tvalid,
    input [S_AXIS_SCALAR_9_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_9_tkeep,
    input [S_AXIS_SCALAR_9_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_9_tstrb,
    input [S_AXIS_SCALAR_9_DIRECT_DMWIDTH-1:0] s_axis_scalar_9_tdata,
    output s_axis_scalar_9_tready,
    //input AXI-Stream to Scalar interface 10
    input s_axis_scalar_10_aclk,
    input s_axis_scalar_10_aresetn,
    input s_axis_scalar_10_tlast,
    input s_axis_scalar_10_tvalid,
    input [S_AXIS_SCALAR_10_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_10_tkeep,
    input [S_AXIS_SCALAR_10_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_10_tstrb,
    input [S_AXIS_SCALAR_10_DIRECT_DMWIDTH-1:0] s_axis_scalar_10_tdata,
    output s_axis_scalar_10_tready,
    //input AXI-Stream to Scalar interface 11
    input s_axis_scalar_11_aclk,
    input s_axis_scalar_11_aresetn,
    input s_axis_scalar_11_tlast,
    input s_axis_scalar_11_tvalid,
    input [S_AXIS_SCALAR_11_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_11_tkeep,
    input [S_AXIS_SCALAR_11_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_11_tstrb,
    input [S_AXIS_SCALAR_11_DIRECT_DMWIDTH-1:0] s_axis_scalar_11_tdata,
    output s_axis_scalar_11_tready,
    //input AXI-Stream to Scalar interface 12
    input s_axis_scalar_12_aclk,
    input s_axis_scalar_12_aresetn,
    input s_axis_scalar_12_tlast,
    input s_axis_scalar_12_tvalid,
    input [S_AXIS_SCALAR_12_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_12_tkeep,
    input [S_AXIS_SCALAR_12_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_12_tstrb,
    input [S_AXIS_SCALAR_12_DIRECT_DMWIDTH-1:0] s_axis_scalar_12_tdata,
    output s_axis_scalar_12_tready,
    //input AXI-Stream to Scalar interface 13
    input s_axis_scalar_13_aclk,
    input s_axis_scalar_13_aresetn,
    input s_axis_scalar_13_tlast,
    input s_axis_scalar_13_tvalid,
    input [S_AXIS_SCALAR_13_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_13_tkeep,
    input [S_AXIS_SCALAR_13_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_13_tstrb,
    input [S_AXIS_SCALAR_13_DIRECT_DMWIDTH-1:0] s_axis_scalar_13_tdata,
    output s_axis_scalar_13_tready,
    //input AXI-Stream to Scalar interface 14
    input s_axis_scalar_14_aclk,
    input s_axis_scalar_14_aresetn,
    input s_axis_scalar_14_tlast,
    input s_axis_scalar_14_tvalid,
    input [S_AXIS_SCALAR_14_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_14_tkeep,
    input [S_AXIS_SCALAR_14_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_14_tstrb,
    input [S_AXIS_SCALAR_14_DIRECT_DMWIDTH-1:0] s_axis_scalar_14_tdata,
    output s_axis_scalar_14_tready,
    //input AXI-Stream to Scalar interface 15
    input s_axis_scalar_15_aclk,
    input s_axis_scalar_15_aresetn,
    input s_axis_scalar_15_tlast,
    input s_axis_scalar_15_tvalid,
    input [S_AXIS_SCALAR_15_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_15_tkeep,
    input [S_AXIS_SCALAR_15_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_15_tstrb,
    input [S_AXIS_SCALAR_15_DIRECT_DMWIDTH-1:0] s_axis_scalar_15_tdata,
    output s_axis_scalar_15_tready,
    //input AXI-Stream to Scalar interface 16
    input s_axis_scalar_16_aclk,
    input s_axis_scalar_16_aresetn,
    input s_axis_scalar_16_tlast,
    input s_axis_scalar_16_tvalid,
    input [S_AXIS_SCALAR_16_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_16_tkeep,
    input [S_AXIS_SCALAR_16_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_16_tstrb,
    input [S_AXIS_SCALAR_16_DIRECT_DMWIDTH-1:0] s_axis_scalar_16_tdata,
    output s_axis_scalar_16_tready,
    //input AXI-Stream to Scalar interface 17
    input s_axis_scalar_17_aclk,
    input s_axis_scalar_17_aresetn,
    input s_axis_scalar_17_tlast,
    input s_axis_scalar_17_tvalid,
    input [S_AXIS_SCALAR_17_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_17_tkeep,
    input [S_AXIS_SCALAR_17_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_17_tstrb,
    input [S_AXIS_SCALAR_17_DIRECT_DMWIDTH-1:0] s_axis_scalar_17_tdata,
    output s_axis_scalar_17_tready,
    //input AXI-Stream to Scalar interface 18
    input s_axis_scalar_18_aclk,
    input s_axis_scalar_18_aresetn,
    input s_axis_scalar_18_tlast,
    input s_axis_scalar_18_tvalid,
    input [S_AXIS_SCALAR_18_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_18_tkeep,
    input [S_AXIS_SCALAR_18_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_18_tstrb,
    input [S_AXIS_SCALAR_18_DIRECT_DMWIDTH-1:0] s_axis_scalar_18_tdata,
    output s_axis_scalar_18_tready,
    //input AXI-Stream to Scalar interface 19
    input s_axis_scalar_19_aclk,
    input s_axis_scalar_19_aresetn,
    input s_axis_scalar_19_tlast,
    input s_axis_scalar_19_tvalid,
    input [S_AXIS_SCALAR_19_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_19_tkeep,
    input [S_AXIS_SCALAR_19_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_19_tstrb,
    input [S_AXIS_SCALAR_19_DIRECT_DMWIDTH-1:0] s_axis_scalar_19_tdata,
    output s_axis_scalar_19_tready,
    //input AXI-Stream to Scalar interface 20
    input s_axis_scalar_20_aclk,
    input s_axis_scalar_20_aresetn,
    input s_axis_scalar_20_tlast,
    input s_axis_scalar_20_tvalid,
    input [S_AXIS_SCALAR_20_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_20_tkeep,
    input [S_AXIS_SCALAR_20_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_20_tstrb,
    input [S_AXIS_SCALAR_20_DIRECT_DMWIDTH-1:0] s_axis_scalar_20_tdata,
    output s_axis_scalar_20_tready,
    //input AXI-Stream to Scalar interface 21
    input s_axis_scalar_21_aclk,
    input s_axis_scalar_21_aresetn,
    input s_axis_scalar_21_tlast,
    input s_axis_scalar_21_tvalid,
    input [S_AXIS_SCALAR_21_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_21_tkeep,
    input [S_AXIS_SCALAR_21_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_21_tstrb,
    input [S_AXIS_SCALAR_21_DIRECT_DMWIDTH-1:0] s_axis_scalar_21_tdata,
    output s_axis_scalar_21_tready,
    //input AXI-Stream to Scalar interface 22
    input s_axis_scalar_22_aclk,
    input s_axis_scalar_22_aresetn,
    input s_axis_scalar_22_tlast,
    input s_axis_scalar_22_tvalid,
    input [S_AXIS_SCALAR_22_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_22_tkeep,
    input [S_AXIS_SCALAR_22_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_22_tstrb,
    input [S_AXIS_SCALAR_22_DIRECT_DMWIDTH-1:0] s_axis_scalar_22_tdata,
    output s_axis_scalar_22_tready,
    //input AXI-Stream to Scalar interface 23
    input s_axis_scalar_23_aclk,
    input s_axis_scalar_23_aresetn,
    input s_axis_scalar_23_tlast,
    input s_axis_scalar_23_tvalid,
    input [S_AXIS_SCALAR_23_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_23_tkeep,
    input [S_AXIS_SCALAR_23_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_23_tstrb,
    input [S_AXIS_SCALAR_23_DIRECT_DMWIDTH-1:0] s_axis_scalar_23_tdata,
    output s_axis_scalar_23_tready,
    //input AXI-Stream to Scalar interface 24
    input s_axis_scalar_24_aclk,
    input s_axis_scalar_24_aresetn,
    input s_axis_scalar_24_tlast,
    input s_axis_scalar_24_tvalid,
    input [S_AXIS_SCALAR_24_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_24_tkeep,
    input [S_AXIS_SCALAR_24_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_24_tstrb,
    input [S_AXIS_SCALAR_24_DIRECT_DMWIDTH-1:0] s_axis_scalar_24_tdata,
    output s_axis_scalar_24_tready,
    //input AXI-Stream to Scalar interface 25
    input s_axis_scalar_25_aclk,
    input s_axis_scalar_25_aresetn,
    input s_axis_scalar_25_tlast,
    input s_axis_scalar_25_tvalid,
    input [S_AXIS_SCALAR_25_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_25_tkeep,
    input [S_AXIS_SCALAR_25_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_25_tstrb,
    input [S_AXIS_SCALAR_25_DIRECT_DMWIDTH-1:0] s_axis_scalar_25_tdata,
    output s_axis_scalar_25_tready,
    //input AXI-Stream to Scalar interface 26
    input s_axis_scalar_26_aclk,
    input s_axis_scalar_26_aresetn,
    input s_axis_scalar_26_tlast,
    input s_axis_scalar_26_tvalid,
    input [S_AXIS_SCALAR_26_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_26_tkeep,
    input [S_AXIS_SCALAR_26_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_26_tstrb,
    input [S_AXIS_SCALAR_26_DIRECT_DMWIDTH-1:0] s_axis_scalar_26_tdata,
    output s_axis_scalar_26_tready,
    //input AXI-Stream to Scalar interface 27
    input s_axis_scalar_27_aclk,
    input s_axis_scalar_27_aresetn,
    input s_axis_scalar_27_tlast,
    input s_axis_scalar_27_tvalid,
    input [S_AXIS_SCALAR_27_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_27_tkeep,
    input [S_AXIS_SCALAR_27_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_27_tstrb,
    input [S_AXIS_SCALAR_27_DIRECT_DMWIDTH-1:0] s_axis_scalar_27_tdata,
    output s_axis_scalar_27_tready,
    //input AXI-Stream to Scalar interface 28
    input s_axis_scalar_28_aclk,
    input s_axis_scalar_28_aresetn,
    input s_axis_scalar_28_tlast,
    input s_axis_scalar_28_tvalid,
    input [S_AXIS_SCALAR_28_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_28_tkeep,
    input [S_AXIS_SCALAR_28_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_28_tstrb,
    input [S_AXIS_SCALAR_28_DIRECT_DMWIDTH-1:0] s_axis_scalar_28_tdata,
    output s_axis_scalar_28_tready,
    //input AXI-Stream to Scalar interface 29
    input s_axis_scalar_29_aclk,
    input s_axis_scalar_29_aresetn,
    input s_axis_scalar_29_tlast,
    input s_axis_scalar_29_tvalid,
    input [S_AXIS_SCALAR_29_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_29_tkeep,
    input [S_AXIS_SCALAR_29_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_29_tstrb,
    input [S_AXIS_SCALAR_29_DIRECT_DMWIDTH-1:0] s_axis_scalar_29_tdata,
    output s_axis_scalar_29_tready,
    //input AXI-Stream to Scalar interface 30
    input s_axis_scalar_30_aclk,
    input s_axis_scalar_30_aresetn,
    input s_axis_scalar_30_tlast,
    input s_axis_scalar_30_tvalid,
    input [S_AXIS_SCALAR_30_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_30_tkeep,
    input [S_AXIS_SCALAR_30_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_30_tstrb,
    input [S_AXIS_SCALAR_30_DIRECT_DMWIDTH-1:0] s_axis_scalar_30_tdata,
    output s_axis_scalar_30_tready,
    //input AXI-Stream to Scalar interface 31
    input s_axis_scalar_31_aclk,
    input s_axis_scalar_31_aresetn,
    input s_axis_scalar_31_tlast,
    input s_axis_scalar_31_tvalid,
    input [S_AXIS_SCALAR_31_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_31_tkeep,
    input [S_AXIS_SCALAR_31_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_31_tstrb,
    input [S_AXIS_SCALAR_31_DIRECT_DMWIDTH-1:0] s_axis_scalar_31_tdata,
    output s_axis_scalar_31_tready,
    //input AXI-Stream to Scalar interface 32
    input s_axis_scalar_32_aclk,
    input s_axis_scalar_32_aresetn,
    input s_axis_scalar_32_tlast,
    input s_axis_scalar_32_tvalid,
    input [S_AXIS_SCALAR_32_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_32_tkeep,
    input [S_AXIS_SCALAR_32_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_32_tstrb,
    input [S_AXIS_SCALAR_32_DIRECT_DMWIDTH-1:0] s_axis_scalar_32_tdata,
    output s_axis_scalar_32_tready,
    //input AXI-Stream to Scalar interface 33
    input s_axis_scalar_33_aclk,
    input s_axis_scalar_33_aresetn,
    input s_axis_scalar_33_tlast,
    input s_axis_scalar_33_tvalid,
    input [S_AXIS_SCALAR_33_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_33_tkeep,
    input [S_AXIS_SCALAR_33_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_33_tstrb,
    input [S_AXIS_SCALAR_33_DIRECT_DMWIDTH-1:0] s_axis_scalar_33_tdata,
    output s_axis_scalar_33_tready,
    //input AXI-Stream to Scalar interface 34
    input s_axis_scalar_34_aclk,
    input s_axis_scalar_34_aresetn,
    input s_axis_scalar_34_tlast,
    input s_axis_scalar_34_tvalid,
    input [S_AXIS_SCALAR_34_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_34_tkeep,
    input [S_AXIS_SCALAR_34_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_34_tstrb,
    input [S_AXIS_SCALAR_34_DIRECT_DMWIDTH-1:0] s_axis_scalar_34_tdata,
    output s_axis_scalar_34_tready,
    //input AXI-Stream to Scalar interface 35
    input s_axis_scalar_35_aclk,
    input s_axis_scalar_35_aresetn,
    input s_axis_scalar_35_tlast,
    input s_axis_scalar_35_tvalid,
    input [S_AXIS_SCALAR_35_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_35_tkeep,
    input [S_AXIS_SCALAR_35_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_35_tstrb,
    input [S_AXIS_SCALAR_35_DIRECT_DMWIDTH-1:0] s_axis_scalar_35_tdata,
    output s_axis_scalar_35_tready,
    //input AXI-Stream to Scalar interface 36
    input s_axis_scalar_36_aclk,
    input s_axis_scalar_36_aresetn,
    input s_axis_scalar_36_tlast,
    input s_axis_scalar_36_tvalid,
    input [S_AXIS_SCALAR_36_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_36_tkeep,
    input [S_AXIS_SCALAR_36_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_36_tstrb,
    input [S_AXIS_SCALAR_36_DIRECT_DMWIDTH-1:0] s_axis_scalar_36_tdata,
    output s_axis_scalar_36_tready,
    //input AXI-Stream to Scalar interface 37
    input s_axis_scalar_37_aclk,
    input s_axis_scalar_37_aresetn,
    input s_axis_scalar_37_tlast,
    input s_axis_scalar_37_tvalid,
    input [S_AXIS_SCALAR_37_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_37_tkeep,
    input [S_AXIS_SCALAR_37_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_37_tstrb,
    input [S_AXIS_SCALAR_37_DIRECT_DMWIDTH-1:0] s_axis_scalar_37_tdata,
    output s_axis_scalar_37_tready,
    //input AXI-Stream to Scalar interface 38
    input s_axis_scalar_38_aclk,
    input s_axis_scalar_38_aresetn,
    input s_axis_scalar_38_tlast,
    input s_axis_scalar_38_tvalid,
    input [S_AXIS_SCALAR_38_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_38_tkeep,
    input [S_AXIS_SCALAR_38_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_38_tstrb,
    input [S_AXIS_SCALAR_38_DIRECT_DMWIDTH-1:0] s_axis_scalar_38_tdata,
    output s_axis_scalar_38_tready,
    //input AXI-Stream to Scalar interface 39
    input s_axis_scalar_39_aclk,
    input s_axis_scalar_39_aresetn,
    input s_axis_scalar_39_tlast,
    input s_axis_scalar_39_tvalid,
    input [S_AXIS_SCALAR_39_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_39_tkeep,
    input [S_AXIS_SCALAR_39_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_39_tstrb,
    input [S_AXIS_SCALAR_39_DIRECT_DMWIDTH-1:0] s_axis_scalar_39_tdata,
    output s_axis_scalar_39_tready,
    //input AXI-Stream to Scalar interface 40
    input s_axis_scalar_40_aclk,
    input s_axis_scalar_40_aresetn,
    input s_axis_scalar_40_tlast,
    input s_axis_scalar_40_tvalid,
    input [S_AXIS_SCALAR_40_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_40_tkeep,
    input [S_AXIS_SCALAR_40_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_40_tstrb,
    input [S_AXIS_SCALAR_40_DIRECT_DMWIDTH-1:0] s_axis_scalar_40_tdata,
    output s_axis_scalar_40_tready,
    //input AXI-Stream to Scalar interface 41
    input s_axis_scalar_41_aclk,
    input s_axis_scalar_41_aresetn,
    input s_axis_scalar_41_tlast,
    input s_axis_scalar_41_tvalid,
    input [S_AXIS_SCALAR_41_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_41_tkeep,
    input [S_AXIS_SCALAR_41_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_41_tstrb,
    input [S_AXIS_SCALAR_41_DIRECT_DMWIDTH-1:0] s_axis_scalar_41_tdata,
    output s_axis_scalar_41_tready,
    //input AXI-Stream to Scalar interface 42
    input s_axis_scalar_42_aclk,
    input s_axis_scalar_42_aresetn,
    input s_axis_scalar_42_tlast,
    input s_axis_scalar_42_tvalid,
    input [S_AXIS_SCALAR_42_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_42_tkeep,
    input [S_AXIS_SCALAR_42_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_42_tstrb,
    input [S_AXIS_SCALAR_42_DIRECT_DMWIDTH-1:0] s_axis_scalar_42_tdata,
    output s_axis_scalar_42_tready,
    //input AXI-Stream to Scalar interface 43
    input s_axis_scalar_43_aclk,
    input s_axis_scalar_43_aresetn,
    input s_axis_scalar_43_tlast,
    input s_axis_scalar_43_tvalid,
    input [S_AXIS_SCALAR_43_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_43_tkeep,
    input [S_AXIS_SCALAR_43_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_43_tstrb,
    input [S_AXIS_SCALAR_43_DIRECT_DMWIDTH-1:0] s_axis_scalar_43_tdata,
    output s_axis_scalar_43_tready,
    //input AXI-Stream to Scalar interface 44
    input s_axis_scalar_44_aclk,
    input s_axis_scalar_44_aresetn,
    input s_axis_scalar_44_tlast,
    input s_axis_scalar_44_tvalid,
    input [S_AXIS_SCALAR_44_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_44_tkeep,
    input [S_AXIS_SCALAR_44_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_44_tstrb,
    input [S_AXIS_SCALAR_44_DIRECT_DMWIDTH-1:0] s_axis_scalar_44_tdata,
    output s_axis_scalar_44_tready,
    //input AXI-Stream to Scalar interface 45
    input s_axis_scalar_45_aclk,
    input s_axis_scalar_45_aresetn,
    input s_axis_scalar_45_tlast,
    input s_axis_scalar_45_tvalid,
    input [S_AXIS_SCALAR_45_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_45_tkeep,
    input [S_AXIS_SCALAR_45_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_45_tstrb,
    input [S_AXIS_SCALAR_45_DIRECT_DMWIDTH-1:0] s_axis_scalar_45_tdata,
    output s_axis_scalar_45_tready,
    //input AXI-Stream to Scalar interface 46
    input s_axis_scalar_46_aclk,
    input s_axis_scalar_46_aresetn,
    input s_axis_scalar_46_tlast,
    input s_axis_scalar_46_tvalid,
    input [S_AXIS_SCALAR_46_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_46_tkeep,
    input [S_AXIS_SCALAR_46_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_46_tstrb,
    input [S_AXIS_SCALAR_46_DIRECT_DMWIDTH-1:0] s_axis_scalar_46_tdata,
    output s_axis_scalar_46_tready,
    //input AXI-Stream to Scalar interface 47
    input s_axis_scalar_47_aclk,
    input s_axis_scalar_47_aresetn,
    input s_axis_scalar_47_tlast,
    input s_axis_scalar_47_tvalid,
    input [S_AXIS_SCALAR_47_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_47_tkeep,
    input [S_AXIS_SCALAR_47_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_47_tstrb,
    input [S_AXIS_SCALAR_47_DIRECT_DMWIDTH-1:0] s_axis_scalar_47_tdata,
    output s_axis_scalar_47_tready,
    //input AXI-Stream to Scalar interface 48
    input s_axis_scalar_48_aclk,
    input s_axis_scalar_48_aresetn,
    input s_axis_scalar_48_tlast,
    input s_axis_scalar_48_tvalid,
    input [S_AXIS_SCALAR_48_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_48_tkeep,
    input [S_AXIS_SCALAR_48_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_48_tstrb,
    input [S_AXIS_SCALAR_48_DIRECT_DMWIDTH-1:0] s_axis_scalar_48_tdata,
    output s_axis_scalar_48_tready,
    //input AXI-Stream to Scalar interface 49
    input s_axis_scalar_49_aclk,
    input s_axis_scalar_49_aresetn,
    input s_axis_scalar_49_tlast,
    input s_axis_scalar_49_tvalid,
    input [S_AXIS_SCALAR_49_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_49_tkeep,
    input [S_AXIS_SCALAR_49_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_49_tstrb,
    input [S_AXIS_SCALAR_49_DIRECT_DMWIDTH-1:0] s_axis_scalar_49_tdata,
    output s_axis_scalar_49_tready,
    //input AXI-Stream to Scalar interface 50
    input s_axis_scalar_50_aclk,
    input s_axis_scalar_50_aresetn,
    input s_axis_scalar_50_tlast,
    input s_axis_scalar_50_tvalid,
    input [S_AXIS_SCALAR_50_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_50_tkeep,
    input [S_AXIS_SCALAR_50_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_50_tstrb,
    input [S_AXIS_SCALAR_50_DIRECT_DMWIDTH-1:0] s_axis_scalar_50_tdata,
    output s_axis_scalar_50_tready,
    //input AXI-Stream to Scalar interface 51
    input s_axis_scalar_51_aclk,
    input s_axis_scalar_51_aresetn,
    input s_axis_scalar_51_tlast,
    input s_axis_scalar_51_tvalid,
    input [S_AXIS_SCALAR_51_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_51_tkeep,
    input [S_AXIS_SCALAR_51_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_51_tstrb,
    input [S_AXIS_SCALAR_51_DIRECT_DMWIDTH-1:0] s_axis_scalar_51_tdata,
    output s_axis_scalar_51_tready,
    //input AXI-Stream to Scalar interface 52
    input s_axis_scalar_52_aclk,
    input s_axis_scalar_52_aresetn,
    input s_axis_scalar_52_tlast,
    input s_axis_scalar_52_tvalid,
    input [S_AXIS_SCALAR_52_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_52_tkeep,
    input [S_AXIS_SCALAR_52_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_52_tstrb,
    input [S_AXIS_SCALAR_52_DIRECT_DMWIDTH-1:0] s_axis_scalar_52_tdata,
    output s_axis_scalar_52_tready,
    //input AXI-Stream to Scalar interface 53
    input s_axis_scalar_53_aclk,
    input s_axis_scalar_53_aresetn,
    input s_axis_scalar_53_tlast,
    input s_axis_scalar_53_tvalid,
    input [S_AXIS_SCALAR_53_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_53_tkeep,
    input [S_AXIS_SCALAR_53_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_53_tstrb,
    input [S_AXIS_SCALAR_53_DIRECT_DMWIDTH-1:0] s_axis_scalar_53_tdata,
    output s_axis_scalar_53_tready,
    //input AXI-Stream to Scalar interface 54
    input s_axis_scalar_54_aclk,
    input s_axis_scalar_54_aresetn,
    input s_axis_scalar_54_tlast,
    input s_axis_scalar_54_tvalid,
    input [S_AXIS_SCALAR_54_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_54_tkeep,
    input [S_AXIS_SCALAR_54_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_54_tstrb,
    input [S_AXIS_SCALAR_54_DIRECT_DMWIDTH-1:0] s_axis_scalar_54_tdata,
    output s_axis_scalar_54_tready,
    //input AXI-Stream to Scalar interface 55
    input s_axis_scalar_55_aclk,
    input s_axis_scalar_55_aresetn,
    input s_axis_scalar_55_tlast,
    input s_axis_scalar_55_tvalid,
    input [S_AXIS_SCALAR_55_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_55_tkeep,
    input [S_AXIS_SCALAR_55_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_55_tstrb,
    input [S_AXIS_SCALAR_55_DIRECT_DMWIDTH-1:0] s_axis_scalar_55_tdata,
    output s_axis_scalar_55_tready,
    //input AXI-Stream to Scalar interface 56
    input s_axis_scalar_56_aclk,
    input s_axis_scalar_56_aresetn,
    input s_axis_scalar_56_tlast,
    input s_axis_scalar_56_tvalid,
    input [S_AXIS_SCALAR_56_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_56_tkeep,
    input [S_AXIS_SCALAR_56_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_56_tstrb,
    input [S_AXIS_SCALAR_56_DIRECT_DMWIDTH-1:0] s_axis_scalar_56_tdata,
    output s_axis_scalar_56_tready,
    //input AXI-Stream to Scalar interface 57
    input s_axis_scalar_57_aclk,
    input s_axis_scalar_57_aresetn,
    input s_axis_scalar_57_tlast,
    input s_axis_scalar_57_tvalid,
    input [S_AXIS_SCALAR_57_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_57_tkeep,
    input [S_AXIS_SCALAR_57_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_57_tstrb,
    input [S_AXIS_SCALAR_57_DIRECT_DMWIDTH-1:0] s_axis_scalar_57_tdata,
    output s_axis_scalar_57_tready,
    //input AXI-Stream to Scalar interface 58
    input s_axis_scalar_58_aclk,
    input s_axis_scalar_58_aresetn,
    input s_axis_scalar_58_tlast,
    input s_axis_scalar_58_tvalid,
    input [S_AXIS_SCALAR_58_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_58_tkeep,
    input [S_AXIS_SCALAR_58_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_58_tstrb,
    input [S_AXIS_SCALAR_58_DIRECT_DMWIDTH-1:0] s_axis_scalar_58_tdata,
    output s_axis_scalar_58_tready,
    //input AXI-Stream to Scalar interface 59
    input s_axis_scalar_59_aclk,
    input s_axis_scalar_59_aresetn,
    input s_axis_scalar_59_tlast,
    input s_axis_scalar_59_tvalid,
    input [S_AXIS_SCALAR_59_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_59_tkeep,
    input [S_AXIS_SCALAR_59_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_59_tstrb,
    input [S_AXIS_SCALAR_59_DIRECT_DMWIDTH-1:0] s_axis_scalar_59_tdata,
    output s_axis_scalar_59_tready,
    //input AXI-Stream to Scalar interface 60
    input s_axis_scalar_60_aclk,
    input s_axis_scalar_60_aresetn,
    input s_axis_scalar_60_tlast,
    input s_axis_scalar_60_tvalid,
    input [S_AXIS_SCALAR_60_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_60_tkeep,
    input [S_AXIS_SCALAR_60_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_60_tstrb,
    input [S_AXIS_SCALAR_60_DIRECT_DMWIDTH-1:0] s_axis_scalar_60_tdata,
    output s_axis_scalar_60_tready,
    //input AXI-Stream to Scalar interface 61
    input s_axis_scalar_61_aclk,
    input s_axis_scalar_61_aresetn,
    input s_axis_scalar_61_tlast,
    input s_axis_scalar_61_tvalid,
    input [S_AXIS_SCALAR_61_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_61_tkeep,
    input [S_AXIS_SCALAR_61_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_61_tstrb,
    input [S_AXIS_SCALAR_61_DIRECT_DMWIDTH-1:0] s_axis_scalar_61_tdata,
    output s_axis_scalar_61_tready,
    //input AXI-Stream to Scalar interface 62
    input s_axis_scalar_62_aclk,
    input s_axis_scalar_62_aresetn,
    input s_axis_scalar_62_tlast,
    input s_axis_scalar_62_tvalid,
    input [S_AXIS_SCALAR_62_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_62_tkeep,
    input [S_AXIS_SCALAR_62_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_62_tstrb,
    input [S_AXIS_SCALAR_62_DIRECT_DMWIDTH-1:0] s_axis_scalar_62_tdata,
    output s_axis_scalar_62_tready,
    //input AXI-Stream to Scalar interface 63
    input s_axis_scalar_63_aclk,
    input s_axis_scalar_63_aresetn,
    input s_axis_scalar_63_tlast,
    input s_axis_scalar_63_tvalid,
    input [S_AXIS_SCALAR_63_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_63_tkeep,
    input [S_AXIS_SCALAR_63_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_63_tstrb,
    input [S_AXIS_SCALAR_63_DIRECT_DMWIDTH-1:0] s_axis_scalar_63_tdata,
    output s_axis_scalar_63_tready,
    //input AXI-Stream to Scalar interface 64
    input s_axis_scalar_64_aclk,
    input s_axis_scalar_64_aresetn,
    input s_axis_scalar_64_tlast,
    input s_axis_scalar_64_tvalid,
    input [S_AXIS_SCALAR_64_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_64_tkeep,
    input [S_AXIS_SCALAR_64_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_64_tstrb,
    input [S_AXIS_SCALAR_64_DIRECT_DMWIDTH-1:0] s_axis_scalar_64_tdata,
    output s_axis_scalar_64_tready,
    //input AXI-Stream to Scalar interface 65
    input s_axis_scalar_65_aclk,
    input s_axis_scalar_65_aresetn,
    input s_axis_scalar_65_tlast,
    input s_axis_scalar_65_tvalid,
    input [S_AXIS_SCALAR_65_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_65_tkeep,
    input [S_AXIS_SCALAR_65_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_65_tstrb,
    input [S_AXIS_SCALAR_65_DIRECT_DMWIDTH-1:0] s_axis_scalar_65_tdata,
    output s_axis_scalar_65_tready,
    //input AXI-Stream to Scalar interface 66
    input s_axis_scalar_66_aclk,
    input s_axis_scalar_66_aresetn,
    input s_axis_scalar_66_tlast,
    input s_axis_scalar_66_tvalid,
    input [S_AXIS_SCALAR_66_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_66_tkeep,
    input [S_AXIS_SCALAR_66_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_66_tstrb,
    input [S_AXIS_SCALAR_66_DIRECT_DMWIDTH-1:0] s_axis_scalar_66_tdata,
    output s_axis_scalar_66_tready,
    //input AXI-Stream to Scalar interface 67
    input s_axis_scalar_67_aclk,
    input s_axis_scalar_67_aresetn,
    input s_axis_scalar_67_tlast,
    input s_axis_scalar_67_tvalid,
    input [S_AXIS_SCALAR_67_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_67_tkeep,
    input [S_AXIS_SCALAR_67_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_67_tstrb,
    input [S_AXIS_SCALAR_67_DIRECT_DMWIDTH-1:0] s_axis_scalar_67_tdata,
    output s_axis_scalar_67_tready,
    //input AXI-Stream to Scalar interface 68
    input s_axis_scalar_68_aclk,
    input s_axis_scalar_68_aresetn,
    input s_axis_scalar_68_tlast,
    input s_axis_scalar_68_tvalid,
    input [S_AXIS_SCALAR_68_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_68_tkeep,
    input [S_AXIS_SCALAR_68_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_68_tstrb,
    input [S_AXIS_SCALAR_68_DIRECT_DMWIDTH-1:0] s_axis_scalar_68_tdata,
    output s_axis_scalar_68_tready,
    //input AXI-Stream to Scalar interface 69
    input s_axis_scalar_69_aclk,
    input s_axis_scalar_69_aresetn,
    input s_axis_scalar_69_tlast,
    input s_axis_scalar_69_tvalid,
    input [S_AXIS_SCALAR_69_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_69_tkeep,
    input [S_AXIS_SCALAR_69_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_69_tstrb,
    input [S_AXIS_SCALAR_69_DIRECT_DMWIDTH-1:0] s_axis_scalar_69_tdata,
    output s_axis_scalar_69_tready,
    //input AXI-Stream to Scalar interface 70
    input s_axis_scalar_70_aclk,
    input s_axis_scalar_70_aresetn,
    input s_axis_scalar_70_tlast,
    input s_axis_scalar_70_tvalid,
    input [S_AXIS_SCALAR_70_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_70_tkeep,
    input [S_AXIS_SCALAR_70_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_70_tstrb,
    input [S_AXIS_SCALAR_70_DIRECT_DMWIDTH-1:0] s_axis_scalar_70_tdata,
    output s_axis_scalar_70_tready,
    //input AXI-Stream to Scalar interface 71
    input s_axis_scalar_71_aclk,
    input s_axis_scalar_71_aresetn,
    input s_axis_scalar_71_tlast,
    input s_axis_scalar_71_tvalid,
    input [S_AXIS_SCALAR_71_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_71_tkeep,
    input [S_AXIS_SCALAR_71_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_71_tstrb,
    input [S_AXIS_SCALAR_71_DIRECT_DMWIDTH-1:0] s_axis_scalar_71_tdata,
    output s_axis_scalar_71_tready,
    //input AXI-Stream to Scalar interface 72
    input s_axis_scalar_72_aclk,
    input s_axis_scalar_72_aresetn,
    input s_axis_scalar_72_tlast,
    input s_axis_scalar_72_tvalid,
    input [S_AXIS_SCALAR_72_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_72_tkeep,
    input [S_AXIS_SCALAR_72_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_72_tstrb,
    input [S_AXIS_SCALAR_72_DIRECT_DMWIDTH-1:0] s_axis_scalar_72_tdata,
    output s_axis_scalar_72_tready,
    //input AXI-Stream to Scalar interface 73
    input s_axis_scalar_73_aclk,
    input s_axis_scalar_73_aresetn,
    input s_axis_scalar_73_tlast,
    input s_axis_scalar_73_tvalid,
    input [S_AXIS_SCALAR_73_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_73_tkeep,
    input [S_AXIS_SCALAR_73_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_73_tstrb,
    input [S_AXIS_SCALAR_73_DIRECT_DMWIDTH-1:0] s_axis_scalar_73_tdata,
    output s_axis_scalar_73_tready,
    //input AXI-Stream to Scalar interface 74
    input s_axis_scalar_74_aclk,
    input s_axis_scalar_74_aresetn,
    input s_axis_scalar_74_tlast,
    input s_axis_scalar_74_tvalid,
    input [S_AXIS_SCALAR_74_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_74_tkeep,
    input [S_AXIS_SCALAR_74_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_74_tstrb,
    input [S_AXIS_SCALAR_74_DIRECT_DMWIDTH-1:0] s_axis_scalar_74_tdata,
    output s_axis_scalar_74_tready,
    //input AXI-Stream to Scalar interface 75
    input s_axis_scalar_75_aclk,
    input s_axis_scalar_75_aresetn,
    input s_axis_scalar_75_tlast,
    input s_axis_scalar_75_tvalid,
    input [S_AXIS_SCALAR_75_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_75_tkeep,
    input [S_AXIS_SCALAR_75_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_75_tstrb,
    input [S_AXIS_SCALAR_75_DIRECT_DMWIDTH-1:0] s_axis_scalar_75_tdata,
    output s_axis_scalar_75_tready,
    //input AXI-Stream to Scalar interface 76
    input s_axis_scalar_76_aclk,
    input s_axis_scalar_76_aresetn,
    input s_axis_scalar_76_tlast,
    input s_axis_scalar_76_tvalid,
    input [S_AXIS_SCALAR_76_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_76_tkeep,
    input [S_AXIS_SCALAR_76_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_76_tstrb,
    input [S_AXIS_SCALAR_76_DIRECT_DMWIDTH-1:0] s_axis_scalar_76_tdata,
    output s_axis_scalar_76_tready,
    //input AXI-Stream to Scalar interface 77
    input s_axis_scalar_77_aclk,
    input s_axis_scalar_77_aresetn,
    input s_axis_scalar_77_tlast,
    input s_axis_scalar_77_tvalid,
    input [S_AXIS_SCALAR_77_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_77_tkeep,
    input [S_AXIS_SCALAR_77_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_77_tstrb,
    input [S_AXIS_SCALAR_77_DIRECT_DMWIDTH-1:0] s_axis_scalar_77_tdata,
    output s_axis_scalar_77_tready,
    //input AXI-Stream to Scalar interface 78
    input s_axis_scalar_78_aclk,
    input s_axis_scalar_78_aresetn,
    input s_axis_scalar_78_tlast,
    input s_axis_scalar_78_tvalid,
    input [S_AXIS_SCALAR_78_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_78_tkeep,
    input [S_AXIS_SCALAR_78_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_78_tstrb,
    input [S_AXIS_SCALAR_78_DIRECT_DMWIDTH-1:0] s_axis_scalar_78_tdata,
    output s_axis_scalar_78_tready,
    //input AXI-Stream to Scalar interface 79
    input s_axis_scalar_79_aclk,
    input s_axis_scalar_79_aresetn,
    input s_axis_scalar_79_tlast,
    input s_axis_scalar_79_tvalid,
    input [S_AXIS_SCALAR_79_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_79_tkeep,
    input [S_AXIS_SCALAR_79_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_79_tstrb,
    input [S_AXIS_SCALAR_79_DIRECT_DMWIDTH-1:0] s_axis_scalar_79_tdata,
    output s_axis_scalar_79_tready,
    //input AXI-Stream to Scalar interface 80
    input s_axis_scalar_80_aclk,
    input s_axis_scalar_80_aresetn,
    input s_axis_scalar_80_tlast,
    input s_axis_scalar_80_tvalid,
    input [S_AXIS_SCALAR_80_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_80_tkeep,
    input [S_AXIS_SCALAR_80_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_80_tstrb,
    input [S_AXIS_SCALAR_80_DIRECT_DMWIDTH-1:0] s_axis_scalar_80_tdata,
    output s_axis_scalar_80_tready,
    //input AXI-Stream to Scalar interface 81
    input s_axis_scalar_81_aclk,
    input s_axis_scalar_81_aresetn,
    input s_axis_scalar_81_tlast,
    input s_axis_scalar_81_tvalid,
    input [S_AXIS_SCALAR_81_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_81_tkeep,
    input [S_AXIS_SCALAR_81_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_81_tstrb,
    input [S_AXIS_SCALAR_81_DIRECT_DMWIDTH-1:0] s_axis_scalar_81_tdata,
    output s_axis_scalar_81_tready,
    //input AXI-Stream to Scalar interface 82
    input s_axis_scalar_82_aclk,
    input s_axis_scalar_82_aresetn,
    input s_axis_scalar_82_tlast,
    input s_axis_scalar_82_tvalid,
    input [S_AXIS_SCALAR_82_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_82_tkeep,
    input [S_AXIS_SCALAR_82_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_82_tstrb,
    input [S_AXIS_SCALAR_82_DIRECT_DMWIDTH-1:0] s_axis_scalar_82_tdata,
    output s_axis_scalar_82_tready,
    //input AXI-Stream to Scalar interface 83
    input s_axis_scalar_83_aclk,
    input s_axis_scalar_83_aresetn,
    input s_axis_scalar_83_tlast,
    input s_axis_scalar_83_tvalid,
    input [S_AXIS_SCALAR_83_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_83_tkeep,
    input [S_AXIS_SCALAR_83_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_83_tstrb,
    input [S_AXIS_SCALAR_83_DIRECT_DMWIDTH-1:0] s_axis_scalar_83_tdata,
    output s_axis_scalar_83_tready,
    //input AXI-Stream to Scalar interface 84
    input s_axis_scalar_84_aclk,
    input s_axis_scalar_84_aresetn,
    input s_axis_scalar_84_tlast,
    input s_axis_scalar_84_tvalid,
    input [S_AXIS_SCALAR_84_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_84_tkeep,
    input [S_AXIS_SCALAR_84_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_84_tstrb,
    input [S_AXIS_SCALAR_84_DIRECT_DMWIDTH-1:0] s_axis_scalar_84_tdata,
    output s_axis_scalar_84_tready,
    //input AXI-Stream to Scalar interface 85
    input s_axis_scalar_85_aclk,
    input s_axis_scalar_85_aresetn,
    input s_axis_scalar_85_tlast,
    input s_axis_scalar_85_tvalid,
    input [S_AXIS_SCALAR_85_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_85_tkeep,
    input [S_AXIS_SCALAR_85_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_85_tstrb,
    input [S_AXIS_SCALAR_85_DIRECT_DMWIDTH-1:0] s_axis_scalar_85_tdata,
    output s_axis_scalar_85_tready,
    //input AXI-Stream to Scalar interface 86
    input s_axis_scalar_86_aclk,
    input s_axis_scalar_86_aresetn,
    input s_axis_scalar_86_tlast,
    input s_axis_scalar_86_tvalid,
    input [S_AXIS_SCALAR_86_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_86_tkeep,
    input [S_AXIS_SCALAR_86_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_86_tstrb,
    input [S_AXIS_SCALAR_86_DIRECT_DMWIDTH-1:0] s_axis_scalar_86_tdata,
    output s_axis_scalar_86_tready,
    //input AXI-Stream to Scalar interface 87
    input s_axis_scalar_87_aclk,
    input s_axis_scalar_87_aresetn,
    input s_axis_scalar_87_tlast,
    input s_axis_scalar_87_tvalid,
    input [S_AXIS_SCALAR_87_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_87_tkeep,
    input [S_AXIS_SCALAR_87_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_87_tstrb,
    input [S_AXIS_SCALAR_87_DIRECT_DMWIDTH-1:0] s_axis_scalar_87_tdata,
    output s_axis_scalar_87_tready,
    //input AXI-Stream to Scalar interface 88
    input s_axis_scalar_88_aclk,
    input s_axis_scalar_88_aresetn,
    input s_axis_scalar_88_tlast,
    input s_axis_scalar_88_tvalid,
    input [S_AXIS_SCALAR_88_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_88_tkeep,
    input [S_AXIS_SCALAR_88_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_88_tstrb,
    input [S_AXIS_SCALAR_88_DIRECT_DMWIDTH-1:0] s_axis_scalar_88_tdata,
    output s_axis_scalar_88_tready,
    //input AXI-Stream to Scalar interface 89
    input s_axis_scalar_89_aclk,
    input s_axis_scalar_89_aresetn,
    input s_axis_scalar_89_tlast,
    input s_axis_scalar_89_tvalid,
    input [S_AXIS_SCALAR_89_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_89_tkeep,
    input [S_AXIS_SCALAR_89_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_89_tstrb,
    input [S_AXIS_SCALAR_89_DIRECT_DMWIDTH-1:0] s_axis_scalar_89_tdata,
    output s_axis_scalar_89_tready,
    //input AXI-Stream to Scalar interface 90
    input s_axis_scalar_90_aclk,
    input s_axis_scalar_90_aresetn,
    input s_axis_scalar_90_tlast,
    input s_axis_scalar_90_tvalid,
    input [S_AXIS_SCALAR_90_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_90_tkeep,
    input [S_AXIS_SCALAR_90_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_90_tstrb,
    input [S_AXIS_SCALAR_90_DIRECT_DMWIDTH-1:0] s_axis_scalar_90_tdata,
    output s_axis_scalar_90_tready,
    //input AXI-Stream to Scalar interface 91
    input s_axis_scalar_91_aclk,
    input s_axis_scalar_91_aresetn,
    input s_axis_scalar_91_tlast,
    input s_axis_scalar_91_tvalid,
    input [S_AXIS_SCALAR_91_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_91_tkeep,
    input [S_AXIS_SCALAR_91_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_91_tstrb,
    input [S_AXIS_SCALAR_91_DIRECT_DMWIDTH-1:0] s_axis_scalar_91_tdata,
    output s_axis_scalar_91_tready,
    //input AXI-Stream to Scalar interface 92
    input s_axis_scalar_92_aclk,
    input s_axis_scalar_92_aresetn,
    input s_axis_scalar_92_tlast,
    input s_axis_scalar_92_tvalid,
    input [S_AXIS_SCALAR_92_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_92_tkeep,
    input [S_AXIS_SCALAR_92_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_92_tstrb,
    input [S_AXIS_SCALAR_92_DIRECT_DMWIDTH-1:0] s_axis_scalar_92_tdata,
    output s_axis_scalar_92_tready,
    //input AXI-Stream to Scalar interface 93
    input s_axis_scalar_93_aclk,
    input s_axis_scalar_93_aresetn,
    input s_axis_scalar_93_tlast,
    input s_axis_scalar_93_tvalid,
    input [S_AXIS_SCALAR_93_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_93_tkeep,
    input [S_AXIS_SCALAR_93_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_93_tstrb,
    input [S_AXIS_SCALAR_93_DIRECT_DMWIDTH-1:0] s_axis_scalar_93_tdata,
    output s_axis_scalar_93_tready,
    //input AXI-Stream to Scalar interface 94
    input s_axis_scalar_94_aclk,
    input s_axis_scalar_94_aresetn,
    input s_axis_scalar_94_tlast,
    input s_axis_scalar_94_tvalid,
    input [S_AXIS_SCALAR_94_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_94_tkeep,
    input [S_AXIS_SCALAR_94_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_94_tstrb,
    input [S_AXIS_SCALAR_94_DIRECT_DMWIDTH-1:0] s_axis_scalar_94_tdata,
    output s_axis_scalar_94_tready,
    //input AXI-Stream to Scalar interface 95
    input s_axis_scalar_95_aclk,
    input s_axis_scalar_95_aresetn,
    input s_axis_scalar_95_tlast,
    input s_axis_scalar_95_tvalid,
    input [S_AXIS_SCALAR_95_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_95_tkeep,
    input [S_AXIS_SCALAR_95_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_95_tstrb,
    input [S_AXIS_SCALAR_95_DIRECT_DMWIDTH-1:0] s_axis_scalar_95_tdata,
    output s_axis_scalar_95_tready,
    //input AXI-Stream to Scalar interface 96
    input s_axis_scalar_96_aclk,
    input s_axis_scalar_96_aresetn,
    input s_axis_scalar_96_tlast,
    input s_axis_scalar_96_tvalid,
    input [S_AXIS_SCALAR_96_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_96_tkeep,
    input [S_AXIS_SCALAR_96_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_96_tstrb,
    input [S_AXIS_SCALAR_96_DIRECT_DMWIDTH-1:0] s_axis_scalar_96_tdata,
    output s_axis_scalar_96_tready,
    //input AXI-Stream to Scalar interface 97
    input s_axis_scalar_97_aclk,
    input s_axis_scalar_97_aresetn,
    input s_axis_scalar_97_tlast,
    input s_axis_scalar_97_tvalid,
    input [S_AXIS_SCALAR_97_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_97_tkeep,
    input [S_AXIS_SCALAR_97_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_97_tstrb,
    input [S_AXIS_SCALAR_97_DIRECT_DMWIDTH-1:0] s_axis_scalar_97_tdata,
    output s_axis_scalar_97_tready,
    //input AXI-Stream to Scalar interface 98
    input s_axis_scalar_98_aclk,
    input s_axis_scalar_98_aresetn,
    input s_axis_scalar_98_tlast,
    input s_axis_scalar_98_tvalid,
    input [S_AXIS_SCALAR_98_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_98_tkeep,
    input [S_AXIS_SCALAR_98_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_98_tstrb,
    input [S_AXIS_SCALAR_98_DIRECT_DMWIDTH-1:0] s_axis_scalar_98_tdata,
    output s_axis_scalar_98_tready,
    //input AXI-Stream to Scalar interface 99
    input s_axis_scalar_99_aclk,
    input s_axis_scalar_99_aresetn,
    input s_axis_scalar_99_tlast,
    input s_axis_scalar_99_tvalid,
    input [S_AXIS_SCALAR_99_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_99_tkeep,
    input [S_AXIS_SCALAR_99_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_99_tstrb,
    input [S_AXIS_SCALAR_99_DIRECT_DMWIDTH-1:0] s_axis_scalar_99_tdata,
    output s_axis_scalar_99_tready,
    //input AXI-Stream to Scalar interface 100
    input s_axis_scalar_100_aclk,
    input s_axis_scalar_100_aresetn,
    input s_axis_scalar_100_tlast,
    input s_axis_scalar_100_tvalid,
    input [S_AXIS_SCALAR_100_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_100_tkeep,
    input [S_AXIS_SCALAR_100_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_100_tstrb,
    input [S_AXIS_SCALAR_100_DIRECT_DMWIDTH-1:0] s_axis_scalar_100_tdata,
    output s_axis_scalar_100_tready,
    //input AXI-Stream to Scalar interface 101
    input s_axis_scalar_101_aclk,
    input s_axis_scalar_101_aresetn,
    input s_axis_scalar_101_tlast,
    input s_axis_scalar_101_tvalid,
    input [S_AXIS_SCALAR_101_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_101_tkeep,
    input [S_AXIS_SCALAR_101_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_101_tstrb,
    input [S_AXIS_SCALAR_101_DIRECT_DMWIDTH-1:0] s_axis_scalar_101_tdata,
    output s_axis_scalar_101_tready,
    //input AXI-Stream to Scalar interface 102
    input s_axis_scalar_102_aclk,
    input s_axis_scalar_102_aresetn,
    input s_axis_scalar_102_tlast,
    input s_axis_scalar_102_tvalid,
    input [S_AXIS_SCALAR_102_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_102_tkeep,
    input [S_AXIS_SCALAR_102_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_102_tstrb,
    input [S_AXIS_SCALAR_102_DIRECT_DMWIDTH-1:0] s_axis_scalar_102_tdata,
    output s_axis_scalar_102_tready,
    //input AXI-Stream to Scalar interface 103
    input s_axis_scalar_103_aclk,
    input s_axis_scalar_103_aresetn,
    input s_axis_scalar_103_tlast,
    input s_axis_scalar_103_tvalid,
    input [S_AXIS_SCALAR_103_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_103_tkeep,
    input [S_AXIS_SCALAR_103_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_103_tstrb,
    input [S_AXIS_SCALAR_103_DIRECT_DMWIDTH-1:0] s_axis_scalar_103_tdata,
    output s_axis_scalar_103_tready,
    //input AXI-Stream to Scalar interface 104
    input s_axis_scalar_104_aclk,
    input s_axis_scalar_104_aresetn,
    input s_axis_scalar_104_tlast,
    input s_axis_scalar_104_tvalid,
    input [S_AXIS_SCALAR_104_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_104_tkeep,
    input [S_AXIS_SCALAR_104_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_104_tstrb,
    input [S_AXIS_SCALAR_104_DIRECT_DMWIDTH-1:0] s_axis_scalar_104_tdata,
    output s_axis_scalar_104_tready,
    //input AXI-Stream to Scalar interface 105
    input s_axis_scalar_105_aclk,
    input s_axis_scalar_105_aresetn,
    input s_axis_scalar_105_tlast,
    input s_axis_scalar_105_tvalid,
    input [S_AXIS_SCALAR_105_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_105_tkeep,
    input [S_AXIS_SCALAR_105_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_105_tstrb,
    input [S_AXIS_SCALAR_105_DIRECT_DMWIDTH-1:0] s_axis_scalar_105_tdata,
    output s_axis_scalar_105_tready,
    //input AXI-Stream to Scalar interface 106
    input s_axis_scalar_106_aclk,
    input s_axis_scalar_106_aresetn,
    input s_axis_scalar_106_tlast,
    input s_axis_scalar_106_tvalid,
    input [S_AXIS_SCALAR_106_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_106_tkeep,
    input [S_AXIS_SCALAR_106_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_106_tstrb,
    input [S_AXIS_SCALAR_106_DIRECT_DMWIDTH-1:0] s_axis_scalar_106_tdata,
    output s_axis_scalar_106_tready,
    //input AXI-Stream to Scalar interface 107
    input s_axis_scalar_107_aclk,
    input s_axis_scalar_107_aresetn,
    input s_axis_scalar_107_tlast,
    input s_axis_scalar_107_tvalid,
    input [S_AXIS_SCALAR_107_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_107_tkeep,
    input [S_AXIS_SCALAR_107_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_107_tstrb,
    input [S_AXIS_SCALAR_107_DIRECT_DMWIDTH-1:0] s_axis_scalar_107_tdata,
    output s_axis_scalar_107_tready,
    //input AXI-Stream to Scalar interface 108
    input s_axis_scalar_108_aclk,
    input s_axis_scalar_108_aresetn,
    input s_axis_scalar_108_tlast,
    input s_axis_scalar_108_tvalid,
    input [S_AXIS_SCALAR_108_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_108_tkeep,
    input [S_AXIS_SCALAR_108_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_108_tstrb,
    input [S_AXIS_SCALAR_108_DIRECT_DMWIDTH-1:0] s_axis_scalar_108_tdata,
    output s_axis_scalar_108_tready,
    //input AXI-Stream to Scalar interface 109
    input s_axis_scalar_109_aclk,
    input s_axis_scalar_109_aresetn,
    input s_axis_scalar_109_tlast,
    input s_axis_scalar_109_tvalid,
    input [S_AXIS_SCALAR_109_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_109_tkeep,
    input [S_AXIS_SCALAR_109_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_109_tstrb,
    input [S_AXIS_SCALAR_109_DIRECT_DMWIDTH-1:0] s_axis_scalar_109_tdata,
    output s_axis_scalar_109_tready,
    //input AXI-Stream to Scalar interface 110
    input s_axis_scalar_110_aclk,
    input s_axis_scalar_110_aresetn,
    input s_axis_scalar_110_tlast,
    input s_axis_scalar_110_tvalid,
    input [S_AXIS_SCALAR_110_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_110_tkeep,
    input [S_AXIS_SCALAR_110_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_110_tstrb,
    input [S_AXIS_SCALAR_110_DIRECT_DMWIDTH-1:0] s_axis_scalar_110_tdata,
    output s_axis_scalar_110_tready,
    //input AXI-Stream to Scalar interface 111
    input s_axis_scalar_111_aclk,
    input s_axis_scalar_111_aresetn,
    input s_axis_scalar_111_tlast,
    input s_axis_scalar_111_tvalid,
    input [S_AXIS_SCALAR_111_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_111_tkeep,
    input [S_AXIS_SCALAR_111_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_111_tstrb,
    input [S_AXIS_SCALAR_111_DIRECT_DMWIDTH-1:0] s_axis_scalar_111_tdata,
    output s_axis_scalar_111_tready,
    //input AXI-Stream to Scalar interface 112
    input s_axis_scalar_112_aclk,
    input s_axis_scalar_112_aresetn,
    input s_axis_scalar_112_tlast,
    input s_axis_scalar_112_tvalid,
    input [S_AXIS_SCALAR_112_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_112_tkeep,
    input [S_AXIS_SCALAR_112_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_112_tstrb,
    input [S_AXIS_SCALAR_112_DIRECT_DMWIDTH-1:0] s_axis_scalar_112_tdata,
    output s_axis_scalar_112_tready,
    //input AXI-Stream to Scalar interface 113
    input s_axis_scalar_113_aclk,
    input s_axis_scalar_113_aresetn,
    input s_axis_scalar_113_tlast,
    input s_axis_scalar_113_tvalid,
    input [S_AXIS_SCALAR_113_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_113_tkeep,
    input [S_AXIS_SCALAR_113_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_113_tstrb,
    input [S_AXIS_SCALAR_113_DIRECT_DMWIDTH-1:0] s_axis_scalar_113_tdata,
    output s_axis_scalar_113_tready,
    //input AXI-Stream to Scalar interface 114
    input s_axis_scalar_114_aclk,
    input s_axis_scalar_114_aresetn,
    input s_axis_scalar_114_tlast,
    input s_axis_scalar_114_tvalid,
    input [S_AXIS_SCALAR_114_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_114_tkeep,
    input [S_AXIS_SCALAR_114_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_114_tstrb,
    input [S_AXIS_SCALAR_114_DIRECT_DMWIDTH-1:0] s_axis_scalar_114_tdata,
    output s_axis_scalar_114_tready,
    //input AXI-Stream to Scalar interface 115
    input s_axis_scalar_115_aclk,
    input s_axis_scalar_115_aresetn,
    input s_axis_scalar_115_tlast,
    input s_axis_scalar_115_tvalid,
    input [S_AXIS_SCALAR_115_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_115_tkeep,
    input [S_AXIS_SCALAR_115_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_115_tstrb,
    input [S_AXIS_SCALAR_115_DIRECT_DMWIDTH-1:0] s_axis_scalar_115_tdata,
    output s_axis_scalar_115_tready,
    //input AXI-Stream to Scalar interface 116
    input s_axis_scalar_116_aclk,
    input s_axis_scalar_116_aresetn,
    input s_axis_scalar_116_tlast,
    input s_axis_scalar_116_tvalid,
    input [S_AXIS_SCALAR_116_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_116_tkeep,
    input [S_AXIS_SCALAR_116_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_116_tstrb,
    input [S_AXIS_SCALAR_116_DIRECT_DMWIDTH-1:0] s_axis_scalar_116_tdata,
    output s_axis_scalar_116_tready,
    //input AXI-Stream to Scalar interface 117
    input s_axis_scalar_117_aclk,
    input s_axis_scalar_117_aresetn,
    input s_axis_scalar_117_tlast,
    input s_axis_scalar_117_tvalid,
    input [S_AXIS_SCALAR_117_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_117_tkeep,
    input [S_AXIS_SCALAR_117_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_117_tstrb,
    input [S_AXIS_SCALAR_117_DIRECT_DMWIDTH-1:0] s_axis_scalar_117_tdata,
    output s_axis_scalar_117_tready,
    //input AXI-Stream to Scalar interface 118
    input s_axis_scalar_118_aclk,
    input s_axis_scalar_118_aresetn,
    input s_axis_scalar_118_tlast,
    input s_axis_scalar_118_tvalid,
    input [S_AXIS_SCALAR_118_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_118_tkeep,
    input [S_AXIS_SCALAR_118_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_118_tstrb,
    input [S_AXIS_SCALAR_118_DIRECT_DMWIDTH-1:0] s_axis_scalar_118_tdata,
    output s_axis_scalar_118_tready,
    //input AXI-Stream to Scalar interface 119
    input s_axis_scalar_119_aclk,
    input s_axis_scalar_119_aresetn,
    input s_axis_scalar_119_tlast,
    input s_axis_scalar_119_tvalid,
    input [S_AXIS_SCALAR_119_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_119_tkeep,
    input [S_AXIS_SCALAR_119_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_119_tstrb,
    input [S_AXIS_SCALAR_119_DIRECT_DMWIDTH-1:0] s_axis_scalar_119_tdata,
    output s_axis_scalar_119_tready,
    //input AXI-Stream to Scalar interface 120
    input s_axis_scalar_120_aclk,
    input s_axis_scalar_120_aresetn,
    input s_axis_scalar_120_tlast,
    input s_axis_scalar_120_tvalid,
    input [S_AXIS_SCALAR_120_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_120_tkeep,
    input [S_AXIS_SCALAR_120_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_120_tstrb,
    input [S_AXIS_SCALAR_120_DIRECT_DMWIDTH-1:0] s_axis_scalar_120_tdata,
    output s_axis_scalar_120_tready,
    //input AXI-Stream to Scalar interface 121
    input s_axis_scalar_121_aclk,
    input s_axis_scalar_121_aresetn,
    input s_axis_scalar_121_tlast,
    input s_axis_scalar_121_tvalid,
    input [S_AXIS_SCALAR_121_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_121_tkeep,
    input [S_AXIS_SCALAR_121_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_121_tstrb,
    input [S_AXIS_SCALAR_121_DIRECT_DMWIDTH-1:0] s_axis_scalar_121_tdata,
    output s_axis_scalar_121_tready,
    //input AXI-Stream to Scalar interface 122
    input s_axis_scalar_122_aclk,
    input s_axis_scalar_122_aresetn,
    input s_axis_scalar_122_tlast,
    input s_axis_scalar_122_tvalid,
    input [S_AXIS_SCALAR_122_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_122_tkeep,
    input [S_AXIS_SCALAR_122_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_122_tstrb,
    input [S_AXIS_SCALAR_122_DIRECT_DMWIDTH-1:0] s_axis_scalar_122_tdata,
    output s_axis_scalar_122_tready,
    //input AXI-Stream to Scalar interface 123
    input s_axis_scalar_123_aclk,
    input s_axis_scalar_123_aresetn,
    input s_axis_scalar_123_tlast,
    input s_axis_scalar_123_tvalid,
    input [S_AXIS_SCALAR_123_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_123_tkeep,
    input [S_AXIS_SCALAR_123_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_123_tstrb,
    input [S_AXIS_SCALAR_123_DIRECT_DMWIDTH-1:0] s_axis_scalar_123_tdata,
    output s_axis_scalar_123_tready,
    //input AXI-Stream to Scalar interface 124
    input s_axis_scalar_124_aclk,
    input s_axis_scalar_124_aresetn,
    input s_axis_scalar_124_tlast,
    input s_axis_scalar_124_tvalid,
    input [S_AXIS_SCALAR_124_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_124_tkeep,
    input [S_AXIS_SCALAR_124_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_124_tstrb,
    input [S_AXIS_SCALAR_124_DIRECT_DMWIDTH-1:0] s_axis_scalar_124_tdata,
    output s_axis_scalar_124_tready,
    //input AXI-Stream to Scalar interface 125
    input s_axis_scalar_125_aclk,
    input s_axis_scalar_125_aresetn,
    input s_axis_scalar_125_tlast,
    input s_axis_scalar_125_tvalid,
    input [S_AXIS_SCALAR_125_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_125_tkeep,
    input [S_AXIS_SCALAR_125_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_125_tstrb,
    input [S_AXIS_SCALAR_125_DIRECT_DMWIDTH-1:0] s_axis_scalar_125_tdata,
    output s_axis_scalar_125_tready,
    //input AXI-Stream to Scalar interface 126
    input s_axis_scalar_126_aclk,
    input s_axis_scalar_126_aresetn,
    input s_axis_scalar_126_tlast,
    input s_axis_scalar_126_tvalid,
    input [S_AXIS_SCALAR_126_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_126_tkeep,
    input [S_AXIS_SCALAR_126_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_126_tstrb,
    input [S_AXIS_SCALAR_126_DIRECT_DMWIDTH-1:0] s_axis_scalar_126_tdata,
    output s_axis_scalar_126_tready,
    //input AXI-Stream to Scalar interface 127
    input s_axis_scalar_127_aclk,
    input s_axis_scalar_127_aresetn,
    input s_axis_scalar_127_tlast,
    input s_axis_scalar_127_tvalid,
    input [S_AXIS_SCALAR_127_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_127_tkeep,
    input [S_AXIS_SCALAR_127_DIRECT_DMWIDTH/8-1:0] s_axis_scalar_127_tstrb,
    input [S_AXIS_SCALAR_127_DIRECT_DMWIDTH-1:0] s_axis_scalar_127_tdata,
    output s_axis_scalar_127_tready,
    //output scalar ports
    input [C_OUTPUT_SCALAR_0_WIDTH-1:0] ap_oscalar_0_din,
    input [C_OUTPUT_SCALAR_1_WIDTH-1:0] ap_oscalar_1_din,
    input [C_OUTPUT_SCALAR_2_WIDTH-1:0] ap_oscalar_2_din,
    input [C_OUTPUT_SCALAR_3_WIDTH-1:0] ap_oscalar_3_din,
    input [C_OUTPUT_SCALAR_4_WIDTH-1:0] ap_oscalar_4_din,
    input [C_OUTPUT_SCALAR_5_WIDTH-1:0] ap_oscalar_5_din,
    input [C_OUTPUT_SCALAR_6_WIDTH-1:0] ap_oscalar_6_din,
    input [C_OUTPUT_SCALAR_7_WIDTH-1:0] ap_oscalar_7_din,
    input [C_OUTPUT_SCALAR_8_WIDTH-1:0] ap_oscalar_8_din,
    input [C_OUTPUT_SCALAR_9_WIDTH-1:0] ap_oscalar_9_din,
    input [C_OUTPUT_SCALAR_10_WIDTH-1:0] ap_oscalar_10_din,
    input [C_OUTPUT_SCALAR_11_WIDTH-1:0] ap_oscalar_11_din,
    input [C_OUTPUT_SCALAR_12_WIDTH-1:0] ap_oscalar_12_din,
    input [C_OUTPUT_SCALAR_13_WIDTH-1:0] ap_oscalar_13_din,
    input [C_OUTPUT_SCALAR_14_WIDTH-1:0] ap_oscalar_14_din,
    input [C_OUTPUT_SCALAR_15_WIDTH-1:0] ap_oscalar_15_din,
    input [C_OUTPUT_SCALAR_16_WIDTH-1:0] ap_oscalar_16_din,
    input [C_OUTPUT_SCALAR_17_WIDTH-1:0] ap_oscalar_17_din,
    input [C_OUTPUT_SCALAR_18_WIDTH-1:0] ap_oscalar_18_din,
    input [C_OUTPUT_SCALAR_19_WIDTH-1:0] ap_oscalar_19_din,
    input [C_OUTPUT_SCALAR_20_WIDTH-1:0] ap_oscalar_20_din,
    input [C_OUTPUT_SCALAR_21_WIDTH-1:0] ap_oscalar_21_din,
    input [C_OUTPUT_SCALAR_22_WIDTH-1:0] ap_oscalar_22_din,
    input [C_OUTPUT_SCALAR_23_WIDTH-1:0] ap_oscalar_23_din,
    input [C_OUTPUT_SCALAR_24_WIDTH-1:0] ap_oscalar_24_din,
    input [C_OUTPUT_SCALAR_25_WIDTH-1:0] ap_oscalar_25_din,
    input [C_OUTPUT_SCALAR_26_WIDTH-1:0] ap_oscalar_26_din,
    input [C_OUTPUT_SCALAR_27_WIDTH-1:0] ap_oscalar_27_din,
    input [C_OUTPUT_SCALAR_28_WIDTH-1:0] ap_oscalar_28_din,
    input [C_OUTPUT_SCALAR_29_WIDTH-1:0] ap_oscalar_29_din,
    input [C_OUTPUT_SCALAR_30_WIDTH-1:0] ap_oscalar_30_din,
    input [C_OUTPUT_SCALAR_31_WIDTH-1:0] ap_oscalar_31_din,
    input [C_OUTPUT_SCALAR_32_WIDTH-1:0] ap_oscalar_32_din,
    input [C_OUTPUT_SCALAR_33_WIDTH-1:0] ap_oscalar_33_din,
    input [C_OUTPUT_SCALAR_34_WIDTH-1:0] ap_oscalar_34_din,
    input [C_OUTPUT_SCALAR_35_WIDTH-1:0] ap_oscalar_35_din,
    input [C_OUTPUT_SCALAR_36_WIDTH-1:0] ap_oscalar_36_din,
    input [C_OUTPUT_SCALAR_37_WIDTH-1:0] ap_oscalar_37_din,
    input [C_OUTPUT_SCALAR_38_WIDTH-1:0] ap_oscalar_38_din,
    input [C_OUTPUT_SCALAR_39_WIDTH-1:0] ap_oscalar_39_din,
    input [C_OUTPUT_SCALAR_40_WIDTH-1:0] ap_oscalar_40_din,
    input [C_OUTPUT_SCALAR_41_WIDTH-1:0] ap_oscalar_41_din,
    input [C_OUTPUT_SCALAR_42_WIDTH-1:0] ap_oscalar_42_din,
    input [C_OUTPUT_SCALAR_43_WIDTH-1:0] ap_oscalar_43_din,
    input [C_OUTPUT_SCALAR_44_WIDTH-1:0] ap_oscalar_44_din,
    input [C_OUTPUT_SCALAR_45_WIDTH-1:0] ap_oscalar_45_din,
    input [C_OUTPUT_SCALAR_46_WIDTH-1:0] ap_oscalar_46_din,
    input [C_OUTPUT_SCALAR_47_WIDTH-1:0] ap_oscalar_47_din,
    input [C_OUTPUT_SCALAR_48_WIDTH-1:0] ap_oscalar_48_din,
    input [C_OUTPUT_SCALAR_49_WIDTH-1:0] ap_oscalar_49_din,
    input [C_OUTPUT_SCALAR_50_WIDTH-1:0] ap_oscalar_50_din,
    input [C_OUTPUT_SCALAR_51_WIDTH-1:0] ap_oscalar_51_din,
    input [C_OUTPUT_SCALAR_52_WIDTH-1:0] ap_oscalar_52_din,
    input [C_OUTPUT_SCALAR_53_WIDTH-1:0] ap_oscalar_53_din,
    input [C_OUTPUT_SCALAR_54_WIDTH-1:0] ap_oscalar_54_din,
    input [C_OUTPUT_SCALAR_55_WIDTH-1:0] ap_oscalar_55_din,
    input [C_OUTPUT_SCALAR_56_WIDTH-1:0] ap_oscalar_56_din,
    input [C_OUTPUT_SCALAR_57_WIDTH-1:0] ap_oscalar_57_din,
    input [C_OUTPUT_SCALAR_58_WIDTH-1:0] ap_oscalar_58_din,
    input [C_OUTPUT_SCALAR_59_WIDTH-1:0] ap_oscalar_59_din,
    input [C_OUTPUT_SCALAR_60_WIDTH-1:0] ap_oscalar_60_din,
    input [C_OUTPUT_SCALAR_61_WIDTH-1:0] ap_oscalar_61_din,
    input [C_OUTPUT_SCALAR_62_WIDTH-1:0] ap_oscalar_62_din,
    input [C_OUTPUT_SCALAR_63_WIDTH-1:0] ap_oscalar_63_din,
    input [C_OUTPUT_SCALAR_64_WIDTH-1:0] ap_oscalar_64_din,
    input [C_OUTPUT_SCALAR_65_WIDTH-1:0] ap_oscalar_65_din,
    input [C_OUTPUT_SCALAR_66_WIDTH-1:0] ap_oscalar_66_din,
    input [C_OUTPUT_SCALAR_67_WIDTH-1:0] ap_oscalar_67_din,
    input [C_OUTPUT_SCALAR_68_WIDTH-1:0] ap_oscalar_68_din,
    input [C_OUTPUT_SCALAR_69_WIDTH-1:0] ap_oscalar_69_din,
    input [C_OUTPUT_SCALAR_70_WIDTH-1:0] ap_oscalar_70_din,
    input [C_OUTPUT_SCALAR_71_WIDTH-1:0] ap_oscalar_71_din,
    input [C_OUTPUT_SCALAR_72_WIDTH-1:0] ap_oscalar_72_din,
    input [C_OUTPUT_SCALAR_73_WIDTH-1:0] ap_oscalar_73_din,
    input [C_OUTPUT_SCALAR_74_WIDTH-1:0] ap_oscalar_74_din,
    input [C_OUTPUT_SCALAR_75_WIDTH-1:0] ap_oscalar_75_din,
    input [C_OUTPUT_SCALAR_76_WIDTH-1:0] ap_oscalar_76_din,
    input [C_OUTPUT_SCALAR_77_WIDTH-1:0] ap_oscalar_77_din,
    input [C_OUTPUT_SCALAR_78_WIDTH-1:0] ap_oscalar_78_din,
    input [C_OUTPUT_SCALAR_79_WIDTH-1:0] ap_oscalar_79_din,
    input [C_OUTPUT_SCALAR_80_WIDTH-1:0] ap_oscalar_80_din,
    input [C_OUTPUT_SCALAR_81_WIDTH-1:0] ap_oscalar_81_din,
    input [C_OUTPUT_SCALAR_82_WIDTH-1:0] ap_oscalar_82_din,
    input [C_OUTPUT_SCALAR_83_WIDTH-1:0] ap_oscalar_83_din,
    input [C_OUTPUT_SCALAR_84_WIDTH-1:0] ap_oscalar_84_din,
    input [C_OUTPUT_SCALAR_85_WIDTH-1:0] ap_oscalar_85_din,
    input [C_OUTPUT_SCALAR_86_WIDTH-1:0] ap_oscalar_86_din,
    input [C_OUTPUT_SCALAR_87_WIDTH-1:0] ap_oscalar_87_din,
    input [C_OUTPUT_SCALAR_88_WIDTH-1:0] ap_oscalar_88_din,
    input [C_OUTPUT_SCALAR_89_WIDTH-1:0] ap_oscalar_89_din,
    input [C_OUTPUT_SCALAR_90_WIDTH-1:0] ap_oscalar_90_din,
    input [C_OUTPUT_SCALAR_91_WIDTH-1:0] ap_oscalar_91_din,
    input [C_OUTPUT_SCALAR_92_WIDTH-1:0] ap_oscalar_92_din,
    input [C_OUTPUT_SCALAR_93_WIDTH-1:0] ap_oscalar_93_din,
    input [C_OUTPUT_SCALAR_94_WIDTH-1:0] ap_oscalar_94_din,
    input [C_OUTPUT_SCALAR_95_WIDTH-1:0] ap_oscalar_95_din,
    input [C_OUTPUT_SCALAR_96_WIDTH-1:0] ap_oscalar_96_din,
    input [C_OUTPUT_SCALAR_97_WIDTH-1:0] ap_oscalar_97_din,
    input [C_OUTPUT_SCALAR_98_WIDTH-1:0] ap_oscalar_98_din,
    input [C_OUTPUT_SCALAR_99_WIDTH-1:0] ap_oscalar_99_din,
    input [C_OUTPUT_SCALAR_100_WIDTH-1:0] ap_oscalar_100_din,
    input [C_OUTPUT_SCALAR_101_WIDTH-1:0] ap_oscalar_101_din,
    input [C_OUTPUT_SCALAR_102_WIDTH-1:0] ap_oscalar_102_din,
    input [C_OUTPUT_SCALAR_103_WIDTH-1:0] ap_oscalar_103_din,
    input [C_OUTPUT_SCALAR_104_WIDTH-1:0] ap_oscalar_104_din,
    input [C_OUTPUT_SCALAR_105_WIDTH-1:0] ap_oscalar_105_din,
    input [C_OUTPUT_SCALAR_106_WIDTH-1:0] ap_oscalar_106_din,
    input [C_OUTPUT_SCALAR_107_WIDTH-1:0] ap_oscalar_107_din,
    input [C_OUTPUT_SCALAR_108_WIDTH-1:0] ap_oscalar_108_din,
    input [C_OUTPUT_SCALAR_109_WIDTH-1:0] ap_oscalar_109_din,
    input [C_OUTPUT_SCALAR_110_WIDTH-1:0] ap_oscalar_110_din,
    input [C_OUTPUT_SCALAR_111_WIDTH-1:0] ap_oscalar_111_din,
    input [C_OUTPUT_SCALAR_112_WIDTH-1:0] ap_oscalar_112_din,
    input [C_OUTPUT_SCALAR_113_WIDTH-1:0] ap_oscalar_113_din,
    input [C_OUTPUT_SCALAR_114_WIDTH-1:0] ap_oscalar_114_din,
    input [C_OUTPUT_SCALAR_115_WIDTH-1:0] ap_oscalar_115_din,
    input [C_OUTPUT_SCALAR_116_WIDTH-1:0] ap_oscalar_116_din,
    input [C_OUTPUT_SCALAR_117_WIDTH-1:0] ap_oscalar_117_din,
    input [C_OUTPUT_SCALAR_118_WIDTH-1:0] ap_oscalar_118_din,
    input [C_OUTPUT_SCALAR_119_WIDTH-1:0] ap_oscalar_119_din,
    input [C_OUTPUT_SCALAR_120_WIDTH-1:0] ap_oscalar_120_din,
    input [C_OUTPUT_SCALAR_121_WIDTH-1:0] ap_oscalar_121_din,
    input [C_OUTPUT_SCALAR_122_WIDTH-1:0] ap_oscalar_122_din,
    input [C_OUTPUT_SCALAR_123_WIDTH-1:0] ap_oscalar_123_din,
    input [C_OUTPUT_SCALAR_124_WIDTH-1:0] ap_oscalar_124_din,
    input [C_OUTPUT_SCALAR_125_WIDTH-1:0] ap_oscalar_125_din,
    input [C_OUTPUT_SCALAR_126_WIDTH-1:0] ap_oscalar_126_din,
    input [C_OUTPUT_SCALAR_127_WIDTH-1:0] ap_oscalar_127_din,
    //output scalar valid ports
    input ap_oscalar_0_vld,
    input ap_oscalar_1_vld,
    input ap_oscalar_2_vld,
    input ap_oscalar_3_vld,
    input ap_oscalar_4_vld,
    input ap_oscalar_5_vld,
    input ap_oscalar_6_vld,
    input ap_oscalar_7_vld,
    input ap_oscalar_8_vld,
    input ap_oscalar_9_vld,
    input ap_oscalar_10_vld,
    input ap_oscalar_11_vld,
    input ap_oscalar_12_vld,
    input ap_oscalar_13_vld,
    input ap_oscalar_14_vld,
    input ap_oscalar_15_vld,
    input ap_oscalar_16_vld,
    input ap_oscalar_17_vld,
    input ap_oscalar_18_vld,
    input ap_oscalar_19_vld,
    input ap_oscalar_20_vld,
    input ap_oscalar_21_vld,
    input ap_oscalar_22_vld,
    input ap_oscalar_23_vld,
    input ap_oscalar_24_vld,
    input ap_oscalar_25_vld,
    input ap_oscalar_26_vld,
    input ap_oscalar_27_vld,
    input ap_oscalar_28_vld,
    input ap_oscalar_29_vld,
    input ap_oscalar_30_vld,
    input ap_oscalar_31_vld,
    input ap_oscalar_32_vld,
    input ap_oscalar_33_vld,
    input ap_oscalar_34_vld,
    input ap_oscalar_35_vld,
    input ap_oscalar_36_vld,
    input ap_oscalar_37_vld,
    input ap_oscalar_38_vld,
    input ap_oscalar_39_vld,
    input ap_oscalar_40_vld,
    input ap_oscalar_41_vld,
    input ap_oscalar_42_vld,
    input ap_oscalar_43_vld,
    input ap_oscalar_44_vld,
    input ap_oscalar_45_vld,
    input ap_oscalar_46_vld,
    input ap_oscalar_47_vld,
    input ap_oscalar_48_vld,
    input ap_oscalar_49_vld,
    input ap_oscalar_50_vld,
    input ap_oscalar_51_vld,
    input ap_oscalar_52_vld,
    input ap_oscalar_53_vld,
    input ap_oscalar_54_vld,
    input ap_oscalar_55_vld,
    input ap_oscalar_56_vld,
    input ap_oscalar_57_vld,
    input ap_oscalar_58_vld,
    input ap_oscalar_59_vld,
    input ap_oscalar_60_vld,
    input ap_oscalar_61_vld,
    input ap_oscalar_62_vld,
    input ap_oscalar_63_vld,
    input ap_oscalar_64_vld,
    input ap_oscalar_65_vld,
    input ap_oscalar_66_vld,
    input ap_oscalar_67_vld,
    input ap_oscalar_68_vld,
    input ap_oscalar_69_vld,
    input ap_oscalar_70_vld,
    input ap_oscalar_71_vld,
    input ap_oscalar_72_vld,
    input ap_oscalar_73_vld,
    input ap_oscalar_74_vld,
    input ap_oscalar_75_vld,
    input ap_oscalar_76_vld,
    input ap_oscalar_77_vld,
    input ap_oscalar_78_vld,
    input ap_oscalar_79_vld,
    input ap_oscalar_80_vld,
    input ap_oscalar_81_vld,
    input ap_oscalar_82_vld,
    input ap_oscalar_83_vld,
    input ap_oscalar_84_vld,
    input ap_oscalar_85_vld,
    input ap_oscalar_86_vld,
    input ap_oscalar_87_vld,
    input ap_oscalar_88_vld,
    input ap_oscalar_89_vld,
    input ap_oscalar_90_vld,
    input ap_oscalar_91_vld,
    input ap_oscalar_92_vld,
    input ap_oscalar_93_vld,
    input ap_oscalar_94_vld,
    input ap_oscalar_95_vld,
    input ap_oscalar_96_vld,
    input ap_oscalar_97_vld,
    input ap_oscalar_98_vld,
    input ap_oscalar_99_vld,
    input ap_oscalar_100_vld,
    input ap_oscalar_101_vld,
    input ap_oscalar_102_vld,
    input ap_oscalar_103_vld,
    input ap_oscalar_104_vld,
    input ap_oscalar_105_vld,
    input ap_oscalar_106_vld,
    input ap_oscalar_107_vld,
    input ap_oscalar_108_vld,
    input ap_oscalar_109_vld,
    input ap_oscalar_110_vld,
    input ap_oscalar_111_vld,
    input ap_oscalar_112_vld,
    input ap_oscalar_113_vld,
    input ap_oscalar_114_vld,
    input ap_oscalar_115_vld,
    input ap_oscalar_116_vld,
    input ap_oscalar_117_vld,
    input ap_oscalar_118_vld,
    input ap_oscalar_119_vld,
    input ap_oscalar_120_vld,
    input ap_oscalar_121_vld,
    input ap_oscalar_122_vld,
    input ap_oscalar_123_vld,
    input ap_oscalar_124_vld,
    input ap_oscalar_125_vld,
    input ap_oscalar_126_vld,
    input ap_oscalar_127_vld,
    //output Scalar to AXI-Stream interface 0
    input m_axis_scalar_0_aclk,
    input m_axis_scalar_0_aresetn,
    output m_axis_scalar_0_tlast,
    output m_axis_scalar_0_tvalid,
    output [M_AXIS_SCALAR_0_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_0_tkeep,
    output [M_AXIS_SCALAR_0_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_0_tstrb,
    output [M_AXIS_SCALAR_0_DIRECT_DMWIDTH-1:0] m_axis_scalar_0_tdata,
    input m_axis_scalar_0_tready,
    //output Scalar to AXI-Stream interface 1
    input m_axis_scalar_1_aclk,
    input m_axis_scalar_1_aresetn,
    output m_axis_scalar_1_tlast,
    output m_axis_scalar_1_tvalid,
    output [M_AXIS_SCALAR_1_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_1_tkeep,
    output [M_AXIS_SCALAR_1_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_1_tstrb,
    output [M_AXIS_SCALAR_1_DIRECT_DMWIDTH-1:0] m_axis_scalar_1_tdata,
    input m_axis_scalar_1_tready,
    //output Scalar to AXI-Stream interface 2
    input m_axis_scalar_2_aclk,
    input m_axis_scalar_2_aresetn,
    output m_axis_scalar_2_tlast,
    output m_axis_scalar_2_tvalid,
    output [M_AXIS_SCALAR_2_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_2_tkeep,
    output [M_AXIS_SCALAR_2_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_2_tstrb,
    output [M_AXIS_SCALAR_2_DIRECT_DMWIDTH-1:0] m_axis_scalar_2_tdata,
    input m_axis_scalar_2_tready,
    //output Scalar to AXI-Stream interface 3
    input m_axis_scalar_3_aclk,
    input m_axis_scalar_3_aresetn,
    output m_axis_scalar_3_tlast,
    output m_axis_scalar_3_tvalid,
    output [M_AXIS_SCALAR_3_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_3_tkeep,
    output [M_AXIS_SCALAR_3_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_3_tstrb,
    output [M_AXIS_SCALAR_3_DIRECT_DMWIDTH-1:0] m_axis_scalar_3_tdata,
    input m_axis_scalar_3_tready,
    //output Scalar to AXI-Stream interface 4
    input m_axis_scalar_4_aclk,
    input m_axis_scalar_4_aresetn,
    output m_axis_scalar_4_tlast,
    output m_axis_scalar_4_tvalid,
    output [M_AXIS_SCALAR_4_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_4_tkeep,
    output [M_AXIS_SCALAR_4_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_4_tstrb,
    output [M_AXIS_SCALAR_4_DIRECT_DMWIDTH-1:0] m_axis_scalar_4_tdata,
    input m_axis_scalar_4_tready,
    //output Scalar to AXI-Stream interface 5
    input m_axis_scalar_5_aclk,
    input m_axis_scalar_5_aresetn,
    output m_axis_scalar_5_tlast,
    output m_axis_scalar_5_tvalid,
    output [M_AXIS_SCALAR_5_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_5_tkeep,
    output [M_AXIS_SCALAR_5_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_5_tstrb,
    output [M_AXIS_SCALAR_5_DIRECT_DMWIDTH-1:0] m_axis_scalar_5_tdata,
    input m_axis_scalar_5_tready,
    //output Scalar to AXI-Stream interface 6
    input m_axis_scalar_6_aclk,
    input m_axis_scalar_6_aresetn,
    output m_axis_scalar_6_tlast,
    output m_axis_scalar_6_tvalid,
    output [M_AXIS_SCALAR_6_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_6_tkeep,
    output [M_AXIS_SCALAR_6_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_6_tstrb,
    output [M_AXIS_SCALAR_6_DIRECT_DMWIDTH-1:0] m_axis_scalar_6_tdata,
    input m_axis_scalar_6_tready,
    //output Scalar to AXI-Stream interface 7
    input m_axis_scalar_7_aclk,
    input m_axis_scalar_7_aresetn,
    output m_axis_scalar_7_tlast,
    output m_axis_scalar_7_tvalid,
    output [M_AXIS_SCALAR_7_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_7_tkeep,
    output [M_AXIS_SCALAR_7_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_7_tstrb,
    output [M_AXIS_SCALAR_7_DIRECT_DMWIDTH-1:0] m_axis_scalar_7_tdata,
    input m_axis_scalar_7_tready,
    //output Scalar to AXI-Stream interface 8
    input m_axis_scalar_8_aclk,
    input m_axis_scalar_8_aresetn,
    output m_axis_scalar_8_tlast,
    output m_axis_scalar_8_tvalid,
    output [M_AXIS_SCALAR_8_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_8_tkeep,
    output [M_AXIS_SCALAR_8_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_8_tstrb,
    output [M_AXIS_SCALAR_8_DIRECT_DMWIDTH-1:0] m_axis_scalar_8_tdata,
    input m_axis_scalar_8_tready,
    //output Scalar to AXI-Stream interface 9
    input m_axis_scalar_9_aclk,
    input m_axis_scalar_9_aresetn,
    output m_axis_scalar_9_tlast,
    output m_axis_scalar_9_tvalid,
    output [M_AXIS_SCALAR_9_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_9_tkeep,
    output [M_AXIS_SCALAR_9_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_9_tstrb,
    output [M_AXIS_SCALAR_9_DIRECT_DMWIDTH-1:0] m_axis_scalar_9_tdata,
    input m_axis_scalar_9_tready,
    //output Scalar to AXI-Stream interface 10
    input m_axis_scalar_10_aclk,
    input m_axis_scalar_10_aresetn,
    output m_axis_scalar_10_tlast,
    output m_axis_scalar_10_tvalid,
    output [M_AXIS_SCALAR_10_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_10_tkeep,
    output [M_AXIS_SCALAR_10_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_10_tstrb,
    output [M_AXIS_SCALAR_10_DIRECT_DMWIDTH-1:0] m_axis_scalar_10_tdata,
    input m_axis_scalar_10_tready,
    //output Scalar to AXI-Stream interface 11
    input m_axis_scalar_11_aclk,
    input m_axis_scalar_11_aresetn,
    output m_axis_scalar_11_tlast,
    output m_axis_scalar_11_tvalid,
    output [M_AXIS_SCALAR_11_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_11_tkeep,
    output [M_AXIS_SCALAR_11_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_11_tstrb,
    output [M_AXIS_SCALAR_11_DIRECT_DMWIDTH-1:0] m_axis_scalar_11_tdata,
    input m_axis_scalar_11_tready,
    //output Scalar to AXI-Stream interface 12
    input m_axis_scalar_12_aclk,
    input m_axis_scalar_12_aresetn,
    output m_axis_scalar_12_tlast,
    output m_axis_scalar_12_tvalid,
    output [M_AXIS_SCALAR_12_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_12_tkeep,
    output [M_AXIS_SCALAR_12_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_12_tstrb,
    output [M_AXIS_SCALAR_12_DIRECT_DMWIDTH-1:0] m_axis_scalar_12_tdata,
    input m_axis_scalar_12_tready,
    //output Scalar to AXI-Stream interface 13
    input m_axis_scalar_13_aclk,
    input m_axis_scalar_13_aresetn,
    output m_axis_scalar_13_tlast,
    output m_axis_scalar_13_tvalid,
    output [M_AXIS_SCALAR_13_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_13_tkeep,
    output [M_AXIS_SCALAR_13_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_13_tstrb,
    output [M_AXIS_SCALAR_13_DIRECT_DMWIDTH-1:0] m_axis_scalar_13_tdata,
    input m_axis_scalar_13_tready,
    //output Scalar to AXI-Stream interface 14
    input m_axis_scalar_14_aclk,
    input m_axis_scalar_14_aresetn,
    output m_axis_scalar_14_tlast,
    output m_axis_scalar_14_tvalid,
    output [M_AXIS_SCALAR_14_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_14_tkeep,
    output [M_AXIS_SCALAR_14_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_14_tstrb,
    output [M_AXIS_SCALAR_14_DIRECT_DMWIDTH-1:0] m_axis_scalar_14_tdata,
    input m_axis_scalar_14_tready,
    //output Scalar to AXI-Stream interface 15
    input m_axis_scalar_15_aclk,
    input m_axis_scalar_15_aresetn,
    output m_axis_scalar_15_tlast,
    output m_axis_scalar_15_tvalid,
    output [M_AXIS_SCALAR_15_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_15_tkeep,
    output [M_AXIS_SCALAR_15_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_15_tstrb,
    output [M_AXIS_SCALAR_15_DIRECT_DMWIDTH-1:0] m_axis_scalar_15_tdata,
    input m_axis_scalar_15_tready,
    //output Scalar to AXI-Stream interface 16
    input m_axis_scalar_16_aclk,
    input m_axis_scalar_16_aresetn,
    output m_axis_scalar_16_tlast,
    output m_axis_scalar_16_tvalid,
    output [M_AXIS_SCALAR_16_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_16_tkeep,
    output [M_AXIS_SCALAR_16_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_16_tstrb,
    output [M_AXIS_SCALAR_16_DIRECT_DMWIDTH-1:0] m_axis_scalar_16_tdata,
    input m_axis_scalar_16_tready,
    //output Scalar to AXI-Stream interface 17
    input m_axis_scalar_17_aclk,
    input m_axis_scalar_17_aresetn,
    output m_axis_scalar_17_tlast,
    output m_axis_scalar_17_tvalid,
    output [M_AXIS_SCALAR_17_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_17_tkeep,
    output [M_AXIS_SCALAR_17_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_17_tstrb,
    output [M_AXIS_SCALAR_17_DIRECT_DMWIDTH-1:0] m_axis_scalar_17_tdata,
    input m_axis_scalar_17_tready,
    //output Scalar to AXI-Stream interface 18
    input m_axis_scalar_18_aclk,
    input m_axis_scalar_18_aresetn,
    output m_axis_scalar_18_tlast,
    output m_axis_scalar_18_tvalid,
    output [M_AXIS_SCALAR_18_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_18_tkeep,
    output [M_AXIS_SCALAR_18_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_18_tstrb,
    output [M_AXIS_SCALAR_18_DIRECT_DMWIDTH-1:0] m_axis_scalar_18_tdata,
    input m_axis_scalar_18_tready,
    //output Scalar to AXI-Stream interface 19
    input m_axis_scalar_19_aclk,
    input m_axis_scalar_19_aresetn,
    output m_axis_scalar_19_tlast,
    output m_axis_scalar_19_tvalid,
    output [M_AXIS_SCALAR_19_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_19_tkeep,
    output [M_AXIS_SCALAR_19_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_19_tstrb,
    output [M_AXIS_SCALAR_19_DIRECT_DMWIDTH-1:0] m_axis_scalar_19_tdata,
    input m_axis_scalar_19_tready,
    //output Scalar to AXI-Stream interface 20
    input m_axis_scalar_20_aclk,
    input m_axis_scalar_20_aresetn,
    output m_axis_scalar_20_tlast,
    output m_axis_scalar_20_tvalid,
    output [M_AXIS_SCALAR_20_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_20_tkeep,
    output [M_AXIS_SCALAR_20_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_20_tstrb,
    output [M_AXIS_SCALAR_20_DIRECT_DMWIDTH-1:0] m_axis_scalar_20_tdata,
    input m_axis_scalar_20_tready,
    //output Scalar to AXI-Stream interface 21
    input m_axis_scalar_21_aclk,
    input m_axis_scalar_21_aresetn,
    output m_axis_scalar_21_tlast,
    output m_axis_scalar_21_tvalid,
    output [M_AXIS_SCALAR_21_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_21_tkeep,
    output [M_AXIS_SCALAR_21_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_21_tstrb,
    output [M_AXIS_SCALAR_21_DIRECT_DMWIDTH-1:0] m_axis_scalar_21_tdata,
    input m_axis_scalar_21_tready,
    //output Scalar to AXI-Stream interface 22
    input m_axis_scalar_22_aclk,
    input m_axis_scalar_22_aresetn,
    output m_axis_scalar_22_tlast,
    output m_axis_scalar_22_tvalid,
    output [M_AXIS_SCALAR_22_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_22_tkeep,
    output [M_AXIS_SCALAR_22_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_22_tstrb,
    output [M_AXIS_SCALAR_22_DIRECT_DMWIDTH-1:0] m_axis_scalar_22_tdata,
    input m_axis_scalar_22_tready,
    //output Scalar to AXI-Stream interface 23
    input m_axis_scalar_23_aclk,
    input m_axis_scalar_23_aresetn,
    output m_axis_scalar_23_tlast,
    output m_axis_scalar_23_tvalid,
    output [M_AXIS_SCALAR_23_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_23_tkeep,
    output [M_AXIS_SCALAR_23_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_23_tstrb,
    output [M_AXIS_SCALAR_23_DIRECT_DMWIDTH-1:0] m_axis_scalar_23_tdata,
    input m_axis_scalar_23_tready,
    //output Scalar to AXI-Stream interface 24
    input m_axis_scalar_24_aclk,
    input m_axis_scalar_24_aresetn,
    output m_axis_scalar_24_tlast,
    output m_axis_scalar_24_tvalid,
    output [M_AXIS_SCALAR_24_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_24_tkeep,
    output [M_AXIS_SCALAR_24_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_24_tstrb,
    output [M_AXIS_SCALAR_24_DIRECT_DMWIDTH-1:0] m_axis_scalar_24_tdata,
    input m_axis_scalar_24_tready,
    //output Scalar to AXI-Stream interface 25
    input m_axis_scalar_25_aclk,
    input m_axis_scalar_25_aresetn,
    output m_axis_scalar_25_tlast,
    output m_axis_scalar_25_tvalid,
    output [M_AXIS_SCALAR_25_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_25_tkeep,
    output [M_AXIS_SCALAR_25_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_25_tstrb,
    output [M_AXIS_SCALAR_25_DIRECT_DMWIDTH-1:0] m_axis_scalar_25_tdata,
    input m_axis_scalar_25_tready,
    //output Scalar to AXI-Stream interface 26
    input m_axis_scalar_26_aclk,
    input m_axis_scalar_26_aresetn,
    output m_axis_scalar_26_tlast,
    output m_axis_scalar_26_tvalid,
    output [M_AXIS_SCALAR_26_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_26_tkeep,
    output [M_AXIS_SCALAR_26_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_26_tstrb,
    output [M_AXIS_SCALAR_26_DIRECT_DMWIDTH-1:0] m_axis_scalar_26_tdata,
    input m_axis_scalar_26_tready,
    //output Scalar to AXI-Stream interface 27
    input m_axis_scalar_27_aclk,
    input m_axis_scalar_27_aresetn,
    output m_axis_scalar_27_tlast,
    output m_axis_scalar_27_tvalid,
    output [M_AXIS_SCALAR_27_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_27_tkeep,
    output [M_AXIS_SCALAR_27_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_27_tstrb,
    output [M_AXIS_SCALAR_27_DIRECT_DMWIDTH-1:0] m_axis_scalar_27_tdata,
    input m_axis_scalar_27_tready,
    //output Scalar to AXI-Stream interface 28
    input m_axis_scalar_28_aclk,
    input m_axis_scalar_28_aresetn,
    output m_axis_scalar_28_tlast,
    output m_axis_scalar_28_tvalid,
    output [M_AXIS_SCALAR_28_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_28_tkeep,
    output [M_AXIS_SCALAR_28_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_28_tstrb,
    output [M_AXIS_SCALAR_28_DIRECT_DMWIDTH-1:0] m_axis_scalar_28_tdata,
    input m_axis_scalar_28_tready,
    //output Scalar to AXI-Stream interface 29
    input m_axis_scalar_29_aclk,
    input m_axis_scalar_29_aresetn,
    output m_axis_scalar_29_tlast,
    output m_axis_scalar_29_tvalid,
    output [M_AXIS_SCALAR_29_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_29_tkeep,
    output [M_AXIS_SCALAR_29_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_29_tstrb,
    output [M_AXIS_SCALAR_29_DIRECT_DMWIDTH-1:0] m_axis_scalar_29_tdata,
    input m_axis_scalar_29_tready,
    //output Scalar to AXI-Stream interface 30
    input m_axis_scalar_30_aclk,
    input m_axis_scalar_30_aresetn,
    output m_axis_scalar_30_tlast,
    output m_axis_scalar_30_tvalid,
    output [M_AXIS_SCALAR_30_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_30_tkeep,
    output [M_AXIS_SCALAR_30_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_30_tstrb,
    output [M_AXIS_SCALAR_30_DIRECT_DMWIDTH-1:0] m_axis_scalar_30_tdata,
    input m_axis_scalar_30_tready,
    //output Scalar to AXI-Stream interface 31
    input m_axis_scalar_31_aclk,
    input m_axis_scalar_31_aresetn,
    output m_axis_scalar_31_tlast,
    output m_axis_scalar_31_tvalid,
    output [M_AXIS_SCALAR_31_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_31_tkeep,
    output [M_AXIS_SCALAR_31_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_31_tstrb,
    output [M_AXIS_SCALAR_31_DIRECT_DMWIDTH-1:0] m_axis_scalar_31_tdata,
    input m_axis_scalar_31_tready,
    //output Scalar to AXI-Stream interface 32
    input m_axis_scalar_32_aclk,
    input m_axis_scalar_32_aresetn,
    output m_axis_scalar_32_tlast,
    output m_axis_scalar_32_tvalid,
    output [M_AXIS_SCALAR_32_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_32_tkeep,
    output [M_AXIS_SCALAR_32_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_32_tstrb,
    output [M_AXIS_SCALAR_32_DIRECT_DMWIDTH-1:0] m_axis_scalar_32_tdata,
    input m_axis_scalar_32_tready,
    //output Scalar to AXI-Stream interface 33
    input m_axis_scalar_33_aclk,
    input m_axis_scalar_33_aresetn,
    output m_axis_scalar_33_tlast,
    output m_axis_scalar_33_tvalid,
    output [M_AXIS_SCALAR_33_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_33_tkeep,
    output [M_AXIS_SCALAR_33_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_33_tstrb,
    output [M_AXIS_SCALAR_33_DIRECT_DMWIDTH-1:0] m_axis_scalar_33_tdata,
    input m_axis_scalar_33_tready,
    //output Scalar to AXI-Stream interface 34
    input m_axis_scalar_34_aclk,
    input m_axis_scalar_34_aresetn,
    output m_axis_scalar_34_tlast,
    output m_axis_scalar_34_tvalid,
    output [M_AXIS_SCALAR_34_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_34_tkeep,
    output [M_AXIS_SCALAR_34_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_34_tstrb,
    output [M_AXIS_SCALAR_34_DIRECT_DMWIDTH-1:0] m_axis_scalar_34_tdata,
    input m_axis_scalar_34_tready,
    //output Scalar to AXI-Stream interface 35
    input m_axis_scalar_35_aclk,
    input m_axis_scalar_35_aresetn,
    output m_axis_scalar_35_tlast,
    output m_axis_scalar_35_tvalid,
    output [M_AXIS_SCALAR_35_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_35_tkeep,
    output [M_AXIS_SCALAR_35_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_35_tstrb,
    output [M_AXIS_SCALAR_35_DIRECT_DMWIDTH-1:0] m_axis_scalar_35_tdata,
    input m_axis_scalar_35_tready,
    //output Scalar to AXI-Stream interface 36
    input m_axis_scalar_36_aclk,
    input m_axis_scalar_36_aresetn,
    output m_axis_scalar_36_tlast,
    output m_axis_scalar_36_tvalid,
    output [M_AXIS_SCALAR_36_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_36_tkeep,
    output [M_AXIS_SCALAR_36_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_36_tstrb,
    output [M_AXIS_SCALAR_36_DIRECT_DMWIDTH-1:0] m_axis_scalar_36_tdata,
    input m_axis_scalar_36_tready,
    //output Scalar to AXI-Stream interface 37
    input m_axis_scalar_37_aclk,
    input m_axis_scalar_37_aresetn,
    output m_axis_scalar_37_tlast,
    output m_axis_scalar_37_tvalid,
    output [M_AXIS_SCALAR_37_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_37_tkeep,
    output [M_AXIS_SCALAR_37_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_37_tstrb,
    output [M_AXIS_SCALAR_37_DIRECT_DMWIDTH-1:0] m_axis_scalar_37_tdata,
    input m_axis_scalar_37_tready,
    //output Scalar to AXI-Stream interface 38
    input m_axis_scalar_38_aclk,
    input m_axis_scalar_38_aresetn,
    output m_axis_scalar_38_tlast,
    output m_axis_scalar_38_tvalid,
    output [M_AXIS_SCALAR_38_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_38_tkeep,
    output [M_AXIS_SCALAR_38_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_38_tstrb,
    output [M_AXIS_SCALAR_38_DIRECT_DMWIDTH-1:0] m_axis_scalar_38_tdata,
    input m_axis_scalar_38_tready,
    //output Scalar to AXI-Stream interface 39
    input m_axis_scalar_39_aclk,
    input m_axis_scalar_39_aresetn,
    output m_axis_scalar_39_tlast,
    output m_axis_scalar_39_tvalid,
    output [M_AXIS_SCALAR_39_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_39_tkeep,
    output [M_AXIS_SCALAR_39_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_39_tstrb,
    output [M_AXIS_SCALAR_39_DIRECT_DMWIDTH-1:0] m_axis_scalar_39_tdata,
    input m_axis_scalar_39_tready,
    //output Scalar to AXI-Stream interface 40
    input m_axis_scalar_40_aclk,
    input m_axis_scalar_40_aresetn,
    output m_axis_scalar_40_tlast,
    output m_axis_scalar_40_tvalid,
    output [M_AXIS_SCALAR_40_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_40_tkeep,
    output [M_AXIS_SCALAR_40_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_40_tstrb,
    output [M_AXIS_SCALAR_40_DIRECT_DMWIDTH-1:0] m_axis_scalar_40_tdata,
    input m_axis_scalar_40_tready,
    //output Scalar to AXI-Stream interface 41
    input m_axis_scalar_41_aclk,
    input m_axis_scalar_41_aresetn,
    output m_axis_scalar_41_tlast,
    output m_axis_scalar_41_tvalid,
    output [M_AXIS_SCALAR_41_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_41_tkeep,
    output [M_AXIS_SCALAR_41_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_41_tstrb,
    output [M_AXIS_SCALAR_41_DIRECT_DMWIDTH-1:0] m_axis_scalar_41_tdata,
    input m_axis_scalar_41_tready,
    //output Scalar to AXI-Stream interface 42
    input m_axis_scalar_42_aclk,
    input m_axis_scalar_42_aresetn,
    output m_axis_scalar_42_tlast,
    output m_axis_scalar_42_tvalid,
    output [M_AXIS_SCALAR_42_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_42_tkeep,
    output [M_AXIS_SCALAR_42_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_42_tstrb,
    output [M_AXIS_SCALAR_42_DIRECT_DMWIDTH-1:0] m_axis_scalar_42_tdata,
    input m_axis_scalar_42_tready,
    //output Scalar to AXI-Stream interface 43
    input m_axis_scalar_43_aclk,
    input m_axis_scalar_43_aresetn,
    output m_axis_scalar_43_tlast,
    output m_axis_scalar_43_tvalid,
    output [M_AXIS_SCALAR_43_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_43_tkeep,
    output [M_AXIS_SCALAR_43_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_43_tstrb,
    output [M_AXIS_SCALAR_43_DIRECT_DMWIDTH-1:0] m_axis_scalar_43_tdata,
    input m_axis_scalar_43_tready,
    //output Scalar to AXI-Stream interface 44
    input m_axis_scalar_44_aclk,
    input m_axis_scalar_44_aresetn,
    output m_axis_scalar_44_tlast,
    output m_axis_scalar_44_tvalid,
    output [M_AXIS_SCALAR_44_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_44_tkeep,
    output [M_AXIS_SCALAR_44_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_44_tstrb,
    output [M_AXIS_SCALAR_44_DIRECT_DMWIDTH-1:0] m_axis_scalar_44_tdata,
    input m_axis_scalar_44_tready,
    //output Scalar to AXI-Stream interface 45
    input m_axis_scalar_45_aclk,
    input m_axis_scalar_45_aresetn,
    output m_axis_scalar_45_tlast,
    output m_axis_scalar_45_tvalid,
    output [M_AXIS_SCALAR_45_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_45_tkeep,
    output [M_AXIS_SCALAR_45_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_45_tstrb,
    output [M_AXIS_SCALAR_45_DIRECT_DMWIDTH-1:0] m_axis_scalar_45_tdata,
    input m_axis_scalar_45_tready,
    //output Scalar to AXI-Stream interface 46
    input m_axis_scalar_46_aclk,
    input m_axis_scalar_46_aresetn,
    output m_axis_scalar_46_tlast,
    output m_axis_scalar_46_tvalid,
    output [M_AXIS_SCALAR_46_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_46_tkeep,
    output [M_AXIS_SCALAR_46_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_46_tstrb,
    output [M_AXIS_SCALAR_46_DIRECT_DMWIDTH-1:0] m_axis_scalar_46_tdata,
    input m_axis_scalar_46_tready,
    //output Scalar to AXI-Stream interface 47
    input m_axis_scalar_47_aclk,
    input m_axis_scalar_47_aresetn,
    output m_axis_scalar_47_tlast,
    output m_axis_scalar_47_tvalid,
    output [M_AXIS_SCALAR_47_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_47_tkeep,
    output [M_AXIS_SCALAR_47_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_47_tstrb,
    output [M_AXIS_SCALAR_47_DIRECT_DMWIDTH-1:0] m_axis_scalar_47_tdata,
    input m_axis_scalar_47_tready,
    //output Scalar to AXI-Stream interface 48
    input m_axis_scalar_48_aclk,
    input m_axis_scalar_48_aresetn,
    output m_axis_scalar_48_tlast,
    output m_axis_scalar_48_tvalid,
    output [M_AXIS_SCALAR_48_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_48_tkeep,
    output [M_AXIS_SCALAR_48_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_48_tstrb,
    output [M_AXIS_SCALAR_48_DIRECT_DMWIDTH-1:0] m_axis_scalar_48_tdata,
    input m_axis_scalar_48_tready,
    //output Scalar to AXI-Stream interface 49
    input m_axis_scalar_49_aclk,
    input m_axis_scalar_49_aresetn,
    output m_axis_scalar_49_tlast,
    output m_axis_scalar_49_tvalid,
    output [M_AXIS_SCALAR_49_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_49_tkeep,
    output [M_AXIS_SCALAR_49_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_49_tstrb,
    output [M_AXIS_SCALAR_49_DIRECT_DMWIDTH-1:0] m_axis_scalar_49_tdata,
    input m_axis_scalar_49_tready,
    //output Scalar to AXI-Stream interface 50
    input m_axis_scalar_50_aclk,
    input m_axis_scalar_50_aresetn,
    output m_axis_scalar_50_tlast,
    output m_axis_scalar_50_tvalid,
    output [M_AXIS_SCALAR_50_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_50_tkeep,
    output [M_AXIS_SCALAR_50_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_50_tstrb,
    output [M_AXIS_SCALAR_50_DIRECT_DMWIDTH-1:0] m_axis_scalar_50_tdata,
    input m_axis_scalar_50_tready,
    //output Scalar to AXI-Stream interface 51
    input m_axis_scalar_51_aclk,
    input m_axis_scalar_51_aresetn,
    output m_axis_scalar_51_tlast,
    output m_axis_scalar_51_tvalid,
    output [M_AXIS_SCALAR_51_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_51_tkeep,
    output [M_AXIS_SCALAR_51_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_51_tstrb,
    output [M_AXIS_SCALAR_51_DIRECT_DMWIDTH-1:0] m_axis_scalar_51_tdata,
    input m_axis_scalar_51_tready,
    //output Scalar to AXI-Stream interface 52
    input m_axis_scalar_52_aclk,
    input m_axis_scalar_52_aresetn,
    output m_axis_scalar_52_tlast,
    output m_axis_scalar_52_tvalid,
    output [M_AXIS_SCALAR_52_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_52_tkeep,
    output [M_AXIS_SCALAR_52_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_52_tstrb,
    output [M_AXIS_SCALAR_52_DIRECT_DMWIDTH-1:0] m_axis_scalar_52_tdata,
    input m_axis_scalar_52_tready,
    //output Scalar to AXI-Stream interface 53
    input m_axis_scalar_53_aclk,
    input m_axis_scalar_53_aresetn,
    output m_axis_scalar_53_tlast,
    output m_axis_scalar_53_tvalid,
    output [M_AXIS_SCALAR_53_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_53_tkeep,
    output [M_AXIS_SCALAR_53_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_53_tstrb,
    output [M_AXIS_SCALAR_53_DIRECT_DMWIDTH-1:0] m_axis_scalar_53_tdata,
    input m_axis_scalar_53_tready,
    //output Scalar to AXI-Stream interface 54
    input m_axis_scalar_54_aclk,
    input m_axis_scalar_54_aresetn,
    output m_axis_scalar_54_tlast,
    output m_axis_scalar_54_tvalid,
    output [M_AXIS_SCALAR_54_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_54_tkeep,
    output [M_AXIS_SCALAR_54_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_54_tstrb,
    output [M_AXIS_SCALAR_54_DIRECT_DMWIDTH-1:0] m_axis_scalar_54_tdata,
    input m_axis_scalar_54_tready,
    //output Scalar to AXI-Stream interface 55
    input m_axis_scalar_55_aclk,
    input m_axis_scalar_55_aresetn,
    output m_axis_scalar_55_tlast,
    output m_axis_scalar_55_tvalid,
    output [M_AXIS_SCALAR_55_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_55_tkeep,
    output [M_AXIS_SCALAR_55_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_55_tstrb,
    output [M_AXIS_SCALAR_55_DIRECT_DMWIDTH-1:0] m_axis_scalar_55_tdata,
    input m_axis_scalar_55_tready,
    //output Scalar to AXI-Stream interface 56
    input m_axis_scalar_56_aclk,
    input m_axis_scalar_56_aresetn,
    output m_axis_scalar_56_tlast,
    output m_axis_scalar_56_tvalid,
    output [M_AXIS_SCALAR_56_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_56_tkeep,
    output [M_AXIS_SCALAR_56_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_56_tstrb,
    output [M_AXIS_SCALAR_56_DIRECT_DMWIDTH-1:0] m_axis_scalar_56_tdata,
    input m_axis_scalar_56_tready,
    //output Scalar to AXI-Stream interface 57
    input m_axis_scalar_57_aclk,
    input m_axis_scalar_57_aresetn,
    output m_axis_scalar_57_tlast,
    output m_axis_scalar_57_tvalid,
    output [M_AXIS_SCALAR_57_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_57_tkeep,
    output [M_AXIS_SCALAR_57_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_57_tstrb,
    output [M_AXIS_SCALAR_57_DIRECT_DMWIDTH-1:0] m_axis_scalar_57_tdata,
    input m_axis_scalar_57_tready,
    //output Scalar to AXI-Stream interface 58
    input m_axis_scalar_58_aclk,
    input m_axis_scalar_58_aresetn,
    output m_axis_scalar_58_tlast,
    output m_axis_scalar_58_tvalid,
    output [M_AXIS_SCALAR_58_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_58_tkeep,
    output [M_AXIS_SCALAR_58_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_58_tstrb,
    output [M_AXIS_SCALAR_58_DIRECT_DMWIDTH-1:0] m_axis_scalar_58_tdata,
    input m_axis_scalar_58_tready,
    //output Scalar to AXI-Stream interface 59
    input m_axis_scalar_59_aclk,
    input m_axis_scalar_59_aresetn,
    output m_axis_scalar_59_tlast,
    output m_axis_scalar_59_tvalid,
    output [M_AXIS_SCALAR_59_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_59_tkeep,
    output [M_AXIS_SCALAR_59_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_59_tstrb,
    output [M_AXIS_SCALAR_59_DIRECT_DMWIDTH-1:0] m_axis_scalar_59_tdata,
    input m_axis_scalar_59_tready,
    //output Scalar to AXI-Stream interface 60
    input m_axis_scalar_60_aclk,
    input m_axis_scalar_60_aresetn,
    output m_axis_scalar_60_tlast,
    output m_axis_scalar_60_tvalid,
    output [M_AXIS_SCALAR_60_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_60_tkeep,
    output [M_AXIS_SCALAR_60_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_60_tstrb,
    output [M_AXIS_SCALAR_60_DIRECT_DMWIDTH-1:0] m_axis_scalar_60_tdata,
    input m_axis_scalar_60_tready,
    //output Scalar to AXI-Stream interface 61
    input m_axis_scalar_61_aclk,
    input m_axis_scalar_61_aresetn,
    output m_axis_scalar_61_tlast,
    output m_axis_scalar_61_tvalid,
    output [M_AXIS_SCALAR_61_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_61_tkeep,
    output [M_AXIS_SCALAR_61_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_61_tstrb,
    output [M_AXIS_SCALAR_61_DIRECT_DMWIDTH-1:0] m_axis_scalar_61_tdata,
    input m_axis_scalar_61_tready,
    //output Scalar to AXI-Stream interface 62
    input m_axis_scalar_62_aclk,
    input m_axis_scalar_62_aresetn,
    output m_axis_scalar_62_tlast,
    output m_axis_scalar_62_tvalid,
    output [M_AXIS_SCALAR_62_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_62_tkeep,
    output [M_AXIS_SCALAR_62_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_62_tstrb,
    output [M_AXIS_SCALAR_62_DIRECT_DMWIDTH-1:0] m_axis_scalar_62_tdata,
    input m_axis_scalar_62_tready,
    //output Scalar to AXI-Stream interface 63
    input m_axis_scalar_63_aclk,
    input m_axis_scalar_63_aresetn,
    output m_axis_scalar_63_tlast,
    output m_axis_scalar_63_tvalid,
    output [M_AXIS_SCALAR_63_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_63_tkeep,
    output [M_AXIS_SCALAR_63_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_63_tstrb,
    output [M_AXIS_SCALAR_63_DIRECT_DMWIDTH-1:0] m_axis_scalar_63_tdata,
    input m_axis_scalar_63_tready,
    //output Scalar to AXI-Stream interface 64
    input m_axis_scalar_64_aclk,
    input m_axis_scalar_64_aresetn,
    output m_axis_scalar_64_tlast,
    output m_axis_scalar_64_tvalid,
    output [M_AXIS_SCALAR_64_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_64_tkeep,
    output [M_AXIS_SCALAR_64_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_64_tstrb,
    output [M_AXIS_SCALAR_64_DIRECT_DMWIDTH-1:0] m_axis_scalar_64_tdata,
    input m_axis_scalar_64_tready,
    //output Scalar to AXI-Stream interface 65
    input m_axis_scalar_65_aclk,
    input m_axis_scalar_65_aresetn,
    output m_axis_scalar_65_tlast,
    output m_axis_scalar_65_tvalid,
    output [M_AXIS_SCALAR_65_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_65_tkeep,
    output [M_AXIS_SCALAR_65_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_65_tstrb,
    output [M_AXIS_SCALAR_65_DIRECT_DMWIDTH-1:0] m_axis_scalar_65_tdata,
    input m_axis_scalar_65_tready,
    //output Scalar to AXI-Stream interface 66
    input m_axis_scalar_66_aclk,
    input m_axis_scalar_66_aresetn,
    output m_axis_scalar_66_tlast,
    output m_axis_scalar_66_tvalid,
    output [M_AXIS_SCALAR_66_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_66_tkeep,
    output [M_AXIS_SCALAR_66_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_66_tstrb,
    output [M_AXIS_SCALAR_66_DIRECT_DMWIDTH-1:0] m_axis_scalar_66_tdata,
    input m_axis_scalar_66_tready,
    //output Scalar to AXI-Stream interface 67
    input m_axis_scalar_67_aclk,
    input m_axis_scalar_67_aresetn,
    output m_axis_scalar_67_tlast,
    output m_axis_scalar_67_tvalid,
    output [M_AXIS_SCALAR_67_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_67_tkeep,
    output [M_AXIS_SCALAR_67_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_67_tstrb,
    output [M_AXIS_SCALAR_67_DIRECT_DMWIDTH-1:0] m_axis_scalar_67_tdata,
    input m_axis_scalar_67_tready,
    //output Scalar to AXI-Stream interface 68
    input m_axis_scalar_68_aclk,
    input m_axis_scalar_68_aresetn,
    output m_axis_scalar_68_tlast,
    output m_axis_scalar_68_tvalid,
    output [M_AXIS_SCALAR_68_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_68_tkeep,
    output [M_AXIS_SCALAR_68_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_68_tstrb,
    output [M_AXIS_SCALAR_68_DIRECT_DMWIDTH-1:0] m_axis_scalar_68_tdata,
    input m_axis_scalar_68_tready,
    //output Scalar to AXI-Stream interface 69
    input m_axis_scalar_69_aclk,
    input m_axis_scalar_69_aresetn,
    output m_axis_scalar_69_tlast,
    output m_axis_scalar_69_tvalid,
    output [M_AXIS_SCALAR_69_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_69_tkeep,
    output [M_AXIS_SCALAR_69_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_69_tstrb,
    output [M_AXIS_SCALAR_69_DIRECT_DMWIDTH-1:0] m_axis_scalar_69_tdata,
    input m_axis_scalar_69_tready,
    //output Scalar to AXI-Stream interface 70
    input m_axis_scalar_70_aclk,
    input m_axis_scalar_70_aresetn,
    output m_axis_scalar_70_tlast,
    output m_axis_scalar_70_tvalid,
    output [M_AXIS_SCALAR_70_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_70_tkeep,
    output [M_AXIS_SCALAR_70_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_70_tstrb,
    output [M_AXIS_SCALAR_70_DIRECT_DMWIDTH-1:0] m_axis_scalar_70_tdata,
    input m_axis_scalar_70_tready,
    //output Scalar to AXI-Stream interface 71
    input m_axis_scalar_71_aclk,
    input m_axis_scalar_71_aresetn,
    output m_axis_scalar_71_tlast,
    output m_axis_scalar_71_tvalid,
    output [M_AXIS_SCALAR_71_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_71_tkeep,
    output [M_AXIS_SCALAR_71_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_71_tstrb,
    output [M_AXIS_SCALAR_71_DIRECT_DMWIDTH-1:0] m_axis_scalar_71_tdata,
    input m_axis_scalar_71_tready,
    //output Scalar to AXI-Stream interface 72
    input m_axis_scalar_72_aclk,
    input m_axis_scalar_72_aresetn,
    output m_axis_scalar_72_tlast,
    output m_axis_scalar_72_tvalid,
    output [M_AXIS_SCALAR_72_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_72_tkeep,
    output [M_AXIS_SCALAR_72_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_72_tstrb,
    output [M_AXIS_SCALAR_72_DIRECT_DMWIDTH-1:0] m_axis_scalar_72_tdata,
    input m_axis_scalar_72_tready,
    //output Scalar to AXI-Stream interface 73
    input m_axis_scalar_73_aclk,
    input m_axis_scalar_73_aresetn,
    output m_axis_scalar_73_tlast,
    output m_axis_scalar_73_tvalid,
    output [M_AXIS_SCALAR_73_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_73_tkeep,
    output [M_AXIS_SCALAR_73_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_73_tstrb,
    output [M_AXIS_SCALAR_73_DIRECT_DMWIDTH-1:0] m_axis_scalar_73_tdata,
    input m_axis_scalar_73_tready,
    //output Scalar to AXI-Stream interface 74
    input m_axis_scalar_74_aclk,
    input m_axis_scalar_74_aresetn,
    output m_axis_scalar_74_tlast,
    output m_axis_scalar_74_tvalid,
    output [M_AXIS_SCALAR_74_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_74_tkeep,
    output [M_AXIS_SCALAR_74_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_74_tstrb,
    output [M_AXIS_SCALAR_74_DIRECT_DMWIDTH-1:0] m_axis_scalar_74_tdata,
    input m_axis_scalar_74_tready,
    //output Scalar to AXI-Stream interface 75
    input m_axis_scalar_75_aclk,
    input m_axis_scalar_75_aresetn,
    output m_axis_scalar_75_tlast,
    output m_axis_scalar_75_tvalid,
    output [M_AXIS_SCALAR_75_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_75_tkeep,
    output [M_AXIS_SCALAR_75_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_75_tstrb,
    output [M_AXIS_SCALAR_75_DIRECT_DMWIDTH-1:0] m_axis_scalar_75_tdata,
    input m_axis_scalar_75_tready,
    //output Scalar to AXI-Stream interface 76
    input m_axis_scalar_76_aclk,
    input m_axis_scalar_76_aresetn,
    output m_axis_scalar_76_tlast,
    output m_axis_scalar_76_tvalid,
    output [M_AXIS_SCALAR_76_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_76_tkeep,
    output [M_AXIS_SCALAR_76_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_76_tstrb,
    output [M_AXIS_SCALAR_76_DIRECT_DMWIDTH-1:0] m_axis_scalar_76_tdata,
    input m_axis_scalar_76_tready,
    //output Scalar to AXI-Stream interface 77
    input m_axis_scalar_77_aclk,
    input m_axis_scalar_77_aresetn,
    output m_axis_scalar_77_tlast,
    output m_axis_scalar_77_tvalid,
    output [M_AXIS_SCALAR_77_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_77_tkeep,
    output [M_AXIS_SCALAR_77_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_77_tstrb,
    output [M_AXIS_SCALAR_77_DIRECT_DMWIDTH-1:0] m_axis_scalar_77_tdata,
    input m_axis_scalar_77_tready,
    //output Scalar to AXI-Stream interface 78
    input m_axis_scalar_78_aclk,
    input m_axis_scalar_78_aresetn,
    output m_axis_scalar_78_tlast,
    output m_axis_scalar_78_tvalid,
    output [M_AXIS_SCALAR_78_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_78_tkeep,
    output [M_AXIS_SCALAR_78_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_78_tstrb,
    output [M_AXIS_SCALAR_78_DIRECT_DMWIDTH-1:0] m_axis_scalar_78_tdata,
    input m_axis_scalar_78_tready,
    //output Scalar to AXI-Stream interface 79
    input m_axis_scalar_79_aclk,
    input m_axis_scalar_79_aresetn,
    output m_axis_scalar_79_tlast,
    output m_axis_scalar_79_tvalid,
    output [M_AXIS_SCALAR_79_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_79_tkeep,
    output [M_AXIS_SCALAR_79_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_79_tstrb,
    output [M_AXIS_SCALAR_79_DIRECT_DMWIDTH-1:0] m_axis_scalar_79_tdata,
    input m_axis_scalar_79_tready,
    //output Scalar to AXI-Stream interface 80
    input m_axis_scalar_80_aclk,
    input m_axis_scalar_80_aresetn,
    output m_axis_scalar_80_tlast,
    output m_axis_scalar_80_tvalid,
    output [M_AXIS_SCALAR_80_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_80_tkeep,
    output [M_AXIS_SCALAR_80_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_80_tstrb,
    output [M_AXIS_SCALAR_80_DIRECT_DMWIDTH-1:0] m_axis_scalar_80_tdata,
    input m_axis_scalar_80_tready,
    //output Scalar to AXI-Stream interface 81
    input m_axis_scalar_81_aclk,
    input m_axis_scalar_81_aresetn,
    output m_axis_scalar_81_tlast,
    output m_axis_scalar_81_tvalid,
    output [M_AXIS_SCALAR_81_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_81_tkeep,
    output [M_AXIS_SCALAR_81_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_81_tstrb,
    output [M_AXIS_SCALAR_81_DIRECT_DMWIDTH-1:0] m_axis_scalar_81_tdata,
    input m_axis_scalar_81_tready,
    //output Scalar to AXI-Stream interface 82
    input m_axis_scalar_82_aclk,
    input m_axis_scalar_82_aresetn,
    output m_axis_scalar_82_tlast,
    output m_axis_scalar_82_tvalid,
    output [M_AXIS_SCALAR_82_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_82_tkeep,
    output [M_AXIS_SCALAR_82_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_82_tstrb,
    output [M_AXIS_SCALAR_82_DIRECT_DMWIDTH-1:0] m_axis_scalar_82_tdata,
    input m_axis_scalar_82_tready,
    //output Scalar to AXI-Stream interface 83
    input m_axis_scalar_83_aclk,
    input m_axis_scalar_83_aresetn,
    output m_axis_scalar_83_tlast,
    output m_axis_scalar_83_tvalid,
    output [M_AXIS_SCALAR_83_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_83_tkeep,
    output [M_AXIS_SCALAR_83_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_83_tstrb,
    output [M_AXIS_SCALAR_83_DIRECT_DMWIDTH-1:0] m_axis_scalar_83_tdata,
    input m_axis_scalar_83_tready,
    //output Scalar to AXI-Stream interface 84
    input m_axis_scalar_84_aclk,
    input m_axis_scalar_84_aresetn,
    output m_axis_scalar_84_tlast,
    output m_axis_scalar_84_tvalid,
    output [M_AXIS_SCALAR_84_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_84_tkeep,
    output [M_AXIS_SCALAR_84_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_84_tstrb,
    output [M_AXIS_SCALAR_84_DIRECT_DMWIDTH-1:0] m_axis_scalar_84_tdata,
    input m_axis_scalar_84_tready,
    //output Scalar to AXI-Stream interface 85
    input m_axis_scalar_85_aclk,
    input m_axis_scalar_85_aresetn,
    output m_axis_scalar_85_tlast,
    output m_axis_scalar_85_tvalid,
    output [M_AXIS_SCALAR_85_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_85_tkeep,
    output [M_AXIS_SCALAR_85_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_85_tstrb,
    output [M_AXIS_SCALAR_85_DIRECT_DMWIDTH-1:0] m_axis_scalar_85_tdata,
    input m_axis_scalar_85_tready,
    //output Scalar to AXI-Stream interface 86
    input m_axis_scalar_86_aclk,
    input m_axis_scalar_86_aresetn,
    output m_axis_scalar_86_tlast,
    output m_axis_scalar_86_tvalid,
    output [M_AXIS_SCALAR_86_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_86_tkeep,
    output [M_AXIS_SCALAR_86_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_86_tstrb,
    output [M_AXIS_SCALAR_86_DIRECT_DMWIDTH-1:0] m_axis_scalar_86_tdata,
    input m_axis_scalar_86_tready,
    //output Scalar to AXI-Stream interface 87
    input m_axis_scalar_87_aclk,
    input m_axis_scalar_87_aresetn,
    output m_axis_scalar_87_tlast,
    output m_axis_scalar_87_tvalid,
    output [M_AXIS_SCALAR_87_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_87_tkeep,
    output [M_AXIS_SCALAR_87_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_87_tstrb,
    output [M_AXIS_SCALAR_87_DIRECT_DMWIDTH-1:0] m_axis_scalar_87_tdata,
    input m_axis_scalar_87_tready,
    //output Scalar to AXI-Stream interface 88
    input m_axis_scalar_88_aclk,
    input m_axis_scalar_88_aresetn,
    output m_axis_scalar_88_tlast,
    output m_axis_scalar_88_tvalid,
    output [M_AXIS_SCALAR_88_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_88_tkeep,
    output [M_AXIS_SCALAR_88_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_88_tstrb,
    output [M_AXIS_SCALAR_88_DIRECT_DMWIDTH-1:0] m_axis_scalar_88_tdata,
    input m_axis_scalar_88_tready,
    //output Scalar to AXI-Stream interface 89
    input m_axis_scalar_89_aclk,
    input m_axis_scalar_89_aresetn,
    output m_axis_scalar_89_tlast,
    output m_axis_scalar_89_tvalid,
    output [M_AXIS_SCALAR_89_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_89_tkeep,
    output [M_AXIS_SCALAR_89_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_89_tstrb,
    output [M_AXIS_SCALAR_89_DIRECT_DMWIDTH-1:0] m_axis_scalar_89_tdata,
    input m_axis_scalar_89_tready,
    //output Scalar to AXI-Stream interface 90
    input m_axis_scalar_90_aclk,
    input m_axis_scalar_90_aresetn,
    output m_axis_scalar_90_tlast,
    output m_axis_scalar_90_tvalid,
    output [M_AXIS_SCALAR_90_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_90_tkeep,
    output [M_AXIS_SCALAR_90_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_90_tstrb,
    output [M_AXIS_SCALAR_90_DIRECT_DMWIDTH-1:0] m_axis_scalar_90_tdata,
    input m_axis_scalar_90_tready,
    //output Scalar to AXI-Stream interface 91
    input m_axis_scalar_91_aclk,
    input m_axis_scalar_91_aresetn,
    output m_axis_scalar_91_tlast,
    output m_axis_scalar_91_tvalid,
    output [M_AXIS_SCALAR_91_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_91_tkeep,
    output [M_AXIS_SCALAR_91_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_91_tstrb,
    output [M_AXIS_SCALAR_91_DIRECT_DMWIDTH-1:0] m_axis_scalar_91_tdata,
    input m_axis_scalar_91_tready,
    //output Scalar to AXI-Stream interface 92
    input m_axis_scalar_92_aclk,
    input m_axis_scalar_92_aresetn,
    output m_axis_scalar_92_tlast,
    output m_axis_scalar_92_tvalid,
    output [M_AXIS_SCALAR_92_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_92_tkeep,
    output [M_AXIS_SCALAR_92_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_92_tstrb,
    output [M_AXIS_SCALAR_92_DIRECT_DMWIDTH-1:0] m_axis_scalar_92_tdata,
    input m_axis_scalar_92_tready,
    //output Scalar to AXI-Stream interface 93
    input m_axis_scalar_93_aclk,
    input m_axis_scalar_93_aresetn,
    output m_axis_scalar_93_tlast,
    output m_axis_scalar_93_tvalid,
    output [M_AXIS_SCALAR_93_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_93_tkeep,
    output [M_AXIS_SCALAR_93_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_93_tstrb,
    output [M_AXIS_SCALAR_93_DIRECT_DMWIDTH-1:0] m_axis_scalar_93_tdata,
    input m_axis_scalar_93_tready,
    //output Scalar to AXI-Stream interface 94
    input m_axis_scalar_94_aclk,
    input m_axis_scalar_94_aresetn,
    output m_axis_scalar_94_tlast,
    output m_axis_scalar_94_tvalid,
    output [M_AXIS_SCALAR_94_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_94_tkeep,
    output [M_AXIS_SCALAR_94_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_94_tstrb,
    output [M_AXIS_SCALAR_94_DIRECT_DMWIDTH-1:0] m_axis_scalar_94_tdata,
    input m_axis_scalar_94_tready,
    //output Scalar to AXI-Stream interface 95
    input m_axis_scalar_95_aclk,
    input m_axis_scalar_95_aresetn,
    output m_axis_scalar_95_tlast,
    output m_axis_scalar_95_tvalid,
    output [M_AXIS_SCALAR_95_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_95_tkeep,
    output [M_AXIS_SCALAR_95_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_95_tstrb,
    output [M_AXIS_SCALAR_95_DIRECT_DMWIDTH-1:0] m_axis_scalar_95_tdata,
    input m_axis_scalar_95_tready,
    //output Scalar to AXI-Stream interface 96
    input m_axis_scalar_96_aclk,
    input m_axis_scalar_96_aresetn,
    output m_axis_scalar_96_tlast,
    output m_axis_scalar_96_tvalid,
    output [M_AXIS_SCALAR_96_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_96_tkeep,
    output [M_AXIS_SCALAR_96_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_96_tstrb,
    output [M_AXIS_SCALAR_96_DIRECT_DMWIDTH-1:0] m_axis_scalar_96_tdata,
    input m_axis_scalar_96_tready,
    //output Scalar to AXI-Stream interface 97
    input m_axis_scalar_97_aclk,
    input m_axis_scalar_97_aresetn,
    output m_axis_scalar_97_tlast,
    output m_axis_scalar_97_tvalid,
    output [M_AXIS_SCALAR_97_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_97_tkeep,
    output [M_AXIS_SCALAR_97_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_97_tstrb,
    output [M_AXIS_SCALAR_97_DIRECT_DMWIDTH-1:0] m_axis_scalar_97_tdata,
    input m_axis_scalar_97_tready,
    //output Scalar to AXI-Stream interface 98
    input m_axis_scalar_98_aclk,
    input m_axis_scalar_98_aresetn,
    output m_axis_scalar_98_tlast,
    output m_axis_scalar_98_tvalid,
    output [M_AXIS_SCALAR_98_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_98_tkeep,
    output [M_AXIS_SCALAR_98_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_98_tstrb,
    output [M_AXIS_SCALAR_98_DIRECT_DMWIDTH-1:0] m_axis_scalar_98_tdata,
    input m_axis_scalar_98_tready,
    //output Scalar to AXI-Stream interface 99
    input m_axis_scalar_99_aclk,
    input m_axis_scalar_99_aresetn,
    output m_axis_scalar_99_tlast,
    output m_axis_scalar_99_tvalid,
    output [M_AXIS_SCALAR_99_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_99_tkeep,
    output [M_AXIS_SCALAR_99_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_99_tstrb,
    output [M_AXIS_SCALAR_99_DIRECT_DMWIDTH-1:0] m_axis_scalar_99_tdata,
    input m_axis_scalar_99_tready,
    //output Scalar to AXI-Stream interface 100
    input m_axis_scalar_100_aclk,
    input m_axis_scalar_100_aresetn,
    output m_axis_scalar_100_tlast,
    output m_axis_scalar_100_tvalid,
    output [M_AXIS_SCALAR_100_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_100_tkeep,
    output [M_AXIS_SCALAR_100_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_100_tstrb,
    output [M_AXIS_SCALAR_100_DIRECT_DMWIDTH-1:0] m_axis_scalar_100_tdata,
    input m_axis_scalar_100_tready,
    //output Scalar to AXI-Stream interface 101
    input m_axis_scalar_101_aclk,
    input m_axis_scalar_101_aresetn,
    output m_axis_scalar_101_tlast,
    output m_axis_scalar_101_tvalid,
    output [M_AXIS_SCALAR_101_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_101_tkeep,
    output [M_AXIS_SCALAR_101_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_101_tstrb,
    output [M_AXIS_SCALAR_101_DIRECT_DMWIDTH-1:0] m_axis_scalar_101_tdata,
    input m_axis_scalar_101_tready,
    //output Scalar to AXI-Stream interface 102
    input m_axis_scalar_102_aclk,
    input m_axis_scalar_102_aresetn,
    output m_axis_scalar_102_tlast,
    output m_axis_scalar_102_tvalid,
    output [M_AXIS_SCALAR_102_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_102_tkeep,
    output [M_AXIS_SCALAR_102_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_102_tstrb,
    output [M_AXIS_SCALAR_102_DIRECT_DMWIDTH-1:0] m_axis_scalar_102_tdata,
    input m_axis_scalar_102_tready,
    //output Scalar to AXI-Stream interface 103
    input m_axis_scalar_103_aclk,
    input m_axis_scalar_103_aresetn,
    output m_axis_scalar_103_tlast,
    output m_axis_scalar_103_tvalid,
    output [M_AXIS_SCALAR_103_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_103_tkeep,
    output [M_AXIS_SCALAR_103_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_103_tstrb,
    output [M_AXIS_SCALAR_103_DIRECT_DMWIDTH-1:0] m_axis_scalar_103_tdata,
    input m_axis_scalar_103_tready,
    //output Scalar to AXI-Stream interface 104
    input m_axis_scalar_104_aclk,
    input m_axis_scalar_104_aresetn,
    output m_axis_scalar_104_tlast,
    output m_axis_scalar_104_tvalid,
    output [M_AXIS_SCALAR_104_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_104_tkeep,
    output [M_AXIS_SCALAR_104_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_104_tstrb,
    output [M_AXIS_SCALAR_104_DIRECT_DMWIDTH-1:0] m_axis_scalar_104_tdata,
    input m_axis_scalar_104_tready,
    //output Scalar to AXI-Stream interface 105
    input m_axis_scalar_105_aclk,
    input m_axis_scalar_105_aresetn,
    output m_axis_scalar_105_tlast,
    output m_axis_scalar_105_tvalid,
    output [M_AXIS_SCALAR_105_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_105_tkeep,
    output [M_AXIS_SCALAR_105_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_105_tstrb,
    output [M_AXIS_SCALAR_105_DIRECT_DMWIDTH-1:0] m_axis_scalar_105_tdata,
    input m_axis_scalar_105_tready,
    //output Scalar to AXI-Stream interface 106
    input m_axis_scalar_106_aclk,
    input m_axis_scalar_106_aresetn,
    output m_axis_scalar_106_tlast,
    output m_axis_scalar_106_tvalid,
    output [M_AXIS_SCALAR_106_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_106_tkeep,
    output [M_AXIS_SCALAR_106_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_106_tstrb,
    output [M_AXIS_SCALAR_106_DIRECT_DMWIDTH-1:0] m_axis_scalar_106_tdata,
    input m_axis_scalar_106_tready,
    //output Scalar to AXI-Stream interface 107
    input m_axis_scalar_107_aclk,
    input m_axis_scalar_107_aresetn,
    output m_axis_scalar_107_tlast,
    output m_axis_scalar_107_tvalid,
    output [M_AXIS_SCALAR_107_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_107_tkeep,
    output [M_AXIS_SCALAR_107_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_107_tstrb,
    output [M_AXIS_SCALAR_107_DIRECT_DMWIDTH-1:0] m_axis_scalar_107_tdata,
    input m_axis_scalar_107_tready,
    //output Scalar to AXI-Stream interface 108
    input m_axis_scalar_108_aclk,
    input m_axis_scalar_108_aresetn,
    output m_axis_scalar_108_tlast,
    output m_axis_scalar_108_tvalid,
    output [M_AXIS_SCALAR_108_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_108_tkeep,
    output [M_AXIS_SCALAR_108_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_108_tstrb,
    output [M_AXIS_SCALAR_108_DIRECT_DMWIDTH-1:0] m_axis_scalar_108_tdata,
    input m_axis_scalar_108_tready,
    //output Scalar to AXI-Stream interface 109
    input m_axis_scalar_109_aclk,
    input m_axis_scalar_109_aresetn,
    output m_axis_scalar_109_tlast,
    output m_axis_scalar_109_tvalid,
    output [M_AXIS_SCALAR_109_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_109_tkeep,
    output [M_AXIS_SCALAR_109_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_109_tstrb,
    output [M_AXIS_SCALAR_109_DIRECT_DMWIDTH-1:0] m_axis_scalar_109_tdata,
    input m_axis_scalar_109_tready,
    //output Scalar to AXI-Stream interface 110
    input m_axis_scalar_110_aclk,
    input m_axis_scalar_110_aresetn,
    output m_axis_scalar_110_tlast,
    output m_axis_scalar_110_tvalid,
    output [M_AXIS_SCALAR_110_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_110_tkeep,
    output [M_AXIS_SCALAR_110_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_110_tstrb,
    output [M_AXIS_SCALAR_110_DIRECT_DMWIDTH-1:0] m_axis_scalar_110_tdata,
    input m_axis_scalar_110_tready,
    //output Scalar to AXI-Stream interface 111
    input m_axis_scalar_111_aclk,
    input m_axis_scalar_111_aresetn,
    output m_axis_scalar_111_tlast,
    output m_axis_scalar_111_tvalid,
    output [M_AXIS_SCALAR_111_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_111_tkeep,
    output [M_AXIS_SCALAR_111_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_111_tstrb,
    output [M_AXIS_SCALAR_111_DIRECT_DMWIDTH-1:0] m_axis_scalar_111_tdata,
    input m_axis_scalar_111_tready,
    //output Scalar to AXI-Stream interface 112
    input m_axis_scalar_112_aclk,
    input m_axis_scalar_112_aresetn,
    output m_axis_scalar_112_tlast,
    output m_axis_scalar_112_tvalid,
    output [M_AXIS_SCALAR_112_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_112_tkeep,
    output [M_AXIS_SCALAR_112_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_112_tstrb,
    output [M_AXIS_SCALAR_112_DIRECT_DMWIDTH-1:0] m_axis_scalar_112_tdata,
    input m_axis_scalar_112_tready,
    //output Scalar to AXI-Stream interface 113
    input m_axis_scalar_113_aclk,
    input m_axis_scalar_113_aresetn,
    output m_axis_scalar_113_tlast,
    output m_axis_scalar_113_tvalid,
    output [M_AXIS_SCALAR_113_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_113_tkeep,
    output [M_AXIS_SCALAR_113_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_113_tstrb,
    output [M_AXIS_SCALAR_113_DIRECT_DMWIDTH-1:0] m_axis_scalar_113_tdata,
    input m_axis_scalar_113_tready,
    //output Scalar to AXI-Stream interface 114
    input m_axis_scalar_114_aclk,
    input m_axis_scalar_114_aresetn,
    output m_axis_scalar_114_tlast,
    output m_axis_scalar_114_tvalid,
    output [M_AXIS_SCALAR_114_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_114_tkeep,
    output [M_AXIS_SCALAR_114_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_114_tstrb,
    output [M_AXIS_SCALAR_114_DIRECT_DMWIDTH-1:0] m_axis_scalar_114_tdata,
    input m_axis_scalar_114_tready,
    //output Scalar to AXI-Stream interface 115
    input m_axis_scalar_115_aclk,
    input m_axis_scalar_115_aresetn,
    output m_axis_scalar_115_tlast,
    output m_axis_scalar_115_tvalid,
    output [M_AXIS_SCALAR_115_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_115_tkeep,
    output [M_AXIS_SCALAR_115_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_115_tstrb,
    output [M_AXIS_SCALAR_115_DIRECT_DMWIDTH-1:0] m_axis_scalar_115_tdata,
    input m_axis_scalar_115_tready,
    //output Scalar to AXI-Stream interface 116
    input m_axis_scalar_116_aclk,
    input m_axis_scalar_116_aresetn,
    output m_axis_scalar_116_tlast,
    output m_axis_scalar_116_tvalid,
    output [M_AXIS_SCALAR_116_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_116_tkeep,
    output [M_AXIS_SCALAR_116_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_116_tstrb,
    output [M_AXIS_SCALAR_116_DIRECT_DMWIDTH-1:0] m_axis_scalar_116_tdata,
    input m_axis_scalar_116_tready,
    //output Scalar to AXI-Stream interface 117
    input m_axis_scalar_117_aclk,
    input m_axis_scalar_117_aresetn,
    output m_axis_scalar_117_tlast,
    output m_axis_scalar_117_tvalid,
    output [M_AXIS_SCALAR_117_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_117_tkeep,
    output [M_AXIS_SCALAR_117_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_117_tstrb,
    output [M_AXIS_SCALAR_117_DIRECT_DMWIDTH-1:0] m_axis_scalar_117_tdata,
    input m_axis_scalar_117_tready,
    //output Scalar to AXI-Stream interface 118
    input m_axis_scalar_118_aclk,
    input m_axis_scalar_118_aresetn,
    output m_axis_scalar_118_tlast,
    output m_axis_scalar_118_tvalid,
    output [M_AXIS_SCALAR_118_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_118_tkeep,
    output [M_AXIS_SCALAR_118_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_118_tstrb,
    output [M_AXIS_SCALAR_118_DIRECT_DMWIDTH-1:0] m_axis_scalar_118_tdata,
    input m_axis_scalar_118_tready,
    //output Scalar to AXI-Stream interface 119
    input m_axis_scalar_119_aclk,
    input m_axis_scalar_119_aresetn,
    output m_axis_scalar_119_tlast,
    output m_axis_scalar_119_tvalid,
    output [M_AXIS_SCALAR_119_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_119_tkeep,
    output [M_AXIS_SCALAR_119_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_119_tstrb,
    output [M_AXIS_SCALAR_119_DIRECT_DMWIDTH-1:0] m_axis_scalar_119_tdata,
    input m_axis_scalar_119_tready,
    //output Scalar to AXI-Stream interface 120
    input m_axis_scalar_120_aclk,
    input m_axis_scalar_120_aresetn,
    output m_axis_scalar_120_tlast,
    output m_axis_scalar_120_tvalid,
    output [M_AXIS_SCALAR_120_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_120_tkeep,
    output [M_AXIS_SCALAR_120_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_120_tstrb,
    output [M_AXIS_SCALAR_120_DIRECT_DMWIDTH-1:0] m_axis_scalar_120_tdata,
    input m_axis_scalar_120_tready,
    //output Scalar to AXI-Stream interface 121
    input m_axis_scalar_121_aclk,
    input m_axis_scalar_121_aresetn,
    output m_axis_scalar_121_tlast,
    output m_axis_scalar_121_tvalid,
    output [M_AXIS_SCALAR_121_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_121_tkeep,
    output [M_AXIS_SCALAR_121_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_121_tstrb,
    output [M_AXIS_SCALAR_121_DIRECT_DMWIDTH-1:0] m_axis_scalar_121_tdata,
    input m_axis_scalar_121_tready,
    //output Scalar to AXI-Stream interface 122
    input m_axis_scalar_122_aclk,
    input m_axis_scalar_122_aresetn,
    output m_axis_scalar_122_tlast,
    output m_axis_scalar_122_tvalid,
    output [M_AXIS_SCALAR_122_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_122_tkeep,
    output [M_AXIS_SCALAR_122_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_122_tstrb,
    output [M_AXIS_SCALAR_122_DIRECT_DMWIDTH-1:0] m_axis_scalar_122_tdata,
    input m_axis_scalar_122_tready,
    //output Scalar to AXI-Stream interface 123
    input m_axis_scalar_123_aclk,
    input m_axis_scalar_123_aresetn,
    output m_axis_scalar_123_tlast,
    output m_axis_scalar_123_tvalid,
    output [M_AXIS_SCALAR_123_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_123_tkeep,
    output [M_AXIS_SCALAR_123_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_123_tstrb,
    output [M_AXIS_SCALAR_123_DIRECT_DMWIDTH-1:0] m_axis_scalar_123_tdata,
    input m_axis_scalar_123_tready,
    //output Scalar to AXI-Stream interface 124
    input m_axis_scalar_124_aclk,
    input m_axis_scalar_124_aresetn,
    output m_axis_scalar_124_tlast,
    output m_axis_scalar_124_tvalid,
    output [M_AXIS_SCALAR_124_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_124_tkeep,
    output [M_AXIS_SCALAR_124_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_124_tstrb,
    output [M_AXIS_SCALAR_124_DIRECT_DMWIDTH-1:0] m_axis_scalar_124_tdata,
    input m_axis_scalar_124_tready,
    //output Scalar to AXI-Stream interface 125
    input m_axis_scalar_125_aclk,
    input m_axis_scalar_125_aresetn,
    output m_axis_scalar_125_tlast,
    output m_axis_scalar_125_tvalid,
    output [M_AXIS_SCALAR_125_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_125_tkeep,
    output [M_AXIS_SCALAR_125_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_125_tstrb,
    output [M_AXIS_SCALAR_125_DIRECT_DMWIDTH-1:0] m_axis_scalar_125_tdata,
    input m_axis_scalar_125_tready,
    //output Scalar to AXI-Stream interface 126
    input m_axis_scalar_126_aclk,
    input m_axis_scalar_126_aresetn,
    output m_axis_scalar_126_tlast,
    output m_axis_scalar_126_tvalid,
    output [M_AXIS_SCALAR_126_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_126_tkeep,
    output [M_AXIS_SCALAR_126_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_126_tstrb,
    output [M_AXIS_SCALAR_126_DIRECT_DMWIDTH-1:0] m_axis_scalar_126_tdata,
    input m_axis_scalar_126_tready,
    //output Scalar to AXI-Stream interface 127
    input m_axis_scalar_127_aclk,
    input m_axis_scalar_127_aresetn,
    output m_axis_scalar_127_tlast,
    output m_axis_scalar_127_tvalid,
    output [M_AXIS_SCALAR_127_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_127_tkeep,
    output [M_AXIS_SCALAR_127_DIRECT_DMWIDTH/8-1:0] m_axis_scalar_127_tstrb,
    output [M_AXIS_SCALAR_127_DIRECT_DMWIDTH-1:0] m_axis_scalar_127_tdata,
    input m_axis_scalar_127_tready,
    //-----------------------------------------------------
    //input AXI-Stream to FIFO interface 0
    input s_axis_fifo_0_aclk,
    input s_axis_fifo_0_aresetn,
    input s_axis_fifo_0_tlast,
    input s_axis_fifo_0_tvalid,
    input [S_AXIS_FIFO_0_DMWIDTH/8-1:0] s_axis_fifo_0_tkeep,
    input [S_AXIS_FIFO_0_DMWIDTH/8-1:0] s_axis_fifo_0_tstrb,
    input [S_AXIS_FIFO_0_DMWIDTH-1:0] s_axis_fifo_0_tdata,
    output s_axis_fifo_0_tready,
    output ap_fifo_iarg_0_empty_n,
    output [S_AXIS_FIFO_0_WIDTH-1:0] ap_fifo_iarg_0_dout,
    input ap_fifo_iarg_0_read,
    //input AXI-Stream to FIFO interface 1
    input s_axis_fifo_1_aclk,
    input s_axis_fifo_1_aresetn,
    input s_axis_fifo_1_tlast,
    input s_axis_fifo_1_tvalid,
    input [S_AXIS_FIFO_1_DMWIDTH/8-1:0] s_axis_fifo_1_tkeep,
    input [S_AXIS_FIFO_1_DMWIDTH/8-1:0] s_axis_fifo_1_tstrb,
    input [S_AXIS_FIFO_1_DMWIDTH-1:0] s_axis_fifo_1_tdata,
    output s_axis_fifo_1_tready,
    output ap_fifo_iarg_1_empty_n,
    output [S_AXIS_FIFO_1_WIDTH-1:0] ap_fifo_iarg_1_dout,
    input ap_fifo_iarg_1_read,
    //input AXI-Stream to FIFO interface 2
    input s_axis_fifo_2_aclk,
    input s_axis_fifo_2_aresetn,
    input s_axis_fifo_2_tlast,
    input s_axis_fifo_2_tvalid,
    input [S_AXIS_FIFO_2_DMWIDTH/8-1:0] s_axis_fifo_2_tkeep,
    input [S_AXIS_FIFO_2_DMWIDTH/8-1:0] s_axis_fifo_2_tstrb,
    input [S_AXIS_FIFO_2_DMWIDTH-1:0] s_axis_fifo_2_tdata,
    output s_axis_fifo_2_tready,
    output ap_fifo_iarg_2_empty_n,
    output [S_AXIS_FIFO_2_WIDTH-1:0] ap_fifo_iarg_2_dout,
    input ap_fifo_iarg_2_read,
    //input AXI-Stream to FIFO interface 3
    input s_axis_fifo_3_aclk,
    input s_axis_fifo_3_aresetn,
    input s_axis_fifo_3_tlast,
    input s_axis_fifo_3_tvalid,
    input [S_AXIS_FIFO_3_DMWIDTH/8-1:0] s_axis_fifo_3_tkeep,
    input [S_AXIS_FIFO_3_DMWIDTH/8-1:0] s_axis_fifo_3_tstrb,
    input [S_AXIS_FIFO_3_DMWIDTH-1:0] s_axis_fifo_3_tdata,
    output s_axis_fifo_3_tready,
    output ap_fifo_iarg_3_empty_n,
    output [S_AXIS_FIFO_3_WIDTH-1:0] ap_fifo_iarg_3_dout,
    input ap_fifo_iarg_3_read,
    //input AXI-Stream to FIFO interface 4
    input s_axis_fifo_4_aclk,
    input s_axis_fifo_4_aresetn,
    input s_axis_fifo_4_tlast,
    input s_axis_fifo_4_tvalid,
    input [S_AXIS_FIFO_4_DMWIDTH/8-1:0] s_axis_fifo_4_tkeep,
    input [S_AXIS_FIFO_4_DMWIDTH/8-1:0] s_axis_fifo_4_tstrb,
    input [S_AXIS_FIFO_4_DMWIDTH-1:0] s_axis_fifo_4_tdata,
    output s_axis_fifo_4_tready,
    output ap_fifo_iarg_4_empty_n,
    output [S_AXIS_FIFO_4_WIDTH-1:0] ap_fifo_iarg_4_dout,
    input ap_fifo_iarg_4_read,
    //input AXI-Stream to FIFO interface 5
    input s_axis_fifo_5_aclk,
    input s_axis_fifo_5_aresetn,
    input s_axis_fifo_5_tlast,
    input s_axis_fifo_5_tvalid,
    input [S_AXIS_FIFO_5_DMWIDTH/8-1:0] s_axis_fifo_5_tkeep,
    input [S_AXIS_FIFO_5_DMWIDTH/8-1:0] s_axis_fifo_5_tstrb,
    input [S_AXIS_FIFO_5_DMWIDTH-1:0] s_axis_fifo_5_tdata,
    output s_axis_fifo_5_tready,
    output ap_fifo_iarg_5_empty_n,
    output [S_AXIS_FIFO_5_WIDTH-1:0] ap_fifo_iarg_5_dout,
    input ap_fifo_iarg_5_read,
    //input AXI-Stream to FIFO interface 6
    input s_axis_fifo_6_aclk,
    input s_axis_fifo_6_aresetn,
    input s_axis_fifo_6_tlast,
    input s_axis_fifo_6_tvalid,
    input [S_AXIS_FIFO_6_DMWIDTH/8-1:0] s_axis_fifo_6_tkeep,
    input [S_AXIS_FIFO_6_DMWIDTH/8-1:0] s_axis_fifo_6_tstrb,
    input [S_AXIS_FIFO_6_DMWIDTH-1:0] s_axis_fifo_6_tdata,
    output s_axis_fifo_6_tready,
    output ap_fifo_iarg_6_empty_n,
    output [S_AXIS_FIFO_6_WIDTH-1:0] ap_fifo_iarg_6_dout,
    input ap_fifo_iarg_6_read,
    //input AXI-Stream to FIFO interface 7
    input s_axis_fifo_7_aclk,
    input s_axis_fifo_7_aresetn,
    input s_axis_fifo_7_tlast,
    input s_axis_fifo_7_tvalid,
    input [S_AXIS_FIFO_7_DMWIDTH/8-1:0] s_axis_fifo_7_tkeep,
    input [S_AXIS_FIFO_7_DMWIDTH/8-1:0] s_axis_fifo_7_tstrb,
    input [S_AXIS_FIFO_7_DMWIDTH-1:0] s_axis_fifo_7_tdata,
    output s_axis_fifo_7_tready,
    output ap_fifo_iarg_7_empty_n,
    output [S_AXIS_FIFO_7_WIDTH-1:0] ap_fifo_iarg_7_dout,
    input ap_fifo_iarg_7_read,
    //input AXI-Stream to FIFO interface 8
    input s_axis_fifo_8_aclk,
    input s_axis_fifo_8_aresetn,
    input s_axis_fifo_8_tlast,
    input s_axis_fifo_8_tvalid,
    input [S_AXIS_FIFO_8_DMWIDTH/8-1:0] s_axis_fifo_8_tkeep,
    input [S_AXIS_FIFO_8_DMWIDTH/8-1:0] s_axis_fifo_8_tstrb,
    input [S_AXIS_FIFO_8_DMWIDTH-1:0] s_axis_fifo_8_tdata,
    output s_axis_fifo_8_tready,
    output ap_fifo_iarg_8_empty_n,
    output [S_AXIS_FIFO_8_WIDTH-1:0] ap_fifo_iarg_8_dout,
    input ap_fifo_iarg_8_read,
    //input AXI-Stream to FIFO interface 9
    input s_axis_fifo_9_aclk,
    input s_axis_fifo_9_aresetn,
    input s_axis_fifo_9_tlast,
    input s_axis_fifo_9_tvalid,
    input [S_AXIS_FIFO_9_DMWIDTH/8-1:0] s_axis_fifo_9_tkeep,
    input [S_AXIS_FIFO_9_DMWIDTH/8-1:0] s_axis_fifo_9_tstrb,
    input [S_AXIS_FIFO_9_DMWIDTH-1:0] s_axis_fifo_9_tdata,
    output s_axis_fifo_9_tready,
    output ap_fifo_iarg_9_empty_n,
    output [S_AXIS_FIFO_9_WIDTH-1:0] ap_fifo_iarg_9_dout,
    input ap_fifo_iarg_9_read,
    //input AXI-Stream to FIFO interface 10
    input s_axis_fifo_10_aclk,
    input s_axis_fifo_10_aresetn,
    input s_axis_fifo_10_tlast,
    input s_axis_fifo_10_tvalid,
    input [S_AXIS_FIFO_10_DMWIDTH/8-1:0] s_axis_fifo_10_tkeep,
    input [S_AXIS_FIFO_10_DMWIDTH/8-1:0] s_axis_fifo_10_tstrb,
    input [S_AXIS_FIFO_10_DMWIDTH-1:0] s_axis_fifo_10_tdata,
    output s_axis_fifo_10_tready,
    output ap_fifo_iarg_10_empty_n,
    output [S_AXIS_FIFO_10_WIDTH-1:0] ap_fifo_iarg_10_dout,
    input ap_fifo_iarg_10_read,
    //input AXI-Stream to FIFO interface 11
    input s_axis_fifo_11_aclk,
    input s_axis_fifo_11_aresetn,
    input s_axis_fifo_11_tlast,
    input s_axis_fifo_11_tvalid,
    input [S_AXIS_FIFO_11_DMWIDTH/8-1:0] s_axis_fifo_11_tkeep,
    input [S_AXIS_FIFO_11_DMWIDTH/8-1:0] s_axis_fifo_11_tstrb,
    input [S_AXIS_FIFO_11_DMWIDTH-1:0] s_axis_fifo_11_tdata,
    output s_axis_fifo_11_tready,
    output ap_fifo_iarg_11_empty_n,
    output [S_AXIS_FIFO_11_WIDTH-1:0] ap_fifo_iarg_11_dout,
    input ap_fifo_iarg_11_read,
    //input AXI-Stream to FIFO interface 12
    input s_axis_fifo_12_aclk,
    input s_axis_fifo_12_aresetn,
    input s_axis_fifo_12_tlast,
    input s_axis_fifo_12_tvalid,
    input [S_AXIS_FIFO_12_DMWIDTH/8-1:0] s_axis_fifo_12_tkeep,
    input [S_AXIS_FIFO_12_DMWIDTH/8-1:0] s_axis_fifo_12_tstrb,
    input [S_AXIS_FIFO_12_DMWIDTH-1:0] s_axis_fifo_12_tdata,
    output s_axis_fifo_12_tready,
    output ap_fifo_iarg_12_empty_n,
    output [S_AXIS_FIFO_12_WIDTH-1:0] ap_fifo_iarg_12_dout,
    input ap_fifo_iarg_12_read,
    //input AXI-Stream to FIFO interface 13
    input s_axis_fifo_13_aclk,
    input s_axis_fifo_13_aresetn,
    input s_axis_fifo_13_tlast,
    input s_axis_fifo_13_tvalid,
    input [S_AXIS_FIFO_13_DMWIDTH/8-1:0] s_axis_fifo_13_tkeep,
    input [S_AXIS_FIFO_13_DMWIDTH/8-1:0] s_axis_fifo_13_tstrb,
    input [S_AXIS_FIFO_13_DMWIDTH-1:0] s_axis_fifo_13_tdata,
    output s_axis_fifo_13_tready,
    output ap_fifo_iarg_13_empty_n,
    output [S_AXIS_FIFO_13_WIDTH-1:0] ap_fifo_iarg_13_dout,
    input ap_fifo_iarg_13_read,
    //input AXI-Stream to FIFO interface 14
    input s_axis_fifo_14_aclk,
    input s_axis_fifo_14_aresetn,
    input s_axis_fifo_14_tlast,
    input s_axis_fifo_14_tvalid,
    input [S_AXIS_FIFO_14_DMWIDTH/8-1:0] s_axis_fifo_14_tkeep,
    input [S_AXIS_FIFO_14_DMWIDTH/8-1:0] s_axis_fifo_14_tstrb,
    input [S_AXIS_FIFO_14_DMWIDTH-1:0] s_axis_fifo_14_tdata,
    output s_axis_fifo_14_tready,
    output ap_fifo_iarg_14_empty_n,
    output [S_AXIS_FIFO_14_WIDTH-1:0] ap_fifo_iarg_14_dout,
    input ap_fifo_iarg_14_read,
    //input AXI-Stream to FIFO interface 15
    input s_axis_fifo_15_aclk,
    input s_axis_fifo_15_aresetn,
    input s_axis_fifo_15_tlast,
    input s_axis_fifo_15_tvalid,
    input [S_AXIS_FIFO_15_DMWIDTH/8-1:0] s_axis_fifo_15_tkeep,
    input [S_AXIS_FIFO_15_DMWIDTH/8-1:0] s_axis_fifo_15_tstrb,
    input [S_AXIS_FIFO_15_DMWIDTH-1:0] s_axis_fifo_15_tdata,
    output s_axis_fifo_15_tready,
    output ap_fifo_iarg_15_empty_n,
    output [S_AXIS_FIFO_15_WIDTH-1:0] ap_fifo_iarg_15_dout,
    input ap_fifo_iarg_15_read,
    //input AXI-Stream to FIFO interface 16
    input s_axis_fifo_16_aclk,
    input s_axis_fifo_16_aresetn,
    input s_axis_fifo_16_tlast,
    input s_axis_fifo_16_tvalid,
    input [S_AXIS_FIFO_16_DMWIDTH/8-1:0] s_axis_fifo_16_tkeep,
    input [S_AXIS_FIFO_16_DMWIDTH/8-1:0] s_axis_fifo_16_tstrb,
    input [S_AXIS_FIFO_16_DMWIDTH-1:0] s_axis_fifo_16_tdata,
    output s_axis_fifo_16_tready,
    output ap_fifo_iarg_16_empty_n,
    output [S_AXIS_FIFO_16_WIDTH-1:0] ap_fifo_iarg_16_dout,
    input ap_fifo_iarg_16_read,
    //input AXI-Stream to FIFO interface 17
    input s_axis_fifo_17_aclk,
    input s_axis_fifo_17_aresetn,
    input s_axis_fifo_17_tlast,
    input s_axis_fifo_17_tvalid,
    input [S_AXIS_FIFO_17_DMWIDTH/8-1:0] s_axis_fifo_17_tkeep,
    input [S_AXIS_FIFO_17_DMWIDTH/8-1:0] s_axis_fifo_17_tstrb,
    input [S_AXIS_FIFO_17_DMWIDTH-1:0] s_axis_fifo_17_tdata,
    output s_axis_fifo_17_tready,
    output ap_fifo_iarg_17_empty_n,
    output [S_AXIS_FIFO_17_WIDTH-1:0] ap_fifo_iarg_17_dout,
    input ap_fifo_iarg_17_read,
    //input AXI-Stream to FIFO interface 18
    input s_axis_fifo_18_aclk,
    input s_axis_fifo_18_aresetn,
    input s_axis_fifo_18_tlast,
    input s_axis_fifo_18_tvalid,
    input [S_AXIS_FIFO_18_DMWIDTH/8-1:0] s_axis_fifo_18_tkeep,
    input [S_AXIS_FIFO_18_DMWIDTH/8-1:0] s_axis_fifo_18_tstrb,
    input [S_AXIS_FIFO_18_DMWIDTH-1:0] s_axis_fifo_18_tdata,
    output s_axis_fifo_18_tready,
    output ap_fifo_iarg_18_empty_n,
    output [S_AXIS_FIFO_18_WIDTH-1:0] ap_fifo_iarg_18_dout,
    input ap_fifo_iarg_18_read,
    //input AXI-Stream to FIFO interface 19
    input s_axis_fifo_19_aclk,
    input s_axis_fifo_19_aresetn,
    input s_axis_fifo_19_tlast,
    input s_axis_fifo_19_tvalid,
    input [S_AXIS_FIFO_19_DMWIDTH/8-1:0] s_axis_fifo_19_tkeep,
    input [S_AXIS_FIFO_19_DMWIDTH/8-1:0] s_axis_fifo_19_tstrb,
    input [S_AXIS_FIFO_19_DMWIDTH-1:0] s_axis_fifo_19_tdata,
    output s_axis_fifo_19_tready,
    output ap_fifo_iarg_19_empty_n,
    output [S_AXIS_FIFO_19_WIDTH-1:0] ap_fifo_iarg_19_dout,
    input ap_fifo_iarg_19_read,
    //input AXI-Stream to FIFO interface 20
    input s_axis_fifo_20_aclk,
    input s_axis_fifo_20_aresetn,
    input s_axis_fifo_20_tlast,
    input s_axis_fifo_20_tvalid,
    input [S_AXIS_FIFO_20_DMWIDTH/8-1:0] s_axis_fifo_20_tkeep,
    input [S_AXIS_FIFO_20_DMWIDTH/8-1:0] s_axis_fifo_20_tstrb,
    input [S_AXIS_FIFO_20_DMWIDTH-1:0] s_axis_fifo_20_tdata,
    output s_axis_fifo_20_tready,
    output ap_fifo_iarg_20_empty_n,
    output [S_AXIS_FIFO_20_WIDTH-1:0] ap_fifo_iarg_20_dout,
    input ap_fifo_iarg_20_read,
    //input AXI-Stream to FIFO interface 21
    input s_axis_fifo_21_aclk,
    input s_axis_fifo_21_aresetn,
    input s_axis_fifo_21_tlast,
    input s_axis_fifo_21_tvalid,
    input [S_AXIS_FIFO_21_DMWIDTH/8-1:0] s_axis_fifo_21_tkeep,
    input [S_AXIS_FIFO_21_DMWIDTH/8-1:0] s_axis_fifo_21_tstrb,
    input [S_AXIS_FIFO_21_DMWIDTH-1:0] s_axis_fifo_21_tdata,
    output s_axis_fifo_21_tready,
    output ap_fifo_iarg_21_empty_n,
    output [S_AXIS_FIFO_21_WIDTH-1:0] ap_fifo_iarg_21_dout,
    input ap_fifo_iarg_21_read,
    //input AXI-Stream to FIFO interface 22
    input s_axis_fifo_22_aclk,
    input s_axis_fifo_22_aresetn,
    input s_axis_fifo_22_tlast,
    input s_axis_fifo_22_tvalid,
    input [S_AXIS_FIFO_22_DMWIDTH/8-1:0] s_axis_fifo_22_tkeep,
    input [S_AXIS_FIFO_22_DMWIDTH/8-1:0] s_axis_fifo_22_tstrb,
    input [S_AXIS_FIFO_22_DMWIDTH-1:0] s_axis_fifo_22_tdata,
    output s_axis_fifo_22_tready,
    output ap_fifo_iarg_22_empty_n,
    output [S_AXIS_FIFO_22_WIDTH-1:0] ap_fifo_iarg_22_dout,
    input ap_fifo_iarg_22_read,
    //input AXI-Stream to FIFO interface 23
    input s_axis_fifo_23_aclk,
    input s_axis_fifo_23_aresetn,
    input s_axis_fifo_23_tlast,
    input s_axis_fifo_23_tvalid,
    input [S_AXIS_FIFO_23_DMWIDTH/8-1:0] s_axis_fifo_23_tkeep,
    input [S_AXIS_FIFO_23_DMWIDTH/8-1:0] s_axis_fifo_23_tstrb,
    input [S_AXIS_FIFO_23_DMWIDTH-1:0] s_axis_fifo_23_tdata,
    output s_axis_fifo_23_tready,
    output ap_fifo_iarg_23_empty_n,
    output [S_AXIS_FIFO_23_WIDTH-1:0] ap_fifo_iarg_23_dout,
    input ap_fifo_iarg_23_read,
    //input AXI-Stream to FIFO interface 24
    input s_axis_fifo_24_aclk,
    input s_axis_fifo_24_aresetn,
    input s_axis_fifo_24_tlast,
    input s_axis_fifo_24_tvalid,
    input [S_AXIS_FIFO_24_DMWIDTH/8-1:0] s_axis_fifo_24_tkeep,
    input [S_AXIS_FIFO_24_DMWIDTH/8-1:0] s_axis_fifo_24_tstrb,
    input [S_AXIS_FIFO_24_DMWIDTH-1:0] s_axis_fifo_24_tdata,
    output s_axis_fifo_24_tready,
    output ap_fifo_iarg_24_empty_n,
    output [S_AXIS_FIFO_24_WIDTH-1:0] ap_fifo_iarg_24_dout,
    input ap_fifo_iarg_24_read,
    //input AXI-Stream to FIFO interface 25
    input s_axis_fifo_25_aclk,
    input s_axis_fifo_25_aresetn,
    input s_axis_fifo_25_tlast,
    input s_axis_fifo_25_tvalid,
    input [S_AXIS_FIFO_25_DMWIDTH/8-1:0] s_axis_fifo_25_tkeep,
    input [S_AXIS_FIFO_25_DMWIDTH/8-1:0] s_axis_fifo_25_tstrb,
    input [S_AXIS_FIFO_25_DMWIDTH-1:0] s_axis_fifo_25_tdata,
    output s_axis_fifo_25_tready,
    output ap_fifo_iarg_25_empty_n,
    output [S_AXIS_FIFO_25_WIDTH-1:0] ap_fifo_iarg_25_dout,
    input ap_fifo_iarg_25_read,
    //input AXI-Stream to FIFO interface 26
    input s_axis_fifo_26_aclk,
    input s_axis_fifo_26_aresetn,
    input s_axis_fifo_26_tlast,
    input s_axis_fifo_26_tvalid,
    input [S_AXIS_FIFO_26_DMWIDTH/8-1:0] s_axis_fifo_26_tkeep,
    input [S_AXIS_FIFO_26_DMWIDTH/8-1:0] s_axis_fifo_26_tstrb,
    input [S_AXIS_FIFO_26_DMWIDTH-1:0] s_axis_fifo_26_tdata,
    output s_axis_fifo_26_tready,
    output ap_fifo_iarg_26_empty_n,
    output [S_AXIS_FIFO_26_WIDTH-1:0] ap_fifo_iarg_26_dout,
    input ap_fifo_iarg_26_read,
    //input AXI-Stream to FIFO interface 27
    input s_axis_fifo_27_aclk,
    input s_axis_fifo_27_aresetn,
    input s_axis_fifo_27_tlast,
    input s_axis_fifo_27_tvalid,
    input [S_AXIS_FIFO_27_DMWIDTH/8-1:0] s_axis_fifo_27_tkeep,
    input [S_AXIS_FIFO_27_DMWIDTH/8-1:0] s_axis_fifo_27_tstrb,
    input [S_AXIS_FIFO_27_DMWIDTH-1:0] s_axis_fifo_27_tdata,
    output s_axis_fifo_27_tready,
    output ap_fifo_iarg_27_empty_n,
    output [S_AXIS_FIFO_27_WIDTH-1:0] ap_fifo_iarg_27_dout,
    input ap_fifo_iarg_27_read,
    //input AXI-Stream to FIFO interface 28
    input s_axis_fifo_28_aclk,
    input s_axis_fifo_28_aresetn,
    input s_axis_fifo_28_tlast,
    input s_axis_fifo_28_tvalid,
    input [S_AXIS_FIFO_28_DMWIDTH/8-1:0] s_axis_fifo_28_tkeep,
    input [S_AXIS_FIFO_28_DMWIDTH/8-1:0] s_axis_fifo_28_tstrb,
    input [S_AXIS_FIFO_28_DMWIDTH-1:0] s_axis_fifo_28_tdata,
    output s_axis_fifo_28_tready,
    output ap_fifo_iarg_28_empty_n,
    output [S_AXIS_FIFO_28_WIDTH-1:0] ap_fifo_iarg_28_dout,
    input ap_fifo_iarg_28_read,
    //input AXI-Stream to FIFO interface 29
    input s_axis_fifo_29_aclk,
    input s_axis_fifo_29_aresetn,
    input s_axis_fifo_29_tlast,
    input s_axis_fifo_29_tvalid,
    input [S_AXIS_FIFO_29_DMWIDTH/8-1:0] s_axis_fifo_29_tkeep,
    input [S_AXIS_FIFO_29_DMWIDTH/8-1:0] s_axis_fifo_29_tstrb,
    input [S_AXIS_FIFO_29_DMWIDTH-1:0] s_axis_fifo_29_tdata,
    output s_axis_fifo_29_tready,
    output ap_fifo_iarg_29_empty_n,
    output [S_AXIS_FIFO_29_WIDTH-1:0] ap_fifo_iarg_29_dout,
    input ap_fifo_iarg_29_read,
    //input AXI-Stream to FIFO interface 30
    input s_axis_fifo_30_aclk,
    input s_axis_fifo_30_aresetn,
    input s_axis_fifo_30_tlast,
    input s_axis_fifo_30_tvalid,
    input [S_AXIS_FIFO_30_DMWIDTH/8-1:0] s_axis_fifo_30_tkeep,
    input [S_AXIS_FIFO_30_DMWIDTH/8-1:0] s_axis_fifo_30_tstrb,
    input [S_AXIS_FIFO_30_DMWIDTH-1:0] s_axis_fifo_30_tdata,
    output s_axis_fifo_30_tready,
    output ap_fifo_iarg_30_empty_n,
    output [S_AXIS_FIFO_30_WIDTH-1:0] ap_fifo_iarg_30_dout,
    input ap_fifo_iarg_30_read,
    //input AXI-Stream to FIFO interface 31
    input s_axis_fifo_31_aclk,
    input s_axis_fifo_31_aresetn,
    input s_axis_fifo_31_tlast,
    input s_axis_fifo_31_tvalid,
    input [S_AXIS_FIFO_31_DMWIDTH/8-1:0] s_axis_fifo_31_tkeep,
    input [S_AXIS_FIFO_31_DMWIDTH/8-1:0] s_axis_fifo_31_tstrb,
    input [S_AXIS_FIFO_31_DMWIDTH-1:0] s_axis_fifo_31_tdata,
    output s_axis_fifo_31_tready,
    output ap_fifo_iarg_31_empty_n,
    output [S_AXIS_FIFO_31_WIDTH-1:0] ap_fifo_iarg_31_dout,
    input ap_fifo_iarg_31_read,
    //input AXI-Stream to FIFO interface 32
    input s_axis_fifo_32_aclk,
    input s_axis_fifo_32_aresetn,
    input s_axis_fifo_32_tlast,
    input s_axis_fifo_32_tvalid,
    input [S_AXIS_FIFO_32_DMWIDTH/8-1:0] s_axis_fifo_32_tkeep,
    input [S_AXIS_FIFO_32_DMWIDTH/8-1:0] s_axis_fifo_32_tstrb,
    input [S_AXIS_FIFO_32_DMWIDTH-1:0] s_axis_fifo_32_tdata,
    output s_axis_fifo_32_tready,
    output ap_fifo_iarg_32_empty_n,
    output [S_AXIS_FIFO_32_WIDTH-1:0] ap_fifo_iarg_32_dout,
    input ap_fifo_iarg_32_read,
    //input AXI-Stream to FIFO interface 33
    input s_axis_fifo_33_aclk,
    input s_axis_fifo_33_aresetn,
    input s_axis_fifo_33_tlast,
    input s_axis_fifo_33_tvalid,
    input [S_AXIS_FIFO_33_DMWIDTH/8-1:0] s_axis_fifo_33_tkeep,
    input [S_AXIS_FIFO_33_DMWIDTH/8-1:0] s_axis_fifo_33_tstrb,
    input [S_AXIS_FIFO_33_DMWIDTH-1:0] s_axis_fifo_33_tdata,
    output s_axis_fifo_33_tready,
    output ap_fifo_iarg_33_empty_n,
    output [S_AXIS_FIFO_33_WIDTH-1:0] ap_fifo_iarg_33_dout,
    input ap_fifo_iarg_33_read,
    //input AXI-Stream to FIFO interface 34
    input s_axis_fifo_34_aclk,
    input s_axis_fifo_34_aresetn,
    input s_axis_fifo_34_tlast,
    input s_axis_fifo_34_tvalid,
    input [S_AXIS_FIFO_34_DMWIDTH/8-1:0] s_axis_fifo_34_tkeep,
    input [S_AXIS_FIFO_34_DMWIDTH/8-1:0] s_axis_fifo_34_tstrb,
    input [S_AXIS_FIFO_34_DMWIDTH-1:0] s_axis_fifo_34_tdata,
    output s_axis_fifo_34_tready,
    output ap_fifo_iarg_34_empty_n,
    output [S_AXIS_FIFO_34_WIDTH-1:0] ap_fifo_iarg_34_dout,
    input ap_fifo_iarg_34_read,
    //input AXI-Stream to FIFO interface 35
    input s_axis_fifo_35_aclk,
    input s_axis_fifo_35_aresetn,
    input s_axis_fifo_35_tlast,
    input s_axis_fifo_35_tvalid,
    input [S_AXIS_FIFO_35_DMWIDTH/8-1:0] s_axis_fifo_35_tkeep,
    input [S_AXIS_FIFO_35_DMWIDTH/8-1:0] s_axis_fifo_35_tstrb,
    input [S_AXIS_FIFO_35_DMWIDTH-1:0] s_axis_fifo_35_tdata,
    output s_axis_fifo_35_tready,
    output ap_fifo_iarg_35_empty_n,
    output [S_AXIS_FIFO_35_WIDTH-1:0] ap_fifo_iarg_35_dout,
    input ap_fifo_iarg_35_read,
    //input AXI-Stream to FIFO interface 36
    input s_axis_fifo_36_aclk,
    input s_axis_fifo_36_aresetn,
    input s_axis_fifo_36_tlast,
    input s_axis_fifo_36_tvalid,
    input [S_AXIS_FIFO_36_DMWIDTH/8-1:0] s_axis_fifo_36_tkeep,
    input [S_AXIS_FIFO_36_DMWIDTH/8-1:0] s_axis_fifo_36_tstrb,
    input [S_AXIS_FIFO_36_DMWIDTH-1:0] s_axis_fifo_36_tdata,
    output s_axis_fifo_36_tready,
    output ap_fifo_iarg_36_empty_n,
    output [S_AXIS_FIFO_36_WIDTH-1:0] ap_fifo_iarg_36_dout,
    input ap_fifo_iarg_36_read,
    //input AXI-Stream to FIFO interface 37
    input s_axis_fifo_37_aclk,
    input s_axis_fifo_37_aresetn,
    input s_axis_fifo_37_tlast,
    input s_axis_fifo_37_tvalid,
    input [S_AXIS_FIFO_37_DMWIDTH/8-1:0] s_axis_fifo_37_tkeep,
    input [S_AXIS_FIFO_37_DMWIDTH/8-1:0] s_axis_fifo_37_tstrb,
    input [S_AXIS_FIFO_37_DMWIDTH-1:0] s_axis_fifo_37_tdata,
    output s_axis_fifo_37_tready,
    output ap_fifo_iarg_37_empty_n,
    output [S_AXIS_FIFO_37_WIDTH-1:0] ap_fifo_iarg_37_dout,
    input ap_fifo_iarg_37_read,
    //input AXI-Stream to FIFO interface 38
    input s_axis_fifo_38_aclk,
    input s_axis_fifo_38_aresetn,
    input s_axis_fifo_38_tlast,
    input s_axis_fifo_38_tvalid,
    input [S_AXIS_FIFO_38_DMWIDTH/8-1:0] s_axis_fifo_38_tkeep,
    input [S_AXIS_FIFO_38_DMWIDTH/8-1:0] s_axis_fifo_38_tstrb,
    input [S_AXIS_FIFO_38_DMWIDTH-1:0] s_axis_fifo_38_tdata,
    output s_axis_fifo_38_tready,
    output ap_fifo_iarg_38_empty_n,
    output [S_AXIS_FIFO_38_WIDTH-1:0] ap_fifo_iarg_38_dout,
    input ap_fifo_iarg_38_read,
    //input AXI-Stream to FIFO interface 39
    input s_axis_fifo_39_aclk,
    input s_axis_fifo_39_aresetn,
    input s_axis_fifo_39_tlast,
    input s_axis_fifo_39_tvalid,
    input [S_AXIS_FIFO_39_DMWIDTH/8-1:0] s_axis_fifo_39_tkeep,
    input [S_AXIS_FIFO_39_DMWIDTH/8-1:0] s_axis_fifo_39_tstrb,
    input [S_AXIS_FIFO_39_DMWIDTH-1:0] s_axis_fifo_39_tdata,
    output s_axis_fifo_39_tready,
    output ap_fifo_iarg_39_empty_n,
    output [S_AXIS_FIFO_39_WIDTH-1:0] ap_fifo_iarg_39_dout,
    input ap_fifo_iarg_39_read,
    //input AXI-Stream to FIFO interface 40
    input s_axis_fifo_40_aclk,
    input s_axis_fifo_40_aresetn,
    input s_axis_fifo_40_tlast,
    input s_axis_fifo_40_tvalid,
    input [S_AXIS_FIFO_40_DMWIDTH/8-1:0] s_axis_fifo_40_tkeep,
    input [S_AXIS_FIFO_40_DMWIDTH/8-1:0] s_axis_fifo_40_tstrb,
    input [S_AXIS_FIFO_40_DMWIDTH-1:0] s_axis_fifo_40_tdata,
    output s_axis_fifo_40_tready,
    output ap_fifo_iarg_40_empty_n,
    output [S_AXIS_FIFO_40_WIDTH-1:0] ap_fifo_iarg_40_dout,
    input ap_fifo_iarg_40_read,
    //input AXI-Stream to FIFO interface 41
    input s_axis_fifo_41_aclk,
    input s_axis_fifo_41_aresetn,
    input s_axis_fifo_41_tlast,
    input s_axis_fifo_41_tvalid,
    input [S_AXIS_FIFO_41_DMWIDTH/8-1:0] s_axis_fifo_41_tkeep,
    input [S_AXIS_FIFO_41_DMWIDTH/8-1:0] s_axis_fifo_41_tstrb,
    input [S_AXIS_FIFO_41_DMWIDTH-1:0] s_axis_fifo_41_tdata,
    output s_axis_fifo_41_tready,
    output ap_fifo_iarg_41_empty_n,
    output [S_AXIS_FIFO_41_WIDTH-1:0] ap_fifo_iarg_41_dout,
    input ap_fifo_iarg_41_read,
    //input AXI-Stream to FIFO interface 42
    input s_axis_fifo_42_aclk,
    input s_axis_fifo_42_aresetn,
    input s_axis_fifo_42_tlast,
    input s_axis_fifo_42_tvalid,
    input [S_AXIS_FIFO_42_DMWIDTH/8-1:0] s_axis_fifo_42_tkeep,
    input [S_AXIS_FIFO_42_DMWIDTH/8-1:0] s_axis_fifo_42_tstrb,
    input [S_AXIS_FIFO_42_DMWIDTH-1:0] s_axis_fifo_42_tdata,
    output s_axis_fifo_42_tready,
    output ap_fifo_iarg_42_empty_n,
    output [S_AXIS_FIFO_42_WIDTH-1:0] ap_fifo_iarg_42_dout,
    input ap_fifo_iarg_42_read,
    //input AXI-Stream to FIFO interface 43
    input s_axis_fifo_43_aclk,
    input s_axis_fifo_43_aresetn,
    input s_axis_fifo_43_tlast,
    input s_axis_fifo_43_tvalid,
    input [S_AXIS_FIFO_43_DMWIDTH/8-1:0] s_axis_fifo_43_tkeep,
    input [S_AXIS_FIFO_43_DMWIDTH/8-1:0] s_axis_fifo_43_tstrb,
    input [S_AXIS_FIFO_43_DMWIDTH-1:0] s_axis_fifo_43_tdata,
    output s_axis_fifo_43_tready,
    output ap_fifo_iarg_43_empty_n,
    output [S_AXIS_FIFO_43_WIDTH-1:0] ap_fifo_iarg_43_dout,
    input ap_fifo_iarg_43_read,
    //input AXI-Stream to FIFO interface 44
    input s_axis_fifo_44_aclk,
    input s_axis_fifo_44_aresetn,
    input s_axis_fifo_44_tlast,
    input s_axis_fifo_44_tvalid,
    input [S_AXIS_FIFO_44_DMWIDTH/8-1:0] s_axis_fifo_44_tkeep,
    input [S_AXIS_FIFO_44_DMWIDTH/8-1:0] s_axis_fifo_44_tstrb,
    input [S_AXIS_FIFO_44_DMWIDTH-1:0] s_axis_fifo_44_tdata,
    output s_axis_fifo_44_tready,
    output ap_fifo_iarg_44_empty_n,
    output [S_AXIS_FIFO_44_WIDTH-1:0] ap_fifo_iarg_44_dout,
    input ap_fifo_iarg_44_read,
    //input AXI-Stream to FIFO interface 45
    input s_axis_fifo_45_aclk,
    input s_axis_fifo_45_aresetn,
    input s_axis_fifo_45_tlast,
    input s_axis_fifo_45_tvalid,
    input [S_AXIS_FIFO_45_DMWIDTH/8-1:0] s_axis_fifo_45_tkeep,
    input [S_AXIS_FIFO_45_DMWIDTH/8-1:0] s_axis_fifo_45_tstrb,
    input [S_AXIS_FIFO_45_DMWIDTH-1:0] s_axis_fifo_45_tdata,
    output s_axis_fifo_45_tready,
    output ap_fifo_iarg_45_empty_n,
    output [S_AXIS_FIFO_45_WIDTH-1:0] ap_fifo_iarg_45_dout,
    input ap_fifo_iarg_45_read,
    //input AXI-Stream to FIFO interface 46
    input s_axis_fifo_46_aclk,
    input s_axis_fifo_46_aresetn,
    input s_axis_fifo_46_tlast,
    input s_axis_fifo_46_tvalid,
    input [S_AXIS_FIFO_46_DMWIDTH/8-1:0] s_axis_fifo_46_tkeep,
    input [S_AXIS_FIFO_46_DMWIDTH/8-1:0] s_axis_fifo_46_tstrb,
    input [S_AXIS_FIFO_46_DMWIDTH-1:0] s_axis_fifo_46_tdata,
    output s_axis_fifo_46_tready,
    output ap_fifo_iarg_46_empty_n,
    output [S_AXIS_FIFO_46_WIDTH-1:0] ap_fifo_iarg_46_dout,
    input ap_fifo_iarg_46_read,
    //input AXI-Stream to FIFO interface 47
    input s_axis_fifo_47_aclk,
    input s_axis_fifo_47_aresetn,
    input s_axis_fifo_47_tlast,
    input s_axis_fifo_47_tvalid,
    input [S_AXIS_FIFO_47_DMWIDTH/8-1:0] s_axis_fifo_47_tkeep,
    input [S_AXIS_FIFO_47_DMWIDTH/8-1:0] s_axis_fifo_47_tstrb,
    input [S_AXIS_FIFO_47_DMWIDTH-1:0] s_axis_fifo_47_tdata,
    output s_axis_fifo_47_tready,
    output ap_fifo_iarg_47_empty_n,
    output [S_AXIS_FIFO_47_WIDTH-1:0] ap_fifo_iarg_47_dout,
    input ap_fifo_iarg_47_read,
    //input AXI-Stream to FIFO interface 48
    input s_axis_fifo_48_aclk,
    input s_axis_fifo_48_aresetn,
    input s_axis_fifo_48_tlast,
    input s_axis_fifo_48_tvalid,
    input [S_AXIS_FIFO_48_DMWIDTH/8-1:0] s_axis_fifo_48_tkeep,
    input [S_AXIS_FIFO_48_DMWIDTH/8-1:0] s_axis_fifo_48_tstrb,
    input [S_AXIS_FIFO_48_DMWIDTH-1:0] s_axis_fifo_48_tdata,
    output s_axis_fifo_48_tready,
    output ap_fifo_iarg_48_empty_n,
    output [S_AXIS_FIFO_48_WIDTH-1:0] ap_fifo_iarg_48_dout,
    input ap_fifo_iarg_48_read,
    //input AXI-Stream to FIFO interface 49
    input s_axis_fifo_49_aclk,
    input s_axis_fifo_49_aresetn,
    input s_axis_fifo_49_tlast,
    input s_axis_fifo_49_tvalid,
    input [S_AXIS_FIFO_49_DMWIDTH/8-1:0] s_axis_fifo_49_tkeep,
    input [S_AXIS_FIFO_49_DMWIDTH/8-1:0] s_axis_fifo_49_tstrb,
    input [S_AXIS_FIFO_49_DMWIDTH-1:0] s_axis_fifo_49_tdata,
    output s_axis_fifo_49_tready,
    output ap_fifo_iarg_49_empty_n,
    output [S_AXIS_FIFO_49_WIDTH-1:0] ap_fifo_iarg_49_dout,
    input ap_fifo_iarg_49_read,
    //input AXI-Stream to FIFO interface 50
    input s_axis_fifo_50_aclk,
    input s_axis_fifo_50_aresetn,
    input s_axis_fifo_50_tlast,
    input s_axis_fifo_50_tvalid,
    input [S_AXIS_FIFO_50_DMWIDTH/8-1:0] s_axis_fifo_50_tkeep,
    input [S_AXIS_FIFO_50_DMWIDTH/8-1:0] s_axis_fifo_50_tstrb,
    input [S_AXIS_FIFO_50_DMWIDTH-1:0] s_axis_fifo_50_tdata,
    output s_axis_fifo_50_tready,
    output ap_fifo_iarg_50_empty_n,
    output [S_AXIS_FIFO_50_WIDTH-1:0] ap_fifo_iarg_50_dout,
    input ap_fifo_iarg_50_read,
    //input AXI-Stream to FIFO interface 51
    input s_axis_fifo_51_aclk,
    input s_axis_fifo_51_aresetn,
    input s_axis_fifo_51_tlast,
    input s_axis_fifo_51_tvalid,
    input [S_AXIS_FIFO_51_DMWIDTH/8-1:0] s_axis_fifo_51_tkeep,
    input [S_AXIS_FIFO_51_DMWIDTH/8-1:0] s_axis_fifo_51_tstrb,
    input [S_AXIS_FIFO_51_DMWIDTH-1:0] s_axis_fifo_51_tdata,
    output s_axis_fifo_51_tready,
    output ap_fifo_iarg_51_empty_n,
    output [S_AXIS_FIFO_51_WIDTH-1:0] ap_fifo_iarg_51_dout,
    input ap_fifo_iarg_51_read,
    //input AXI-Stream to FIFO interface 52
    input s_axis_fifo_52_aclk,
    input s_axis_fifo_52_aresetn,
    input s_axis_fifo_52_tlast,
    input s_axis_fifo_52_tvalid,
    input [S_AXIS_FIFO_52_DMWIDTH/8-1:0] s_axis_fifo_52_tkeep,
    input [S_AXIS_FIFO_52_DMWIDTH/8-1:0] s_axis_fifo_52_tstrb,
    input [S_AXIS_FIFO_52_DMWIDTH-1:0] s_axis_fifo_52_tdata,
    output s_axis_fifo_52_tready,
    output ap_fifo_iarg_52_empty_n,
    output [S_AXIS_FIFO_52_WIDTH-1:0] ap_fifo_iarg_52_dout,
    input ap_fifo_iarg_52_read,
    //input AXI-Stream to FIFO interface 53
    input s_axis_fifo_53_aclk,
    input s_axis_fifo_53_aresetn,
    input s_axis_fifo_53_tlast,
    input s_axis_fifo_53_tvalid,
    input [S_AXIS_FIFO_53_DMWIDTH/8-1:0] s_axis_fifo_53_tkeep,
    input [S_AXIS_FIFO_53_DMWIDTH/8-1:0] s_axis_fifo_53_tstrb,
    input [S_AXIS_FIFO_53_DMWIDTH-1:0] s_axis_fifo_53_tdata,
    output s_axis_fifo_53_tready,
    output ap_fifo_iarg_53_empty_n,
    output [S_AXIS_FIFO_53_WIDTH-1:0] ap_fifo_iarg_53_dout,
    input ap_fifo_iarg_53_read,
    //input AXI-Stream to FIFO interface 54
    input s_axis_fifo_54_aclk,
    input s_axis_fifo_54_aresetn,
    input s_axis_fifo_54_tlast,
    input s_axis_fifo_54_tvalid,
    input [S_AXIS_FIFO_54_DMWIDTH/8-1:0] s_axis_fifo_54_tkeep,
    input [S_AXIS_FIFO_54_DMWIDTH/8-1:0] s_axis_fifo_54_tstrb,
    input [S_AXIS_FIFO_54_DMWIDTH-1:0] s_axis_fifo_54_tdata,
    output s_axis_fifo_54_tready,
    output ap_fifo_iarg_54_empty_n,
    output [S_AXIS_FIFO_54_WIDTH-1:0] ap_fifo_iarg_54_dout,
    input ap_fifo_iarg_54_read,
    //input AXI-Stream to FIFO interface 55
    input s_axis_fifo_55_aclk,
    input s_axis_fifo_55_aresetn,
    input s_axis_fifo_55_tlast,
    input s_axis_fifo_55_tvalid,
    input [S_AXIS_FIFO_55_DMWIDTH/8-1:0] s_axis_fifo_55_tkeep,
    input [S_AXIS_FIFO_55_DMWIDTH/8-1:0] s_axis_fifo_55_tstrb,
    input [S_AXIS_FIFO_55_DMWIDTH-1:0] s_axis_fifo_55_tdata,
    output s_axis_fifo_55_tready,
    output ap_fifo_iarg_55_empty_n,
    output [S_AXIS_FIFO_55_WIDTH-1:0] ap_fifo_iarg_55_dout,
    input ap_fifo_iarg_55_read,
    //input AXI-Stream to FIFO interface 56
    input s_axis_fifo_56_aclk,
    input s_axis_fifo_56_aresetn,
    input s_axis_fifo_56_tlast,
    input s_axis_fifo_56_tvalid,
    input [S_AXIS_FIFO_56_DMWIDTH/8-1:0] s_axis_fifo_56_tkeep,
    input [S_AXIS_FIFO_56_DMWIDTH/8-1:0] s_axis_fifo_56_tstrb,
    input [S_AXIS_FIFO_56_DMWIDTH-1:0] s_axis_fifo_56_tdata,
    output s_axis_fifo_56_tready,
    output ap_fifo_iarg_56_empty_n,
    output [S_AXIS_FIFO_56_WIDTH-1:0] ap_fifo_iarg_56_dout,
    input ap_fifo_iarg_56_read,
    //input AXI-Stream to FIFO interface 57
    input s_axis_fifo_57_aclk,
    input s_axis_fifo_57_aresetn,
    input s_axis_fifo_57_tlast,
    input s_axis_fifo_57_tvalid,
    input [S_AXIS_FIFO_57_DMWIDTH/8-1:0] s_axis_fifo_57_tkeep,
    input [S_AXIS_FIFO_57_DMWIDTH/8-1:0] s_axis_fifo_57_tstrb,
    input [S_AXIS_FIFO_57_DMWIDTH-1:0] s_axis_fifo_57_tdata,
    output s_axis_fifo_57_tready,
    output ap_fifo_iarg_57_empty_n,
    output [S_AXIS_FIFO_57_WIDTH-1:0] ap_fifo_iarg_57_dout,
    input ap_fifo_iarg_57_read,
    //input AXI-Stream to FIFO interface 58
    input s_axis_fifo_58_aclk,
    input s_axis_fifo_58_aresetn,
    input s_axis_fifo_58_tlast,
    input s_axis_fifo_58_tvalid,
    input [S_AXIS_FIFO_58_DMWIDTH/8-1:0] s_axis_fifo_58_tkeep,
    input [S_AXIS_FIFO_58_DMWIDTH/8-1:0] s_axis_fifo_58_tstrb,
    input [S_AXIS_FIFO_58_DMWIDTH-1:0] s_axis_fifo_58_tdata,
    output s_axis_fifo_58_tready,
    output ap_fifo_iarg_58_empty_n,
    output [S_AXIS_FIFO_58_WIDTH-1:0] ap_fifo_iarg_58_dout,
    input ap_fifo_iarg_58_read,
    //input AXI-Stream to FIFO interface 59
    input s_axis_fifo_59_aclk,
    input s_axis_fifo_59_aresetn,
    input s_axis_fifo_59_tlast,
    input s_axis_fifo_59_tvalid,
    input [S_AXIS_FIFO_59_DMWIDTH/8-1:0] s_axis_fifo_59_tkeep,
    input [S_AXIS_FIFO_59_DMWIDTH/8-1:0] s_axis_fifo_59_tstrb,
    input [S_AXIS_FIFO_59_DMWIDTH-1:0] s_axis_fifo_59_tdata,
    output s_axis_fifo_59_tready,
    output ap_fifo_iarg_59_empty_n,
    output [S_AXIS_FIFO_59_WIDTH-1:0] ap_fifo_iarg_59_dout,
    input ap_fifo_iarg_59_read,
    //input AXI-Stream to FIFO interface 60
    input s_axis_fifo_60_aclk,
    input s_axis_fifo_60_aresetn,
    input s_axis_fifo_60_tlast,
    input s_axis_fifo_60_tvalid,
    input [S_AXIS_FIFO_60_DMWIDTH/8-1:0] s_axis_fifo_60_tkeep,
    input [S_AXIS_FIFO_60_DMWIDTH/8-1:0] s_axis_fifo_60_tstrb,
    input [S_AXIS_FIFO_60_DMWIDTH-1:0] s_axis_fifo_60_tdata,
    output s_axis_fifo_60_tready,
    output ap_fifo_iarg_60_empty_n,
    output [S_AXIS_FIFO_60_WIDTH-1:0] ap_fifo_iarg_60_dout,
    input ap_fifo_iarg_60_read,
    //input AXI-Stream to FIFO interface 61
    input s_axis_fifo_61_aclk,
    input s_axis_fifo_61_aresetn,
    input s_axis_fifo_61_tlast,
    input s_axis_fifo_61_tvalid,
    input [S_AXIS_FIFO_61_DMWIDTH/8-1:0] s_axis_fifo_61_tkeep,
    input [S_AXIS_FIFO_61_DMWIDTH/8-1:0] s_axis_fifo_61_tstrb,
    input [S_AXIS_FIFO_61_DMWIDTH-1:0] s_axis_fifo_61_tdata,
    output s_axis_fifo_61_tready,
    output ap_fifo_iarg_61_empty_n,
    output [S_AXIS_FIFO_61_WIDTH-1:0] ap_fifo_iarg_61_dout,
    input ap_fifo_iarg_61_read,
    //input AXI-Stream to FIFO interface 62
    input s_axis_fifo_62_aclk,
    input s_axis_fifo_62_aresetn,
    input s_axis_fifo_62_tlast,
    input s_axis_fifo_62_tvalid,
    input [S_AXIS_FIFO_62_DMWIDTH/8-1:0] s_axis_fifo_62_tkeep,
    input [S_AXIS_FIFO_62_DMWIDTH/8-1:0] s_axis_fifo_62_tstrb,
    input [S_AXIS_FIFO_62_DMWIDTH-1:0] s_axis_fifo_62_tdata,
    output s_axis_fifo_62_tready,
    output ap_fifo_iarg_62_empty_n,
    output [S_AXIS_FIFO_62_WIDTH-1:0] ap_fifo_iarg_62_dout,
    input ap_fifo_iarg_62_read,
    //input AXI-Stream to FIFO interface 63
    input s_axis_fifo_63_aclk,
    input s_axis_fifo_63_aresetn,
    input s_axis_fifo_63_tlast,
    input s_axis_fifo_63_tvalid,
    input [S_AXIS_FIFO_63_DMWIDTH/8-1:0] s_axis_fifo_63_tkeep,
    input [S_AXIS_FIFO_63_DMWIDTH/8-1:0] s_axis_fifo_63_tstrb,
    input [S_AXIS_FIFO_63_DMWIDTH-1:0] s_axis_fifo_63_tdata,
    output s_axis_fifo_63_tready,
    output ap_fifo_iarg_63_empty_n,
    output [S_AXIS_FIFO_63_WIDTH-1:0] ap_fifo_iarg_63_dout,
    input ap_fifo_iarg_63_read,
    //input AXI-Stream to FIFO interface 64
    input s_axis_fifo_64_aclk,
    input s_axis_fifo_64_aresetn,
    input s_axis_fifo_64_tlast,
    input s_axis_fifo_64_tvalid,
    input [S_AXIS_FIFO_64_DMWIDTH/8-1:0] s_axis_fifo_64_tkeep,
    input [S_AXIS_FIFO_64_DMWIDTH/8-1:0] s_axis_fifo_64_tstrb,
    input [S_AXIS_FIFO_64_DMWIDTH-1:0] s_axis_fifo_64_tdata,
    output s_axis_fifo_64_tready,
    output ap_fifo_iarg_64_empty_n,
    output [S_AXIS_FIFO_64_WIDTH-1:0] ap_fifo_iarg_64_dout,
    input ap_fifo_iarg_64_read,
    //input AXI-Stream to FIFO interface 65
    input s_axis_fifo_65_aclk,
    input s_axis_fifo_65_aresetn,
    input s_axis_fifo_65_tlast,
    input s_axis_fifo_65_tvalid,
    input [S_AXIS_FIFO_65_DMWIDTH/8-1:0] s_axis_fifo_65_tkeep,
    input [S_AXIS_FIFO_65_DMWIDTH/8-1:0] s_axis_fifo_65_tstrb,
    input [S_AXIS_FIFO_65_DMWIDTH-1:0] s_axis_fifo_65_tdata,
    output s_axis_fifo_65_tready,
    output ap_fifo_iarg_65_empty_n,
    output [S_AXIS_FIFO_65_WIDTH-1:0] ap_fifo_iarg_65_dout,
    input ap_fifo_iarg_65_read,
    //input AXI-Stream to FIFO interface 66
    input s_axis_fifo_66_aclk,
    input s_axis_fifo_66_aresetn,
    input s_axis_fifo_66_tlast,
    input s_axis_fifo_66_tvalid,
    input [S_AXIS_FIFO_66_DMWIDTH/8-1:0] s_axis_fifo_66_tkeep,
    input [S_AXIS_FIFO_66_DMWIDTH/8-1:0] s_axis_fifo_66_tstrb,
    input [S_AXIS_FIFO_66_DMWIDTH-1:0] s_axis_fifo_66_tdata,
    output s_axis_fifo_66_tready,
    output ap_fifo_iarg_66_empty_n,
    output [S_AXIS_FIFO_66_WIDTH-1:0] ap_fifo_iarg_66_dout,
    input ap_fifo_iarg_66_read,
    //input AXI-Stream to FIFO interface 67
    input s_axis_fifo_67_aclk,
    input s_axis_fifo_67_aresetn,
    input s_axis_fifo_67_tlast,
    input s_axis_fifo_67_tvalid,
    input [S_AXIS_FIFO_67_DMWIDTH/8-1:0] s_axis_fifo_67_tkeep,
    input [S_AXIS_FIFO_67_DMWIDTH/8-1:0] s_axis_fifo_67_tstrb,
    input [S_AXIS_FIFO_67_DMWIDTH-1:0] s_axis_fifo_67_tdata,
    output s_axis_fifo_67_tready,
    output ap_fifo_iarg_67_empty_n,
    output [S_AXIS_FIFO_67_WIDTH-1:0] ap_fifo_iarg_67_dout,
    input ap_fifo_iarg_67_read,
    //input AXI-Stream to FIFO interface 68
    input s_axis_fifo_68_aclk,
    input s_axis_fifo_68_aresetn,
    input s_axis_fifo_68_tlast,
    input s_axis_fifo_68_tvalid,
    input [S_AXIS_FIFO_68_DMWIDTH/8-1:0] s_axis_fifo_68_tkeep,
    input [S_AXIS_FIFO_68_DMWIDTH/8-1:0] s_axis_fifo_68_tstrb,
    input [S_AXIS_FIFO_68_DMWIDTH-1:0] s_axis_fifo_68_tdata,
    output s_axis_fifo_68_tready,
    output ap_fifo_iarg_68_empty_n,
    output [S_AXIS_FIFO_68_WIDTH-1:0] ap_fifo_iarg_68_dout,
    input ap_fifo_iarg_68_read,
    //input AXI-Stream to FIFO interface 69
    input s_axis_fifo_69_aclk,
    input s_axis_fifo_69_aresetn,
    input s_axis_fifo_69_tlast,
    input s_axis_fifo_69_tvalid,
    input [S_AXIS_FIFO_69_DMWIDTH/8-1:0] s_axis_fifo_69_tkeep,
    input [S_AXIS_FIFO_69_DMWIDTH/8-1:0] s_axis_fifo_69_tstrb,
    input [S_AXIS_FIFO_69_DMWIDTH-1:0] s_axis_fifo_69_tdata,
    output s_axis_fifo_69_tready,
    output ap_fifo_iarg_69_empty_n,
    output [S_AXIS_FIFO_69_WIDTH-1:0] ap_fifo_iarg_69_dout,
    input ap_fifo_iarg_69_read,
    //input AXI-Stream to FIFO interface 70
    input s_axis_fifo_70_aclk,
    input s_axis_fifo_70_aresetn,
    input s_axis_fifo_70_tlast,
    input s_axis_fifo_70_tvalid,
    input [S_AXIS_FIFO_70_DMWIDTH/8-1:0] s_axis_fifo_70_tkeep,
    input [S_AXIS_FIFO_70_DMWIDTH/8-1:0] s_axis_fifo_70_tstrb,
    input [S_AXIS_FIFO_70_DMWIDTH-1:0] s_axis_fifo_70_tdata,
    output s_axis_fifo_70_tready,
    output ap_fifo_iarg_70_empty_n,
    output [S_AXIS_FIFO_70_WIDTH-1:0] ap_fifo_iarg_70_dout,
    input ap_fifo_iarg_70_read,
    //input AXI-Stream to FIFO interface 71
    input s_axis_fifo_71_aclk,
    input s_axis_fifo_71_aresetn,
    input s_axis_fifo_71_tlast,
    input s_axis_fifo_71_tvalid,
    input [S_AXIS_FIFO_71_DMWIDTH/8-1:0] s_axis_fifo_71_tkeep,
    input [S_AXIS_FIFO_71_DMWIDTH/8-1:0] s_axis_fifo_71_tstrb,
    input [S_AXIS_FIFO_71_DMWIDTH-1:0] s_axis_fifo_71_tdata,
    output s_axis_fifo_71_tready,
    output ap_fifo_iarg_71_empty_n,
    output [S_AXIS_FIFO_71_WIDTH-1:0] ap_fifo_iarg_71_dout,
    input ap_fifo_iarg_71_read,
    //input AXI-Stream to FIFO interface 72
    input s_axis_fifo_72_aclk,
    input s_axis_fifo_72_aresetn,
    input s_axis_fifo_72_tlast,
    input s_axis_fifo_72_tvalid,
    input [S_AXIS_FIFO_72_DMWIDTH/8-1:0] s_axis_fifo_72_tkeep,
    input [S_AXIS_FIFO_72_DMWIDTH/8-1:0] s_axis_fifo_72_tstrb,
    input [S_AXIS_FIFO_72_DMWIDTH-1:0] s_axis_fifo_72_tdata,
    output s_axis_fifo_72_tready,
    output ap_fifo_iarg_72_empty_n,
    output [S_AXIS_FIFO_72_WIDTH-1:0] ap_fifo_iarg_72_dout,
    input ap_fifo_iarg_72_read,
    //input AXI-Stream to FIFO interface 73
    input s_axis_fifo_73_aclk,
    input s_axis_fifo_73_aresetn,
    input s_axis_fifo_73_tlast,
    input s_axis_fifo_73_tvalid,
    input [S_AXIS_FIFO_73_DMWIDTH/8-1:0] s_axis_fifo_73_tkeep,
    input [S_AXIS_FIFO_73_DMWIDTH/8-1:0] s_axis_fifo_73_tstrb,
    input [S_AXIS_FIFO_73_DMWIDTH-1:0] s_axis_fifo_73_tdata,
    output s_axis_fifo_73_tready,
    output ap_fifo_iarg_73_empty_n,
    output [S_AXIS_FIFO_73_WIDTH-1:0] ap_fifo_iarg_73_dout,
    input ap_fifo_iarg_73_read,
    //input AXI-Stream to FIFO interface 74
    input s_axis_fifo_74_aclk,
    input s_axis_fifo_74_aresetn,
    input s_axis_fifo_74_tlast,
    input s_axis_fifo_74_tvalid,
    input [S_AXIS_FIFO_74_DMWIDTH/8-1:0] s_axis_fifo_74_tkeep,
    input [S_AXIS_FIFO_74_DMWIDTH/8-1:0] s_axis_fifo_74_tstrb,
    input [S_AXIS_FIFO_74_DMWIDTH-1:0] s_axis_fifo_74_tdata,
    output s_axis_fifo_74_tready,
    output ap_fifo_iarg_74_empty_n,
    output [S_AXIS_FIFO_74_WIDTH-1:0] ap_fifo_iarg_74_dout,
    input ap_fifo_iarg_74_read,
    //input AXI-Stream to FIFO interface 75
    input s_axis_fifo_75_aclk,
    input s_axis_fifo_75_aresetn,
    input s_axis_fifo_75_tlast,
    input s_axis_fifo_75_tvalid,
    input [S_AXIS_FIFO_75_DMWIDTH/8-1:0] s_axis_fifo_75_tkeep,
    input [S_AXIS_FIFO_75_DMWIDTH/8-1:0] s_axis_fifo_75_tstrb,
    input [S_AXIS_FIFO_75_DMWIDTH-1:0] s_axis_fifo_75_tdata,
    output s_axis_fifo_75_tready,
    output ap_fifo_iarg_75_empty_n,
    output [S_AXIS_FIFO_75_WIDTH-1:0] ap_fifo_iarg_75_dout,
    input ap_fifo_iarg_75_read,
    //input AXI-Stream to FIFO interface 76
    input s_axis_fifo_76_aclk,
    input s_axis_fifo_76_aresetn,
    input s_axis_fifo_76_tlast,
    input s_axis_fifo_76_tvalid,
    input [S_AXIS_FIFO_76_DMWIDTH/8-1:0] s_axis_fifo_76_tkeep,
    input [S_AXIS_FIFO_76_DMWIDTH/8-1:0] s_axis_fifo_76_tstrb,
    input [S_AXIS_FIFO_76_DMWIDTH-1:0] s_axis_fifo_76_tdata,
    output s_axis_fifo_76_tready,
    output ap_fifo_iarg_76_empty_n,
    output [S_AXIS_FIFO_76_WIDTH-1:0] ap_fifo_iarg_76_dout,
    input ap_fifo_iarg_76_read,
    //input AXI-Stream to FIFO interface 77
    input s_axis_fifo_77_aclk,
    input s_axis_fifo_77_aresetn,
    input s_axis_fifo_77_tlast,
    input s_axis_fifo_77_tvalid,
    input [S_AXIS_FIFO_77_DMWIDTH/8-1:0] s_axis_fifo_77_tkeep,
    input [S_AXIS_FIFO_77_DMWIDTH/8-1:0] s_axis_fifo_77_tstrb,
    input [S_AXIS_FIFO_77_DMWIDTH-1:0] s_axis_fifo_77_tdata,
    output s_axis_fifo_77_tready,
    output ap_fifo_iarg_77_empty_n,
    output [S_AXIS_FIFO_77_WIDTH-1:0] ap_fifo_iarg_77_dout,
    input ap_fifo_iarg_77_read,
    //input AXI-Stream to FIFO interface 78
    input s_axis_fifo_78_aclk,
    input s_axis_fifo_78_aresetn,
    input s_axis_fifo_78_tlast,
    input s_axis_fifo_78_tvalid,
    input [S_AXIS_FIFO_78_DMWIDTH/8-1:0] s_axis_fifo_78_tkeep,
    input [S_AXIS_FIFO_78_DMWIDTH/8-1:0] s_axis_fifo_78_tstrb,
    input [S_AXIS_FIFO_78_DMWIDTH-1:0] s_axis_fifo_78_tdata,
    output s_axis_fifo_78_tready,
    output ap_fifo_iarg_78_empty_n,
    output [S_AXIS_FIFO_78_WIDTH-1:0] ap_fifo_iarg_78_dout,
    input ap_fifo_iarg_78_read,
    //input AXI-Stream to FIFO interface 79
    input s_axis_fifo_79_aclk,
    input s_axis_fifo_79_aresetn,
    input s_axis_fifo_79_tlast,
    input s_axis_fifo_79_tvalid,
    input [S_AXIS_FIFO_79_DMWIDTH/8-1:0] s_axis_fifo_79_tkeep,
    input [S_AXIS_FIFO_79_DMWIDTH/8-1:0] s_axis_fifo_79_tstrb,
    input [S_AXIS_FIFO_79_DMWIDTH-1:0] s_axis_fifo_79_tdata,
    output s_axis_fifo_79_tready,
    output ap_fifo_iarg_79_empty_n,
    output [S_AXIS_FIFO_79_WIDTH-1:0] ap_fifo_iarg_79_dout,
    input ap_fifo_iarg_79_read,
    //input AXI-Stream to FIFO interface 80
    input s_axis_fifo_80_aclk,
    input s_axis_fifo_80_aresetn,
    input s_axis_fifo_80_tlast,
    input s_axis_fifo_80_tvalid,
    input [S_AXIS_FIFO_80_DMWIDTH/8-1:0] s_axis_fifo_80_tkeep,
    input [S_AXIS_FIFO_80_DMWIDTH/8-1:0] s_axis_fifo_80_tstrb,
    input [S_AXIS_FIFO_80_DMWIDTH-1:0] s_axis_fifo_80_tdata,
    output s_axis_fifo_80_tready,
    output ap_fifo_iarg_80_empty_n,
    output [S_AXIS_FIFO_80_WIDTH-1:0] ap_fifo_iarg_80_dout,
    input ap_fifo_iarg_80_read,
    //input AXI-Stream to FIFO interface 81
    input s_axis_fifo_81_aclk,
    input s_axis_fifo_81_aresetn,
    input s_axis_fifo_81_tlast,
    input s_axis_fifo_81_tvalid,
    input [S_AXIS_FIFO_81_DMWIDTH/8-1:0] s_axis_fifo_81_tkeep,
    input [S_AXIS_FIFO_81_DMWIDTH/8-1:0] s_axis_fifo_81_tstrb,
    input [S_AXIS_FIFO_81_DMWIDTH-1:0] s_axis_fifo_81_tdata,
    output s_axis_fifo_81_tready,
    output ap_fifo_iarg_81_empty_n,
    output [S_AXIS_FIFO_81_WIDTH-1:0] ap_fifo_iarg_81_dout,
    input ap_fifo_iarg_81_read,
    //input AXI-Stream to FIFO interface 82
    input s_axis_fifo_82_aclk,
    input s_axis_fifo_82_aresetn,
    input s_axis_fifo_82_tlast,
    input s_axis_fifo_82_tvalid,
    input [S_AXIS_FIFO_82_DMWIDTH/8-1:0] s_axis_fifo_82_tkeep,
    input [S_AXIS_FIFO_82_DMWIDTH/8-1:0] s_axis_fifo_82_tstrb,
    input [S_AXIS_FIFO_82_DMWIDTH-1:0] s_axis_fifo_82_tdata,
    output s_axis_fifo_82_tready,
    output ap_fifo_iarg_82_empty_n,
    output [S_AXIS_FIFO_82_WIDTH-1:0] ap_fifo_iarg_82_dout,
    input ap_fifo_iarg_82_read,
    //input AXI-Stream to FIFO interface 83
    input s_axis_fifo_83_aclk,
    input s_axis_fifo_83_aresetn,
    input s_axis_fifo_83_tlast,
    input s_axis_fifo_83_tvalid,
    input [S_AXIS_FIFO_83_DMWIDTH/8-1:0] s_axis_fifo_83_tkeep,
    input [S_AXIS_FIFO_83_DMWIDTH/8-1:0] s_axis_fifo_83_tstrb,
    input [S_AXIS_FIFO_83_DMWIDTH-1:0] s_axis_fifo_83_tdata,
    output s_axis_fifo_83_tready,
    output ap_fifo_iarg_83_empty_n,
    output [S_AXIS_FIFO_83_WIDTH-1:0] ap_fifo_iarg_83_dout,
    input ap_fifo_iarg_83_read,
    //input AXI-Stream to FIFO interface 84
    input s_axis_fifo_84_aclk,
    input s_axis_fifo_84_aresetn,
    input s_axis_fifo_84_tlast,
    input s_axis_fifo_84_tvalid,
    input [S_AXIS_FIFO_84_DMWIDTH/8-1:0] s_axis_fifo_84_tkeep,
    input [S_AXIS_FIFO_84_DMWIDTH/8-1:0] s_axis_fifo_84_tstrb,
    input [S_AXIS_FIFO_84_DMWIDTH-1:0] s_axis_fifo_84_tdata,
    output s_axis_fifo_84_tready,
    output ap_fifo_iarg_84_empty_n,
    output [S_AXIS_FIFO_84_WIDTH-1:0] ap_fifo_iarg_84_dout,
    input ap_fifo_iarg_84_read,
    //input AXI-Stream to FIFO interface 85
    input s_axis_fifo_85_aclk,
    input s_axis_fifo_85_aresetn,
    input s_axis_fifo_85_tlast,
    input s_axis_fifo_85_tvalid,
    input [S_AXIS_FIFO_85_DMWIDTH/8-1:0] s_axis_fifo_85_tkeep,
    input [S_AXIS_FIFO_85_DMWIDTH/8-1:0] s_axis_fifo_85_tstrb,
    input [S_AXIS_FIFO_85_DMWIDTH-1:0] s_axis_fifo_85_tdata,
    output s_axis_fifo_85_tready,
    output ap_fifo_iarg_85_empty_n,
    output [S_AXIS_FIFO_85_WIDTH-1:0] ap_fifo_iarg_85_dout,
    input ap_fifo_iarg_85_read,
    //input AXI-Stream to FIFO interface 86
    input s_axis_fifo_86_aclk,
    input s_axis_fifo_86_aresetn,
    input s_axis_fifo_86_tlast,
    input s_axis_fifo_86_tvalid,
    input [S_AXIS_FIFO_86_DMWIDTH/8-1:0] s_axis_fifo_86_tkeep,
    input [S_AXIS_FIFO_86_DMWIDTH/8-1:0] s_axis_fifo_86_tstrb,
    input [S_AXIS_FIFO_86_DMWIDTH-1:0] s_axis_fifo_86_tdata,
    output s_axis_fifo_86_tready,
    output ap_fifo_iarg_86_empty_n,
    output [S_AXIS_FIFO_86_WIDTH-1:0] ap_fifo_iarg_86_dout,
    input ap_fifo_iarg_86_read,
    //input AXI-Stream to FIFO interface 87
    input s_axis_fifo_87_aclk,
    input s_axis_fifo_87_aresetn,
    input s_axis_fifo_87_tlast,
    input s_axis_fifo_87_tvalid,
    input [S_AXIS_FIFO_87_DMWIDTH/8-1:0] s_axis_fifo_87_tkeep,
    input [S_AXIS_FIFO_87_DMWIDTH/8-1:0] s_axis_fifo_87_tstrb,
    input [S_AXIS_FIFO_87_DMWIDTH-1:0] s_axis_fifo_87_tdata,
    output s_axis_fifo_87_tready,
    output ap_fifo_iarg_87_empty_n,
    output [S_AXIS_FIFO_87_WIDTH-1:0] ap_fifo_iarg_87_dout,
    input ap_fifo_iarg_87_read,
    //input AXI-Stream to FIFO interface 88
    input s_axis_fifo_88_aclk,
    input s_axis_fifo_88_aresetn,
    input s_axis_fifo_88_tlast,
    input s_axis_fifo_88_tvalid,
    input [S_AXIS_FIFO_88_DMWIDTH/8-1:0] s_axis_fifo_88_tkeep,
    input [S_AXIS_FIFO_88_DMWIDTH/8-1:0] s_axis_fifo_88_tstrb,
    input [S_AXIS_FIFO_88_DMWIDTH-1:0] s_axis_fifo_88_tdata,
    output s_axis_fifo_88_tready,
    output ap_fifo_iarg_88_empty_n,
    output [S_AXIS_FIFO_88_WIDTH-1:0] ap_fifo_iarg_88_dout,
    input ap_fifo_iarg_88_read,
    //input AXI-Stream to FIFO interface 89
    input s_axis_fifo_89_aclk,
    input s_axis_fifo_89_aresetn,
    input s_axis_fifo_89_tlast,
    input s_axis_fifo_89_tvalid,
    input [S_AXIS_FIFO_89_DMWIDTH/8-1:0] s_axis_fifo_89_tkeep,
    input [S_AXIS_FIFO_89_DMWIDTH/8-1:0] s_axis_fifo_89_tstrb,
    input [S_AXIS_FIFO_89_DMWIDTH-1:0] s_axis_fifo_89_tdata,
    output s_axis_fifo_89_tready,
    output ap_fifo_iarg_89_empty_n,
    output [S_AXIS_FIFO_89_WIDTH-1:0] ap_fifo_iarg_89_dout,
    input ap_fifo_iarg_89_read,
    //input AXI-Stream to FIFO interface 90
    input s_axis_fifo_90_aclk,
    input s_axis_fifo_90_aresetn,
    input s_axis_fifo_90_tlast,
    input s_axis_fifo_90_tvalid,
    input [S_AXIS_FIFO_90_DMWIDTH/8-1:0] s_axis_fifo_90_tkeep,
    input [S_AXIS_FIFO_90_DMWIDTH/8-1:0] s_axis_fifo_90_tstrb,
    input [S_AXIS_FIFO_90_DMWIDTH-1:0] s_axis_fifo_90_tdata,
    output s_axis_fifo_90_tready,
    output ap_fifo_iarg_90_empty_n,
    output [S_AXIS_FIFO_90_WIDTH-1:0] ap_fifo_iarg_90_dout,
    input ap_fifo_iarg_90_read,
    //input AXI-Stream to FIFO interface 91
    input s_axis_fifo_91_aclk,
    input s_axis_fifo_91_aresetn,
    input s_axis_fifo_91_tlast,
    input s_axis_fifo_91_tvalid,
    input [S_AXIS_FIFO_91_DMWIDTH/8-1:0] s_axis_fifo_91_tkeep,
    input [S_AXIS_FIFO_91_DMWIDTH/8-1:0] s_axis_fifo_91_tstrb,
    input [S_AXIS_FIFO_91_DMWIDTH-1:0] s_axis_fifo_91_tdata,
    output s_axis_fifo_91_tready,
    output ap_fifo_iarg_91_empty_n,
    output [S_AXIS_FIFO_91_WIDTH-1:0] ap_fifo_iarg_91_dout,
    input ap_fifo_iarg_91_read,
    //input AXI-Stream to FIFO interface 92
    input s_axis_fifo_92_aclk,
    input s_axis_fifo_92_aresetn,
    input s_axis_fifo_92_tlast,
    input s_axis_fifo_92_tvalid,
    input [S_AXIS_FIFO_92_DMWIDTH/8-1:0] s_axis_fifo_92_tkeep,
    input [S_AXIS_FIFO_92_DMWIDTH/8-1:0] s_axis_fifo_92_tstrb,
    input [S_AXIS_FIFO_92_DMWIDTH-1:0] s_axis_fifo_92_tdata,
    output s_axis_fifo_92_tready,
    output ap_fifo_iarg_92_empty_n,
    output [S_AXIS_FIFO_92_WIDTH-1:0] ap_fifo_iarg_92_dout,
    input ap_fifo_iarg_92_read,
    //input AXI-Stream to FIFO interface 93
    input s_axis_fifo_93_aclk,
    input s_axis_fifo_93_aresetn,
    input s_axis_fifo_93_tlast,
    input s_axis_fifo_93_tvalid,
    input [S_AXIS_FIFO_93_DMWIDTH/8-1:0] s_axis_fifo_93_tkeep,
    input [S_AXIS_FIFO_93_DMWIDTH/8-1:0] s_axis_fifo_93_tstrb,
    input [S_AXIS_FIFO_93_DMWIDTH-1:0] s_axis_fifo_93_tdata,
    output s_axis_fifo_93_tready,
    output ap_fifo_iarg_93_empty_n,
    output [S_AXIS_FIFO_93_WIDTH-1:0] ap_fifo_iarg_93_dout,
    input ap_fifo_iarg_93_read,
    //input AXI-Stream to FIFO interface 94
    input s_axis_fifo_94_aclk,
    input s_axis_fifo_94_aresetn,
    input s_axis_fifo_94_tlast,
    input s_axis_fifo_94_tvalid,
    input [S_AXIS_FIFO_94_DMWIDTH/8-1:0] s_axis_fifo_94_tkeep,
    input [S_AXIS_FIFO_94_DMWIDTH/8-1:0] s_axis_fifo_94_tstrb,
    input [S_AXIS_FIFO_94_DMWIDTH-1:0] s_axis_fifo_94_tdata,
    output s_axis_fifo_94_tready,
    output ap_fifo_iarg_94_empty_n,
    output [S_AXIS_FIFO_94_WIDTH-1:0] ap_fifo_iarg_94_dout,
    input ap_fifo_iarg_94_read,
    //input AXI-Stream to FIFO interface 95
    input s_axis_fifo_95_aclk,
    input s_axis_fifo_95_aresetn,
    input s_axis_fifo_95_tlast,
    input s_axis_fifo_95_tvalid,
    input [S_AXIS_FIFO_95_DMWIDTH/8-1:0] s_axis_fifo_95_tkeep,
    input [S_AXIS_FIFO_95_DMWIDTH/8-1:0] s_axis_fifo_95_tstrb,
    input [S_AXIS_FIFO_95_DMWIDTH-1:0] s_axis_fifo_95_tdata,
    output s_axis_fifo_95_tready,
    output ap_fifo_iarg_95_empty_n,
    output [S_AXIS_FIFO_95_WIDTH-1:0] ap_fifo_iarg_95_dout,
    input ap_fifo_iarg_95_read,
    //input AXI-Stream to FIFO interface 96
    input s_axis_fifo_96_aclk,
    input s_axis_fifo_96_aresetn,
    input s_axis_fifo_96_tlast,
    input s_axis_fifo_96_tvalid,
    input [S_AXIS_FIFO_96_DMWIDTH/8-1:0] s_axis_fifo_96_tkeep,
    input [S_AXIS_FIFO_96_DMWIDTH/8-1:0] s_axis_fifo_96_tstrb,
    input [S_AXIS_FIFO_96_DMWIDTH-1:0] s_axis_fifo_96_tdata,
    output s_axis_fifo_96_tready,
    output ap_fifo_iarg_96_empty_n,
    output [S_AXIS_FIFO_96_WIDTH-1:0] ap_fifo_iarg_96_dout,
    input ap_fifo_iarg_96_read,
    //input AXI-Stream to FIFO interface 97
    input s_axis_fifo_97_aclk,
    input s_axis_fifo_97_aresetn,
    input s_axis_fifo_97_tlast,
    input s_axis_fifo_97_tvalid,
    input [S_AXIS_FIFO_97_DMWIDTH/8-1:0] s_axis_fifo_97_tkeep,
    input [S_AXIS_FIFO_97_DMWIDTH/8-1:0] s_axis_fifo_97_tstrb,
    input [S_AXIS_FIFO_97_DMWIDTH-1:0] s_axis_fifo_97_tdata,
    output s_axis_fifo_97_tready,
    output ap_fifo_iarg_97_empty_n,
    output [S_AXIS_FIFO_97_WIDTH-1:0] ap_fifo_iarg_97_dout,
    input ap_fifo_iarg_97_read,
    //input AXI-Stream to FIFO interface 98
    input s_axis_fifo_98_aclk,
    input s_axis_fifo_98_aresetn,
    input s_axis_fifo_98_tlast,
    input s_axis_fifo_98_tvalid,
    input [S_AXIS_FIFO_98_DMWIDTH/8-1:0] s_axis_fifo_98_tkeep,
    input [S_AXIS_FIFO_98_DMWIDTH/8-1:0] s_axis_fifo_98_tstrb,
    input [S_AXIS_FIFO_98_DMWIDTH-1:0] s_axis_fifo_98_tdata,
    output s_axis_fifo_98_tready,
    output ap_fifo_iarg_98_empty_n,
    output [S_AXIS_FIFO_98_WIDTH-1:0] ap_fifo_iarg_98_dout,
    input ap_fifo_iarg_98_read,
    //input AXI-Stream to FIFO interface 99
    input s_axis_fifo_99_aclk,
    input s_axis_fifo_99_aresetn,
    input s_axis_fifo_99_tlast,
    input s_axis_fifo_99_tvalid,
    input [S_AXIS_FIFO_99_DMWIDTH/8-1:0] s_axis_fifo_99_tkeep,
    input [S_AXIS_FIFO_99_DMWIDTH/8-1:0] s_axis_fifo_99_tstrb,
    input [S_AXIS_FIFO_99_DMWIDTH-1:0] s_axis_fifo_99_tdata,
    output s_axis_fifo_99_tready,
    output ap_fifo_iarg_99_empty_n,
    output [S_AXIS_FIFO_99_WIDTH-1:0] ap_fifo_iarg_99_dout,
    input ap_fifo_iarg_99_read,
    //input AXI-Stream to FIFO interface 100
    input s_axis_fifo_100_aclk,
    input s_axis_fifo_100_aresetn,
    input s_axis_fifo_100_tlast,
    input s_axis_fifo_100_tvalid,
    input [S_AXIS_FIFO_100_DMWIDTH/8-1:0] s_axis_fifo_100_tkeep,
    input [S_AXIS_FIFO_100_DMWIDTH/8-1:0] s_axis_fifo_100_tstrb,
    input [S_AXIS_FIFO_100_DMWIDTH-1:0] s_axis_fifo_100_tdata,
    output s_axis_fifo_100_tready,
    output ap_fifo_iarg_100_empty_n,
    output [S_AXIS_FIFO_100_WIDTH-1:0] ap_fifo_iarg_100_dout,
    input ap_fifo_iarg_100_read,
    //input AXI-Stream to FIFO interface 101
    input s_axis_fifo_101_aclk,
    input s_axis_fifo_101_aresetn,
    input s_axis_fifo_101_tlast,
    input s_axis_fifo_101_tvalid,
    input [S_AXIS_FIFO_101_DMWIDTH/8-1:0] s_axis_fifo_101_tkeep,
    input [S_AXIS_FIFO_101_DMWIDTH/8-1:0] s_axis_fifo_101_tstrb,
    input [S_AXIS_FIFO_101_DMWIDTH-1:0] s_axis_fifo_101_tdata,
    output s_axis_fifo_101_tready,
    output ap_fifo_iarg_101_empty_n,
    output [S_AXIS_FIFO_101_WIDTH-1:0] ap_fifo_iarg_101_dout,
    input ap_fifo_iarg_101_read,
    //input AXI-Stream to FIFO interface 102
    input s_axis_fifo_102_aclk,
    input s_axis_fifo_102_aresetn,
    input s_axis_fifo_102_tlast,
    input s_axis_fifo_102_tvalid,
    input [S_AXIS_FIFO_102_DMWIDTH/8-1:0] s_axis_fifo_102_tkeep,
    input [S_AXIS_FIFO_102_DMWIDTH/8-1:0] s_axis_fifo_102_tstrb,
    input [S_AXIS_FIFO_102_DMWIDTH-1:0] s_axis_fifo_102_tdata,
    output s_axis_fifo_102_tready,
    output ap_fifo_iarg_102_empty_n,
    output [S_AXIS_FIFO_102_WIDTH-1:0] ap_fifo_iarg_102_dout,
    input ap_fifo_iarg_102_read,
    //input AXI-Stream to FIFO interface 103
    input s_axis_fifo_103_aclk,
    input s_axis_fifo_103_aresetn,
    input s_axis_fifo_103_tlast,
    input s_axis_fifo_103_tvalid,
    input [S_AXIS_FIFO_103_DMWIDTH/8-1:0] s_axis_fifo_103_tkeep,
    input [S_AXIS_FIFO_103_DMWIDTH/8-1:0] s_axis_fifo_103_tstrb,
    input [S_AXIS_FIFO_103_DMWIDTH-1:0] s_axis_fifo_103_tdata,
    output s_axis_fifo_103_tready,
    output ap_fifo_iarg_103_empty_n,
    output [S_AXIS_FIFO_103_WIDTH-1:0] ap_fifo_iarg_103_dout,
    input ap_fifo_iarg_103_read,
    //input AXI-Stream to FIFO interface 104
    input s_axis_fifo_104_aclk,
    input s_axis_fifo_104_aresetn,
    input s_axis_fifo_104_tlast,
    input s_axis_fifo_104_tvalid,
    input [S_AXIS_FIFO_104_DMWIDTH/8-1:0] s_axis_fifo_104_tkeep,
    input [S_AXIS_FIFO_104_DMWIDTH/8-1:0] s_axis_fifo_104_tstrb,
    input [S_AXIS_FIFO_104_DMWIDTH-1:0] s_axis_fifo_104_tdata,
    output s_axis_fifo_104_tready,
    output ap_fifo_iarg_104_empty_n,
    output [S_AXIS_FIFO_104_WIDTH-1:0] ap_fifo_iarg_104_dout,
    input ap_fifo_iarg_104_read,
    //input AXI-Stream to FIFO interface 105
    input s_axis_fifo_105_aclk,
    input s_axis_fifo_105_aresetn,
    input s_axis_fifo_105_tlast,
    input s_axis_fifo_105_tvalid,
    input [S_AXIS_FIFO_105_DMWIDTH/8-1:0] s_axis_fifo_105_tkeep,
    input [S_AXIS_FIFO_105_DMWIDTH/8-1:0] s_axis_fifo_105_tstrb,
    input [S_AXIS_FIFO_105_DMWIDTH-1:0] s_axis_fifo_105_tdata,
    output s_axis_fifo_105_tready,
    output ap_fifo_iarg_105_empty_n,
    output [S_AXIS_FIFO_105_WIDTH-1:0] ap_fifo_iarg_105_dout,
    input ap_fifo_iarg_105_read,
    //input AXI-Stream to FIFO interface 106
    input s_axis_fifo_106_aclk,
    input s_axis_fifo_106_aresetn,
    input s_axis_fifo_106_tlast,
    input s_axis_fifo_106_tvalid,
    input [S_AXIS_FIFO_106_DMWIDTH/8-1:0] s_axis_fifo_106_tkeep,
    input [S_AXIS_FIFO_106_DMWIDTH/8-1:0] s_axis_fifo_106_tstrb,
    input [S_AXIS_FIFO_106_DMWIDTH-1:0] s_axis_fifo_106_tdata,
    output s_axis_fifo_106_tready,
    output ap_fifo_iarg_106_empty_n,
    output [S_AXIS_FIFO_106_WIDTH-1:0] ap_fifo_iarg_106_dout,
    input ap_fifo_iarg_106_read,
    //input AXI-Stream to FIFO interface 107
    input s_axis_fifo_107_aclk,
    input s_axis_fifo_107_aresetn,
    input s_axis_fifo_107_tlast,
    input s_axis_fifo_107_tvalid,
    input [S_AXIS_FIFO_107_DMWIDTH/8-1:0] s_axis_fifo_107_tkeep,
    input [S_AXIS_FIFO_107_DMWIDTH/8-1:0] s_axis_fifo_107_tstrb,
    input [S_AXIS_FIFO_107_DMWIDTH-1:0] s_axis_fifo_107_tdata,
    output s_axis_fifo_107_tready,
    output ap_fifo_iarg_107_empty_n,
    output [S_AXIS_FIFO_107_WIDTH-1:0] ap_fifo_iarg_107_dout,
    input ap_fifo_iarg_107_read,
    //input AXI-Stream to FIFO interface 108
    input s_axis_fifo_108_aclk,
    input s_axis_fifo_108_aresetn,
    input s_axis_fifo_108_tlast,
    input s_axis_fifo_108_tvalid,
    input [S_AXIS_FIFO_108_DMWIDTH/8-1:0] s_axis_fifo_108_tkeep,
    input [S_AXIS_FIFO_108_DMWIDTH/8-1:0] s_axis_fifo_108_tstrb,
    input [S_AXIS_FIFO_108_DMWIDTH-1:0] s_axis_fifo_108_tdata,
    output s_axis_fifo_108_tready,
    output ap_fifo_iarg_108_empty_n,
    output [S_AXIS_FIFO_108_WIDTH-1:0] ap_fifo_iarg_108_dout,
    input ap_fifo_iarg_108_read,
    //input AXI-Stream to FIFO interface 109
    input s_axis_fifo_109_aclk,
    input s_axis_fifo_109_aresetn,
    input s_axis_fifo_109_tlast,
    input s_axis_fifo_109_tvalid,
    input [S_AXIS_FIFO_109_DMWIDTH/8-1:0] s_axis_fifo_109_tkeep,
    input [S_AXIS_FIFO_109_DMWIDTH/8-1:0] s_axis_fifo_109_tstrb,
    input [S_AXIS_FIFO_109_DMWIDTH-1:0] s_axis_fifo_109_tdata,
    output s_axis_fifo_109_tready,
    output ap_fifo_iarg_109_empty_n,
    output [S_AXIS_FIFO_109_WIDTH-1:0] ap_fifo_iarg_109_dout,
    input ap_fifo_iarg_109_read,
    //input AXI-Stream to FIFO interface 110
    input s_axis_fifo_110_aclk,
    input s_axis_fifo_110_aresetn,
    input s_axis_fifo_110_tlast,
    input s_axis_fifo_110_tvalid,
    input [S_AXIS_FIFO_110_DMWIDTH/8-1:0] s_axis_fifo_110_tkeep,
    input [S_AXIS_FIFO_110_DMWIDTH/8-1:0] s_axis_fifo_110_tstrb,
    input [S_AXIS_FIFO_110_DMWIDTH-1:0] s_axis_fifo_110_tdata,
    output s_axis_fifo_110_tready,
    output ap_fifo_iarg_110_empty_n,
    output [S_AXIS_FIFO_110_WIDTH-1:0] ap_fifo_iarg_110_dout,
    input ap_fifo_iarg_110_read,
    //input AXI-Stream to FIFO interface 111
    input s_axis_fifo_111_aclk,
    input s_axis_fifo_111_aresetn,
    input s_axis_fifo_111_tlast,
    input s_axis_fifo_111_tvalid,
    input [S_AXIS_FIFO_111_DMWIDTH/8-1:0] s_axis_fifo_111_tkeep,
    input [S_AXIS_FIFO_111_DMWIDTH/8-1:0] s_axis_fifo_111_tstrb,
    input [S_AXIS_FIFO_111_DMWIDTH-1:0] s_axis_fifo_111_tdata,
    output s_axis_fifo_111_tready,
    output ap_fifo_iarg_111_empty_n,
    output [S_AXIS_FIFO_111_WIDTH-1:0] ap_fifo_iarg_111_dout,
    input ap_fifo_iarg_111_read,
    //input AXI-Stream to FIFO interface 112
    input s_axis_fifo_112_aclk,
    input s_axis_fifo_112_aresetn,
    input s_axis_fifo_112_tlast,
    input s_axis_fifo_112_tvalid,
    input [S_AXIS_FIFO_112_DMWIDTH/8-1:0] s_axis_fifo_112_tkeep,
    input [S_AXIS_FIFO_112_DMWIDTH/8-1:0] s_axis_fifo_112_tstrb,
    input [S_AXIS_FIFO_112_DMWIDTH-1:0] s_axis_fifo_112_tdata,
    output s_axis_fifo_112_tready,
    output ap_fifo_iarg_112_empty_n,
    output [S_AXIS_FIFO_112_WIDTH-1:0] ap_fifo_iarg_112_dout,
    input ap_fifo_iarg_112_read,
    //input AXI-Stream to FIFO interface 113
    input s_axis_fifo_113_aclk,
    input s_axis_fifo_113_aresetn,
    input s_axis_fifo_113_tlast,
    input s_axis_fifo_113_tvalid,
    input [S_AXIS_FIFO_113_DMWIDTH/8-1:0] s_axis_fifo_113_tkeep,
    input [S_AXIS_FIFO_113_DMWIDTH/8-1:0] s_axis_fifo_113_tstrb,
    input [S_AXIS_FIFO_113_DMWIDTH-1:0] s_axis_fifo_113_tdata,
    output s_axis_fifo_113_tready,
    output ap_fifo_iarg_113_empty_n,
    output [S_AXIS_FIFO_113_WIDTH-1:0] ap_fifo_iarg_113_dout,
    input ap_fifo_iarg_113_read,
    //input AXI-Stream to FIFO interface 114
    input s_axis_fifo_114_aclk,
    input s_axis_fifo_114_aresetn,
    input s_axis_fifo_114_tlast,
    input s_axis_fifo_114_tvalid,
    input [S_AXIS_FIFO_114_DMWIDTH/8-1:0] s_axis_fifo_114_tkeep,
    input [S_AXIS_FIFO_114_DMWIDTH/8-1:0] s_axis_fifo_114_tstrb,
    input [S_AXIS_FIFO_114_DMWIDTH-1:0] s_axis_fifo_114_tdata,
    output s_axis_fifo_114_tready,
    output ap_fifo_iarg_114_empty_n,
    output [S_AXIS_FIFO_114_WIDTH-1:0] ap_fifo_iarg_114_dout,
    input ap_fifo_iarg_114_read,
    //input AXI-Stream to FIFO interface 115
    input s_axis_fifo_115_aclk,
    input s_axis_fifo_115_aresetn,
    input s_axis_fifo_115_tlast,
    input s_axis_fifo_115_tvalid,
    input [S_AXIS_FIFO_115_DMWIDTH/8-1:0] s_axis_fifo_115_tkeep,
    input [S_AXIS_FIFO_115_DMWIDTH/8-1:0] s_axis_fifo_115_tstrb,
    input [S_AXIS_FIFO_115_DMWIDTH-1:0] s_axis_fifo_115_tdata,
    output s_axis_fifo_115_tready,
    output ap_fifo_iarg_115_empty_n,
    output [S_AXIS_FIFO_115_WIDTH-1:0] ap_fifo_iarg_115_dout,
    input ap_fifo_iarg_115_read,
    //input AXI-Stream to FIFO interface 116
    input s_axis_fifo_116_aclk,
    input s_axis_fifo_116_aresetn,
    input s_axis_fifo_116_tlast,
    input s_axis_fifo_116_tvalid,
    input [S_AXIS_FIFO_116_DMWIDTH/8-1:0] s_axis_fifo_116_tkeep,
    input [S_AXIS_FIFO_116_DMWIDTH/8-1:0] s_axis_fifo_116_tstrb,
    input [S_AXIS_FIFO_116_DMWIDTH-1:0] s_axis_fifo_116_tdata,
    output s_axis_fifo_116_tready,
    output ap_fifo_iarg_116_empty_n,
    output [S_AXIS_FIFO_116_WIDTH-1:0] ap_fifo_iarg_116_dout,
    input ap_fifo_iarg_116_read,
    //input AXI-Stream to FIFO interface 117
    input s_axis_fifo_117_aclk,
    input s_axis_fifo_117_aresetn,
    input s_axis_fifo_117_tlast,
    input s_axis_fifo_117_tvalid,
    input [S_AXIS_FIFO_117_DMWIDTH/8-1:0] s_axis_fifo_117_tkeep,
    input [S_AXIS_FIFO_117_DMWIDTH/8-1:0] s_axis_fifo_117_tstrb,
    input [S_AXIS_FIFO_117_DMWIDTH-1:0] s_axis_fifo_117_tdata,
    output s_axis_fifo_117_tready,
    output ap_fifo_iarg_117_empty_n,
    output [S_AXIS_FIFO_117_WIDTH-1:0] ap_fifo_iarg_117_dout,
    input ap_fifo_iarg_117_read,
    //input AXI-Stream to FIFO interface 118
    input s_axis_fifo_118_aclk,
    input s_axis_fifo_118_aresetn,
    input s_axis_fifo_118_tlast,
    input s_axis_fifo_118_tvalid,
    input [S_AXIS_FIFO_118_DMWIDTH/8-1:0] s_axis_fifo_118_tkeep,
    input [S_AXIS_FIFO_118_DMWIDTH/8-1:0] s_axis_fifo_118_tstrb,
    input [S_AXIS_FIFO_118_DMWIDTH-1:0] s_axis_fifo_118_tdata,
    output s_axis_fifo_118_tready,
    output ap_fifo_iarg_118_empty_n,
    output [S_AXIS_FIFO_118_WIDTH-1:0] ap_fifo_iarg_118_dout,
    input ap_fifo_iarg_118_read,
    //input AXI-Stream to FIFO interface 119
    input s_axis_fifo_119_aclk,
    input s_axis_fifo_119_aresetn,
    input s_axis_fifo_119_tlast,
    input s_axis_fifo_119_tvalid,
    input [S_AXIS_FIFO_119_DMWIDTH/8-1:0] s_axis_fifo_119_tkeep,
    input [S_AXIS_FIFO_119_DMWIDTH/8-1:0] s_axis_fifo_119_tstrb,
    input [S_AXIS_FIFO_119_DMWIDTH-1:0] s_axis_fifo_119_tdata,
    output s_axis_fifo_119_tready,
    output ap_fifo_iarg_119_empty_n,
    output [S_AXIS_FIFO_119_WIDTH-1:0] ap_fifo_iarg_119_dout,
    input ap_fifo_iarg_119_read,
    //input AXI-Stream to FIFO interface 120
    input s_axis_fifo_120_aclk,
    input s_axis_fifo_120_aresetn,
    input s_axis_fifo_120_tlast,
    input s_axis_fifo_120_tvalid,
    input [S_AXIS_FIFO_120_DMWIDTH/8-1:0] s_axis_fifo_120_tkeep,
    input [S_AXIS_FIFO_120_DMWIDTH/8-1:0] s_axis_fifo_120_tstrb,
    input [S_AXIS_FIFO_120_DMWIDTH-1:0] s_axis_fifo_120_tdata,
    output s_axis_fifo_120_tready,
    output ap_fifo_iarg_120_empty_n,
    output [S_AXIS_FIFO_120_WIDTH-1:0] ap_fifo_iarg_120_dout,
    input ap_fifo_iarg_120_read,
    //input AXI-Stream to FIFO interface 121
    input s_axis_fifo_121_aclk,
    input s_axis_fifo_121_aresetn,
    input s_axis_fifo_121_tlast,
    input s_axis_fifo_121_tvalid,
    input [S_AXIS_FIFO_121_DMWIDTH/8-1:0] s_axis_fifo_121_tkeep,
    input [S_AXIS_FIFO_121_DMWIDTH/8-1:0] s_axis_fifo_121_tstrb,
    input [S_AXIS_FIFO_121_DMWIDTH-1:0] s_axis_fifo_121_tdata,
    output s_axis_fifo_121_tready,
    output ap_fifo_iarg_121_empty_n,
    output [S_AXIS_FIFO_121_WIDTH-1:0] ap_fifo_iarg_121_dout,
    input ap_fifo_iarg_121_read,
    //input AXI-Stream to FIFO interface 122
    input s_axis_fifo_122_aclk,
    input s_axis_fifo_122_aresetn,
    input s_axis_fifo_122_tlast,
    input s_axis_fifo_122_tvalid,
    input [S_AXIS_FIFO_122_DMWIDTH/8-1:0] s_axis_fifo_122_tkeep,
    input [S_AXIS_FIFO_122_DMWIDTH/8-1:0] s_axis_fifo_122_tstrb,
    input [S_AXIS_FIFO_122_DMWIDTH-1:0] s_axis_fifo_122_tdata,
    output s_axis_fifo_122_tready,
    output ap_fifo_iarg_122_empty_n,
    output [S_AXIS_FIFO_122_WIDTH-1:0] ap_fifo_iarg_122_dout,
    input ap_fifo_iarg_122_read,
    //input AXI-Stream to FIFO interface 123
    input s_axis_fifo_123_aclk,
    input s_axis_fifo_123_aresetn,
    input s_axis_fifo_123_tlast,
    input s_axis_fifo_123_tvalid,
    input [S_AXIS_FIFO_123_DMWIDTH/8-1:0] s_axis_fifo_123_tkeep,
    input [S_AXIS_FIFO_123_DMWIDTH/8-1:0] s_axis_fifo_123_tstrb,
    input [S_AXIS_FIFO_123_DMWIDTH-1:0] s_axis_fifo_123_tdata,
    output s_axis_fifo_123_tready,
    output ap_fifo_iarg_123_empty_n,
    output [S_AXIS_FIFO_123_WIDTH-1:0] ap_fifo_iarg_123_dout,
    input ap_fifo_iarg_123_read,
    //input AXI-Stream to FIFO interface 124
    input s_axis_fifo_124_aclk,
    input s_axis_fifo_124_aresetn,
    input s_axis_fifo_124_tlast,
    input s_axis_fifo_124_tvalid,
    input [S_AXIS_FIFO_124_DMWIDTH/8-1:0] s_axis_fifo_124_tkeep,
    input [S_AXIS_FIFO_124_DMWIDTH/8-1:0] s_axis_fifo_124_tstrb,
    input [S_AXIS_FIFO_124_DMWIDTH-1:0] s_axis_fifo_124_tdata,
    output s_axis_fifo_124_tready,
    output ap_fifo_iarg_124_empty_n,
    output [S_AXIS_FIFO_124_WIDTH-1:0] ap_fifo_iarg_124_dout,
    input ap_fifo_iarg_124_read,
    //input AXI-Stream to FIFO interface 125
    input s_axis_fifo_125_aclk,
    input s_axis_fifo_125_aresetn,
    input s_axis_fifo_125_tlast,
    input s_axis_fifo_125_tvalid,
    input [S_AXIS_FIFO_125_DMWIDTH/8-1:0] s_axis_fifo_125_tkeep,
    input [S_AXIS_FIFO_125_DMWIDTH/8-1:0] s_axis_fifo_125_tstrb,
    input [S_AXIS_FIFO_125_DMWIDTH-1:0] s_axis_fifo_125_tdata,
    output s_axis_fifo_125_tready,
    output ap_fifo_iarg_125_empty_n,
    output [S_AXIS_FIFO_125_WIDTH-1:0] ap_fifo_iarg_125_dout,
    input ap_fifo_iarg_125_read,
    //input AXI-Stream to FIFO interface 126
    input s_axis_fifo_126_aclk,
    input s_axis_fifo_126_aresetn,
    input s_axis_fifo_126_tlast,
    input s_axis_fifo_126_tvalid,
    input [S_AXIS_FIFO_126_DMWIDTH/8-1:0] s_axis_fifo_126_tkeep,
    input [S_AXIS_FIFO_126_DMWIDTH/8-1:0] s_axis_fifo_126_tstrb,
    input [S_AXIS_FIFO_126_DMWIDTH-1:0] s_axis_fifo_126_tdata,
    output s_axis_fifo_126_tready,
    output ap_fifo_iarg_126_empty_n,
    output [S_AXIS_FIFO_126_WIDTH-1:0] ap_fifo_iarg_126_dout,
    input ap_fifo_iarg_126_read,
    //input AXI-Stream to FIFO interface 127
    input s_axis_fifo_127_aclk,
    input s_axis_fifo_127_aresetn,
    input s_axis_fifo_127_tlast,
    input s_axis_fifo_127_tvalid,
    input [S_AXIS_FIFO_127_DMWIDTH/8-1:0] s_axis_fifo_127_tkeep,
    input [S_AXIS_FIFO_127_DMWIDTH/8-1:0] s_axis_fifo_127_tstrb,
    input [S_AXIS_FIFO_127_DMWIDTH-1:0] s_axis_fifo_127_tdata,
    output s_axis_fifo_127_tready,
    output ap_fifo_iarg_127_empty_n,
    output [S_AXIS_FIFO_127_WIDTH-1:0] ap_fifo_iarg_127_dout,
    input ap_fifo_iarg_127_read,
    //-----------------------------------------------------
    //output FIFO to AXI-Stream interface 0
    input m_axis_fifo_0_aclk,
    input m_axis_fifo_0_aresetn,
    output m_axis_fifo_0_tlast,
    output m_axis_fifo_0_tvalid,
    output [M_AXIS_FIFO_0_DMWIDTH/8-1:0] m_axis_fifo_0_tkeep,
    output [M_AXIS_FIFO_0_DMWIDTH/8-1:0] m_axis_fifo_0_tstrb,
    output [M_AXIS_FIFO_0_DMWIDTH-1:0] m_axis_fifo_0_tdata,
    input m_axis_fifo_0_tready,
    output ap_fifo_oarg_0_full_n,
    input [M_AXIS_FIFO_0_WIDTH-1:0] ap_fifo_oarg_0_din,
    input ap_fifo_oarg_0_write,
    //output FIFO to AXI-Stream interface 1
    input m_axis_fifo_1_aclk,
    input m_axis_fifo_1_aresetn,
    output m_axis_fifo_1_tlast,
    output m_axis_fifo_1_tvalid,
    output [M_AXIS_FIFO_1_DMWIDTH/8-1:0] m_axis_fifo_1_tkeep,
    output [M_AXIS_FIFO_1_DMWIDTH/8-1:0] m_axis_fifo_1_tstrb,
    output [M_AXIS_FIFO_1_DMWIDTH-1:0] m_axis_fifo_1_tdata,
    input m_axis_fifo_1_tready,
    output ap_fifo_oarg_1_full_n,
    input [M_AXIS_FIFO_1_WIDTH-1:0] ap_fifo_oarg_1_din,
    input ap_fifo_oarg_1_write,
    //output FIFO to AXI-Stream interface 2
    input m_axis_fifo_2_aclk,
    input m_axis_fifo_2_aresetn,
    output m_axis_fifo_2_tlast,
    output m_axis_fifo_2_tvalid,
    output [M_AXIS_FIFO_2_DMWIDTH/8-1:0] m_axis_fifo_2_tkeep,
    output [M_AXIS_FIFO_2_DMWIDTH/8-1:0] m_axis_fifo_2_tstrb,
    output [M_AXIS_FIFO_2_DMWIDTH-1:0] m_axis_fifo_2_tdata,
    input m_axis_fifo_2_tready,
    output ap_fifo_oarg_2_full_n,
    input [M_AXIS_FIFO_2_WIDTH-1:0] ap_fifo_oarg_2_din,
    input ap_fifo_oarg_2_write,
    //output FIFO to AXI-Stream interface 3
    input m_axis_fifo_3_aclk,
    input m_axis_fifo_3_aresetn,
    output m_axis_fifo_3_tlast,
    output m_axis_fifo_3_tvalid,
    output [M_AXIS_FIFO_3_DMWIDTH/8-1:0] m_axis_fifo_3_tkeep,
    output [M_AXIS_FIFO_3_DMWIDTH/8-1:0] m_axis_fifo_3_tstrb,
    output [M_AXIS_FIFO_3_DMWIDTH-1:0] m_axis_fifo_3_tdata,
    input m_axis_fifo_3_tready,
    output ap_fifo_oarg_3_full_n,
    input [M_AXIS_FIFO_3_WIDTH-1:0] ap_fifo_oarg_3_din,
    input ap_fifo_oarg_3_write,
    //output FIFO to AXI-Stream interface 4
    input m_axis_fifo_4_aclk,
    input m_axis_fifo_4_aresetn,
    output m_axis_fifo_4_tlast,
    output m_axis_fifo_4_tvalid,
    output [M_AXIS_FIFO_4_DMWIDTH/8-1:0] m_axis_fifo_4_tkeep,
    output [M_AXIS_FIFO_4_DMWIDTH/8-1:0] m_axis_fifo_4_tstrb,
    output [M_AXIS_FIFO_4_DMWIDTH-1:0] m_axis_fifo_4_tdata,
    input m_axis_fifo_4_tready,
    output ap_fifo_oarg_4_full_n,
    input [M_AXIS_FIFO_4_WIDTH-1:0] ap_fifo_oarg_4_din,
    input ap_fifo_oarg_4_write,
    //output FIFO to AXI-Stream interface 5
    input m_axis_fifo_5_aclk,
    input m_axis_fifo_5_aresetn,
    output m_axis_fifo_5_tlast,
    output m_axis_fifo_5_tvalid,
    output [M_AXIS_FIFO_5_DMWIDTH/8-1:0] m_axis_fifo_5_tkeep,
    output [M_AXIS_FIFO_5_DMWIDTH/8-1:0] m_axis_fifo_5_tstrb,
    output [M_AXIS_FIFO_5_DMWIDTH-1:0] m_axis_fifo_5_tdata,
    input m_axis_fifo_5_tready,
    output ap_fifo_oarg_5_full_n,
    input [M_AXIS_FIFO_5_WIDTH-1:0] ap_fifo_oarg_5_din,
    input ap_fifo_oarg_5_write,
    //output FIFO to AXI-Stream interface 6
    input m_axis_fifo_6_aclk,
    input m_axis_fifo_6_aresetn,
    output m_axis_fifo_6_tlast,
    output m_axis_fifo_6_tvalid,
    output [M_AXIS_FIFO_6_DMWIDTH/8-1:0] m_axis_fifo_6_tkeep,
    output [M_AXIS_FIFO_6_DMWIDTH/8-1:0] m_axis_fifo_6_tstrb,
    output [M_AXIS_FIFO_6_DMWIDTH-1:0] m_axis_fifo_6_tdata,
    input m_axis_fifo_6_tready,
    output ap_fifo_oarg_6_full_n,
    input [M_AXIS_FIFO_6_WIDTH-1:0] ap_fifo_oarg_6_din,
    input ap_fifo_oarg_6_write,
    //output FIFO to AXI-Stream interface 7
    input m_axis_fifo_7_aclk,
    input m_axis_fifo_7_aresetn,
    output m_axis_fifo_7_tlast,
    output m_axis_fifo_7_tvalid,
    output [M_AXIS_FIFO_7_DMWIDTH/8-1:0] m_axis_fifo_7_tkeep,
    output [M_AXIS_FIFO_7_DMWIDTH/8-1:0] m_axis_fifo_7_tstrb,
    output [M_AXIS_FIFO_7_DMWIDTH-1:0] m_axis_fifo_7_tdata,
    input m_axis_fifo_7_tready,
    output ap_fifo_oarg_7_full_n,
    input [M_AXIS_FIFO_7_WIDTH-1:0] ap_fifo_oarg_7_din,
    input ap_fifo_oarg_7_write,
    //output FIFO to AXI-Stream interface 8
    input m_axis_fifo_8_aclk,
    input m_axis_fifo_8_aresetn,
    output m_axis_fifo_8_tlast,
    output m_axis_fifo_8_tvalid,
    output [M_AXIS_FIFO_8_DMWIDTH/8-1:0] m_axis_fifo_8_tkeep,
    output [M_AXIS_FIFO_8_DMWIDTH/8-1:0] m_axis_fifo_8_tstrb,
    output [M_AXIS_FIFO_8_DMWIDTH-1:0] m_axis_fifo_8_tdata,
    input m_axis_fifo_8_tready,
    output ap_fifo_oarg_8_full_n,
    input [M_AXIS_FIFO_8_WIDTH-1:0] ap_fifo_oarg_8_din,
    input ap_fifo_oarg_8_write,
    //output FIFO to AXI-Stream interface 9
    input m_axis_fifo_9_aclk,
    input m_axis_fifo_9_aresetn,
    output m_axis_fifo_9_tlast,
    output m_axis_fifo_9_tvalid,
    output [M_AXIS_FIFO_9_DMWIDTH/8-1:0] m_axis_fifo_9_tkeep,
    output [M_AXIS_FIFO_9_DMWIDTH/8-1:0] m_axis_fifo_9_tstrb,
    output [M_AXIS_FIFO_9_DMWIDTH-1:0] m_axis_fifo_9_tdata,
    input m_axis_fifo_9_tready,
    output ap_fifo_oarg_9_full_n,
    input [M_AXIS_FIFO_9_WIDTH-1:0] ap_fifo_oarg_9_din,
    input ap_fifo_oarg_9_write,
    //output FIFO to AXI-Stream interface 10
    input m_axis_fifo_10_aclk,
    input m_axis_fifo_10_aresetn,
    output m_axis_fifo_10_tlast,
    output m_axis_fifo_10_tvalid,
    output [M_AXIS_FIFO_10_DMWIDTH/8-1:0] m_axis_fifo_10_tkeep,
    output [M_AXIS_FIFO_10_DMWIDTH/8-1:0] m_axis_fifo_10_tstrb,
    output [M_AXIS_FIFO_10_DMWIDTH-1:0] m_axis_fifo_10_tdata,
    input m_axis_fifo_10_tready,
    output ap_fifo_oarg_10_full_n,
    input [M_AXIS_FIFO_10_WIDTH-1:0] ap_fifo_oarg_10_din,
    input ap_fifo_oarg_10_write,
    //output FIFO to AXI-Stream interface 11
    input m_axis_fifo_11_aclk,
    input m_axis_fifo_11_aresetn,
    output m_axis_fifo_11_tlast,
    output m_axis_fifo_11_tvalid,
    output [M_AXIS_FIFO_11_DMWIDTH/8-1:0] m_axis_fifo_11_tkeep,
    output [M_AXIS_FIFO_11_DMWIDTH/8-1:0] m_axis_fifo_11_tstrb,
    output [M_AXIS_FIFO_11_DMWIDTH-1:0] m_axis_fifo_11_tdata,
    input m_axis_fifo_11_tready,
    output ap_fifo_oarg_11_full_n,
    input [M_AXIS_FIFO_11_WIDTH-1:0] ap_fifo_oarg_11_din,
    input ap_fifo_oarg_11_write,
    //output FIFO to AXI-Stream interface 12
    input m_axis_fifo_12_aclk,
    input m_axis_fifo_12_aresetn,
    output m_axis_fifo_12_tlast,
    output m_axis_fifo_12_tvalid,
    output [M_AXIS_FIFO_12_DMWIDTH/8-1:0] m_axis_fifo_12_tkeep,
    output [M_AXIS_FIFO_12_DMWIDTH/8-1:0] m_axis_fifo_12_tstrb,
    output [M_AXIS_FIFO_12_DMWIDTH-1:0] m_axis_fifo_12_tdata,
    input m_axis_fifo_12_tready,
    output ap_fifo_oarg_12_full_n,
    input [M_AXIS_FIFO_12_WIDTH-1:0] ap_fifo_oarg_12_din,
    input ap_fifo_oarg_12_write,
    //output FIFO to AXI-Stream interface 13
    input m_axis_fifo_13_aclk,
    input m_axis_fifo_13_aresetn,
    output m_axis_fifo_13_tlast,
    output m_axis_fifo_13_tvalid,
    output [M_AXIS_FIFO_13_DMWIDTH/8-1:0] m_axis_fifo_13_tkeep,
    output [M_AXIS_FIFO_13_DMWIDTH/8-1:0] m_axis_fifo_13_tstrb,
    output [M_AXIS_FIFO_13_DMWIDTH-1:0] m_axis_fifo_13_tdata,
    input m_axis_fifo_13_tready,
    output ap_fifo_oarg_13_full_n,
    input [M_AXIS_FIFO_13_WIDTH-1:0] ap_fifo_oarg_13_din,
    input ap_fifo_oarg_13_write,
    //output FIFO to AXI-Stream interface 14
    input m_axis_fifo_14_aclk,
    input m_axis_fifo_14_aresetn,
    output m_axis_fifo_14_tlast,
    output m_axis_fifo_14_tvalid,
    output [M_AXIS_FIFO_14_DMWIDTH/8-1:0] m_axis_fifo_14_tkeep,
    output [M_AXIS_FIFO_14_DMWIDTH/8-1:0] m_axis_fifo_14_tstrb,
    output [M_AXIS_FIFO_14_DMWIDTH-1:0] m_axis_fifo_14_tdata,
    input m_axis_fifo_14_tready,
    output ap_fifo_oarg_14_full_n,
    input [M_AXIS_FIFO_14_WIDTH-1:0] ap_fifo_oarg_14_din,
    input ap_fifo_oarg_14_write,
    //output FIFO to AXI-Stream interface 15
    input m_axis_fifo_15_aclk,
    input m_axis_fifo_15_aresetn,
    output m_axis_fifo_15_tlast,
    output m_axis_fifo_15_tvalid,
    output [M_AXIS_FIFO_15_DMWIDTH/8-1:0] m_axis_fifo_15_tkeep,
    output [M_AXIS_FIFO_15_DMWIDTH/8-1:0] m_axis_fifo_15_tstrb,
    output [M_AXIS_FIFO_15_DMWIDTH-1:0] m_axis_fifo_15_tdata,
    input m_axis_fifo_15_tready,
    output ap_fifo_oarg_15_full_n,
    input [M_AXIS_FIFO_15_WIDTH-1:0] ap_fifo_oarg_15_din,
    input ap_fifo_oarg_15_write,
    //output FIFO to AXI-Stream interface 16
    input m_axis_fifo_16_aclk,
    input m_axis_fifo_16_aresetn,
    output m_axis_fifo_16_tlast,
    output m_axis_fifo_16_tvalid,
    output [M_AXIS_FIFO_16_DMWIDTH/8-1:0] m_axis_fifo_16_tkeep,
    output [M_AXIS_FIFO_16_DMWIDTH/8-1:0] m_axis_fifo_16_tstrb,
    output [M_AXIS_FIFO_16_DMWIDTH-1:0] m_axis_fifo_16_tdata,
    input m_axis_fifo_16_tready,
    output ap_fifo_oarg_16_full_n,
    input [M_AXIS_FIFO_16_WIDTH-1:0] ap_fifo_oarg_16_din,
    input ap_fifo_oarg_16_write,
    //output FIFO to AXI-Stream interface 17
    input m_axis_fifo_17_aclk,
    input m_axis_fifo_17_aresetn,
    output m_axis_fifo_17_tlast,
    output m_axis_fifo_17_tvalid,
    output [M_AXIS_FIFO_17_DMWIDTH/8-1:0] m_axis_fifo_17_tkeep,
    output [M_AXIS_FIFO_17_DMWIDTH/8-1:0] m_axis_fifo_17_tstrb,
    output [M_AXIS_FIFO_17_DMWIDTH-1:0] m_axis_fifo_17_tdata,
    input m_axis_fifo_17_tready,
    output ap_fifo_oarg_17_full_n,
    input [M_AXIS_FIFO_17_WIDTH-1:0] ap_fifo_oarg_17_din,
    input ap_fifo_oarg_17_write,
    //output FIFO to AXI-Stream interface 18
    input m_axis_fifo_18_aclk,
    input m_axis_fifo_18_aresetn,
    output m_axis_fifo_18_tlast,
    output m_axis_fifo_18_tvalid,
    output [M_AXIS_FIFO_18_DMWIDTH/8-1:0] m_axis_fifo_18_tkeep,
    output [M_AXIS_FIFO_18_DMWIDTH/8-1:0] m_axis_fifo_18_tstrb,
    output [M_AXIS_FIFO_18_DMWIDTH-1:0] m_axis_fifo_18_tdata,
    input m_axis_fifo_18_tready,
    output ap_fifo_oarg_18_full_n,
    input [M_AXIS_FIFO_18_WIDTH-1:0] ap_fifo_oarg_18_din,
    input ap_fifo_oarg_18_write,
    //output FIFO to AXI-Stream interface 19
    input m_axis_fifo_19_aclk,
    input m_axis_fifo_19_aresetn,
    output m_axis_fifo_19_tlast,
    output m_axis_fifo_19_tvalid,
    output [M_AXIS_FIFO_19_DMWIDTH/8-1:0] m_axis_fifo_19_tkeep,
    output [M_AXIS_FIFO_19_DMWIDTH/8-1:0] m_axis_fifo_19_tstrb,
    output [M_AXIS_FIFO_19_DMWIDTH-1:0] m_axis_fifo_19_tdata,
    input m_axis_fifo_19_tready,
    output ap_fifo_oarg_19_full_n,
    input [M_AXIS_FIFO_19_WIDTH-1:0] ap_fifo_oarg_19_din,
    input ap_fifo_oarg_19_write,
    //output FIFO to AXI-Stream interface 20
    input m_axis_fifo_20_aclk,
    input m_axis_fifo_20_aresetn,
    output m_axis_fifo_20_tlast,
    output m_axis_fifo_20_tvalid,
    output [M_AXIS_FIFO_20_DMWIDTH/8-1:0] m_axis_fifo_20_tkeep,
    output [M_AXIS_FIFO_20_DMWIDTH/8-1:0] m_axis_fifo_20_tstrb,
    output [M_AXIS_FIFO_20_DMWIDTH-1:0] m_axis_fifo_20_tdata,
    input m_axis_fifo_20_tready,
    output ap_fifo_oarg_20_full_n,
    input [M_AXIS_FIFO_20_WIDTH-1:0] ap_fifo_oarg_20_din,
    input ap_fifo_oarg_20_write,
    //output FIFO to AXI-Stream interface 21
    input m_axis_fifo_21_aclk,
    input m_axis_fifo_21_aresetn,
    output m_axis_fifo_21_tlast,
    output m_axis_fifo_21_tvalid,
    output [M_AXIS_FIFO_21_DMWIDTH/8-1:0] m_axis_fifo_21_tkeep,
    output [M_AXIS_FIFO_21_DMWIDTH/8-1:0] m_axis_fifo_21_tstrb,
    output [M_AXIS_FIFO_21_DMWIDTH-1:0] m_axis_fifo_21_tdata,
    input m_axis_fifo_21_tready,
    output ap_fifo_oarg_21_full_n,
    input [M_AXIS_FIFO_21_WIDTH-1:0] ap_fifo_oarg_21_din,
    input ap_fifo_oarg_21_write,
    //output FIFO to AXI-Stream interface 22
    input m_axis_fifo_22_aclk,
    input m_axis_fifo_22_aresetn,
    output m_axis_fifo_22_tlast,
    output m_axis_fifo_22_tvalid,
    output [M_AXIS_FIFO_22_DMWIDTH/8-1:0] m_axis_fifo_22_tkeep,
    output [M_AXIS_FIFO_22_DMWIDTH/8-1:0] m_axis_fifo_22_tstrb,
    output [M_AXIS_FIFO_22_DMWIDTH-1:0] m_axis_fifo_22_tdata,
    input m_axis_fifo_22_tready,
    output ap_fifo_oarg_22_full_n,
    input [M_AXIS_FIFO_22_WIDTH-1:0] ap_fifo_oarg_22_din,
    input ap_fifo_oarg_22_write,
    //output FIFO to AXI-Stream interface 23
    input m_axis_fifo_23_aclk,
    input m_axis_fifo_23_aresetn,
    output m_axis_fifo_23_tlast,
    output m_axis_fifo_23_tvalid,
    output [M_AXIS_FIFO_23_DMWIDTH/8-1:0] m_axis_fifo_23_tkeep,
    output [M_AXIS_FIFO_23_DMWIDTH/8-1:0] m_axis_fifo_23_tstrb,
    output [M_AXIS_FIFO_23_DMWIDTH-1:0] m_axis_fifo_23_tdata,
    input m_axis_fifo_23_tready,
    output ap_fifo_oarg_23_full_n,
    input [M_AXIS_FIFO_23_WIDTH-1:0] ap_fifo_oarg_23_din,
    input ap_fifo_oarg_23_write,
    //output FIFO to AXI-Stream interface 24
    input m_axis_fifo_24_aclk,
    input m_axis_fifo_24_aresetn,
    output m_axis_fifo_24_tlast,
    output m_axis_fifo_24_tvalid,
    output [M_AXIS_FIFO_24_DMWIDTH/8-1:0] m_axis_fifo_24_tkeep,
    output [M_AXIS_FIFO_24_DMWIDTH/8-1:0] m_axis_fifo_24_tstrb,
    output [M_AXIS_FIFO_24_DMWIDTH-1:0] m_axis_fifo_24_tdata,
    input m_axis_fifo_24_tready,
    output ap_fifo_oarg_24_full_n,
    input [M_AXIS_FIFO_24_WIDTH-1:0] ap_fifo_oarg_24_din,
    input ap_fifo_oarg_24_write,
    //output FIFO to AXI-Stream interface 25
    input m_axis_fifo_25_aclk,
    input m_axis_fifo_25_aresetn,
    output m_axis_fifo_25_tlast,
    output m_axis_fifo_25_tvalid,
    output [M_AXIS_FIFO_25_DMWIDTH/8-1:0] m_axis_fifo_25_tkeep,
    output [M_AXIS_FIFO_25_DMWIDTH/8-1:0] m_axis_fifo_25_tstrb,
    output [M_AXIS_FIFO_25_DMWIDTH-1:0] m_axis_fifo_25_tdata,
    input m_axis_fifo_25_tready,
    output ap_fifo_oarg_25_full_n,
    input [M_AXIS_FIFO_25_WIDTH-1:0] ap_fifo_oarg_25_din,
    input ap_fifo_oarg_25_write,
    //output FIFO to AXI-Stream interface 26
    input m_axis_fifo_26_aclk,
    input m_axis_fifo_26_aresetn,
    output m_axis_fifo_26_tlast,
    output m_axis_fifo_26_tvalid,
    output [M_AXIS_FIFO_26_DMWIDTH/8-1:0] m_axis_fifo_26_tkeep,
    output [M_AXIS_FIFO_26_DMWIDTH/8-1:0] m_axis_fifo_26_tstrb,
    output [M_AXIS_FIFO_26_DMWIDTH-1:0] m_axis_fifo_26_tdata,
    input m_axis_fifo_26_tready,
    output ap_fifo_oarg_26_full_n,
    input [M_AXIS_FIFO_26_WIDTH-1:0] ap_fifo_oarg_26_din,
    input ap_fifo_oarg_26_write,
    //output FIFO to AXI-Stream interface 27
    input m_axis_fifo_27_aclk,
    input m_axis_fifo_27_aresetn,
    output m_axis_fifo_27_tlast,
    output m_axis_fifo_27_tvalid,
    output [M_AXIS_FIFO_27_DMWIDTH/8-1:0] m_axis_fifo_27_tkeep,
    output [M_AXIS_FIFO_27_DMWIDTH/8-1:0] m_axis_fifo_27_tstrb,
    output [M_AXIS_FIFO_27_DMWIDTH-1:0] m_axis_fifo_27_tdata,
    input m_axis_fifo_27_tready,
    output ap_fifo_oarg_27_full_n,
    input [M_AXIS_FIFO_27_WIDTH-1:0] ap_fifo_oarg_27_din,
    input ap_fifo_oarg_27_write,
    //output FIFO to AXI-Stream interface 28
    input m_axis_fifo_28_aclk,
    input m_axis_fifo_28_aresetn,
    output m_axis_fifo_28_tlast,
    output m_axis_fifo_28_tvalid,
    output [M_AXIS_FIFO_28_DMWIDTH/8-1:0] m_axis_fifo_28_tkeep,
    output [M_AXIS_FIFO_28_DMWIDTH/8-1:0] m_axis_fifo_28_tstrb,
    output [M_AXIS_FIFO_28_DMWIDTH-1:0] m_axis_fifo_28_tdata,
    input m_axis_fifo_28_tready,
    output ap_fifo_oarg_28_full_n,
    input [M_AXIS_FIFO_28_WIDTH-1:0] ap_fifo_oarg_28_din,
    input ap_fifo_oarg_28_write,
    //output FIFO to AXI-Stream interface 29
    input m_axis_fifo_29_aclk,
    input m_axis_fifo_29_aresetn,
    output m_axis_fifo_29_tlast,
    output m_axis_fifo_29_tvalid,
    output [M_AXIS_FIFO_29_DMWIDTH/8-1:0] m_axis_fifo_29_tkeep,
    output [M_AXIS_FIFO_29_DMWIDTH/8-1:0] m_axis_fifo_29_tstrb,
    output [M_AXIS_FIFO_29_DMWIDTH-1:0] m_axis_fifo_29_tdata,
    input m_axis_fifo_29_tready,
    output ap_fifo_oarg_29_full_n,
    input [M_AXIS_FIFO_29_WIDTH-1:0] ap_fifo_oarg_29_din,
    input ap_fifo_oarg_29_write,
    //output FIFO to AXI-Stream interface 30
    input m_axis_fifo_30_aclk,
    input m_axis_fifo_30_aresetn,
    output m_axis_fifo_30_tlast,
    output m_axis_fifo_30_tvalid,
    output [M_AXIS_FIFO_30_DMWIDTH/8-1:0] m_axis_fifo_30_tkeep,
    output [M_AXIS_FIFO_30_DMWIDTH/8-1:0] m_axis_fifo_30_tstrb,
    output [M_AXIS_FIFO_30_DMWIDTH-1:0] m_axis_fifo_30_tdata,
    input m_axis_fifo_30_tready,
    output ap_fifo_oarg_30_full_n,
    input [M_AXIS_FIFO_30_WIDTH-1:0] ap_fifo_oarg_30_din,
    input ap_fifo_oarg_30_write,
    //output FIFO to AXI-Stream interface 31
    input m_axis_fifo_31_aclk,
    input m_axis_fifo_31_aresetn,
    output m_axis_fifo_31_tlast,
    output m_axis_fifo_31_tvalid,
    output [M_AXIS_FIFO_31_DMWIDTH/8-1:0] m_axis_fifo_31_tkeep,
    output [M_AXIS_FIFO_31_DMWIDTH/8-1:0] m_axis_fifo_31_tstrb,
    output [M_AXIS_FIFO_31_DMWIDTH-1:0] m_axis_fifo_31_tdata,
    input m_axis_fifo_31_tready,
    output ap_fifo_oarg_31_full_n,
    input [M_AXIS_FIFO_31_WIDTH-1:0] ap_fifo_oarg_31_din,
    input ap_fifo_oarg_31_write,
    //output FIFO to AXI-Stream interface 32
    input m_axis_fifo_32_aclk,
    input m_axis_fifo_32_aresetn,
    output m_axis_fifo_32_tlast,
    output m_axis_fifo_32_tvalid,
    output [M_AXIS_FIFO_32_DMWIDTH/8-1:0] m_axis_fifo_32_tkeep,
    output [M_AXIS_FIFO_32_DMWIDTH/8-1:0] m_axis_fifo_32_tstrb,
    output [M_AXIS_FIFO_32_DMWIDTH-1:0] m_axis_fifo_32_tdata,
    input m_axis_fifo_32_tready,
    output ap_fifo_oarg_32_full_n,
    input [M_AXIS_FIFO_32_WIDTH-1:0] ap_fifo_oarg_32_din,
    input ap_fifo_oarg_32_write,
    //output FIFO to AXI-Stream interface 33
    input m_axis_fifo_33_aclk,
    input m_axis_fifo_33_aresetn,
    output m_axis_fifo_33_tlast,
    output m_axis_fifo_33_tvalid,
    output [M_AXIS_FIFO_33_DMWIDTH/8-1:0] m_axis_fifo_33_tkeep,
    output [M_AXIS_FIFO_33_DMWIDTH/8-1:0] m_axis_fifo_33_tstrb,
    output [M_AXIS_FIFO_33_DMWIDTH-1:0] m_axis_fifo_33_tdata,
    input m_axis_fifo_33_tready,
    output ap_fifo_oarg_33_full_n,
    input [M_AXIS_FIFO_33_WIDTH-1:0] ap_fifo_oarg_33_din,
    input ap_fifo_oarg_33_write,
    //output FIFO to AXI-Stream interface 34
    input m_axis_fifo_34_aclk,
    input m_axis_fifo_34_aresetn,
    output m_axis_fifo_34_tlast,
    output m_axis_fifo_34_tvalid,
    output [M_AXIS_FIFO_34_DMWIDTH/8-1:0] m_axis_fifo_34_tkeep,
    output [M_AXIS_FIFO_34_DMWIDTH/8-1:0] m_axis_fifo_34_tstrb,
    output [M_AXIS_FIFO_34_DMWIDTH-1:0] m_axis_fifo_34_tdata,
    input m_axis_fifo_34_tready,
    output ap_fifo_oarg_34_full_n,
    input [M_AXIS_FIFO_34_WIDTH-1:0] ap_fifo_oarg_34_din,
    input ap_fifo_oarg_34_write,
    //output FIFO to AXI-Stream interface 35
    input m_axis_fifo_35_aclk,
    input m_axis_fifo_35_aresetn,
    output m_axis_fifo_35_tlast,
    output m_axis_fifo_35_tvalid,
    output [M_AXIS_FIFO_35_DMWIDTH/8-1:0] m_axis_fifo_35_tkeep,
    output [M_AXIS_FIFO_35_DMWIDTH/8-1:0] m_axis_fifo_35_tstrb,
    output [M_AXIS_FIFO_35_DMWIDTH-1:0] m_axis_fifo_35_tdata,
    input m_axis_fifo_35_tready,
    output ap_fifo_oarg_35_full_n,
    input [M_AXIS_FIFO_35_WIDTH-1:0] ap_fifo_oarg_35_din,
    input ap_fifo_oarg_35_write,
    //output FIFO to AXI-Stream interface 36
    input m_axis_fifo_36_aclk,
    input m_axis_fifo_36_aresetn,
    output m_axis_fifo_36_tlast,
    output m_axis_fifo_36_tvalid,
    output [M_AXIS_FIFO_36_DMWIDTH/8-1:0] m_axis_fifo_36_tkeep,
    output [M_AXIS_FIFO_36_DMWIDTH/8-1:0] m_axis_fifo_36_tstrb,
    output [M_AXIS_FIFO_36_DMWIDTH-1:0] m_axis_fifo_36_tdata,
    input m_axis_fifo_36_tready,
    output ap_fifo_oarg_36_full_n,
    input [M_AXIS_FIFO_36_WIDTH-1:0] ap_fifo_oarg_36_din,
    input ap_fifo_oarg_36_write,
    //output FIFO to AXI-Stream interface 37
    input m_axis_fifo_37_aclk,
    input m_axis_fifo_37_aresetn,
    output m_axis_fifo_37_tlast,
    output m_axis_fifo_37_tvalid,
    output [M_AXIS_FIFO_37_DMWIDTH/8-1:0] m_axis_fifo_37_tkeep,
    output [M_AXIS_FIFO_37_DMWIDTH/8-1:0] m_axis_fifo_37_tstrb,
    output [M_AXIS_FIFO_37_DMWIDTH-1:0] m_axis_fifo_37_tdata,
    input m_axis_fifo_37_tready,
    output ap_fifo_oarg_37_full_n,
    input [M_AXIS_FIFO_37_WIDTH-1:0] ap_fifo_oarg_37_din,
    input ap_fifo_oarg_37_write,
    //output FIFO to AXI-Stream interface 38
    input m_axis_fifo_38_aclk,
    input m_axis_fifo_38_aresetn,
    output m_axis_fifo_38_tlast,
    output m_axis_fifo_38_tvalid,
    output [M_AXIS_FIFO_38_DMWIDTH/8-1:0] m_axis_fifo_38_tkeep,
    output [M_AXIS_FIFO_38_DMWIDTH/8-1:0] m_axis_fifo_38_tstrb,
    output [M_AXIS_FIFO_38_DMWIDTH-1:0] m_axis_fifo_38_tdata,
    input m_axis_fifo_38_tready,
    output ap_fifo_oarg_38_full_n,
    input [M_AXIS_FIFO_38_WIDTH-1:0] ap_fifo_oarg_38_din,
    input ap_fifo_oarg_38_write,
    //output FIFO to AXI-Stream interface 39
    input m_axis_fifo_39_aclk,
    input m_axis_fifo_39_aresetn,
    output m_axis_fifo_39_tlast,
    output m_axis_fifo_39_tvalid,
    output [M_AXIS_FIFO_39_DMWIDTH/8-1:0] m_axis_fifo_39_tkeep,
    output [M_AXIS_FIFO_39_DMWIDTH/8-1:0] m_axis_fifo_39_tstrb,
    output [M_AXIS_FIFO_39_DMWIDTH-1:0] m_axis_fifo_39_tdata,
    input m_axis_fifo_39_tready,
    output ap_fifo_oarg_39_full_n,
    input [M_AXIS_FIFO_39_WIDTH-1:0] ap_fifo_oarg_39_din,
    input ap_fifo_oarg_39_write,
    //output FIFO to AXI-Stream interface 40
    input m_axis_fifo_40_aclk,
    input m_axis_fifo_40_aresetn,
    output m_axis_fifo_40_tlast,
    output m_axis_fifo_40_tvalid,
    output [M_AXIS_FIFO_40_DMWIDTH/8-1:0] m_axis_fifo_40_tkeep,
    output [M_AXIS_FIFO_40_DMWIDTH/8-1:0] m_axis_fifo_40_tstrb,
    output [M_AXIS_FIFO_40_DMWIDTH-1:0] m_axis_fifo_40_tdata,
    input m_axis_fifo_40_tready,
    output ap_fifo_oarg_40_full_n,
    input [M_AXIS_FIFO_40_WIDTH-1:0] ap_fifo_oarg_40_din,
    input ap_fifo_oarg_40_write,
    //output FIFO to AXI-Stream interface 41
    input m_axis_fifo_41_aclk,
    input m_axis_fifo_41_aresetn,
    output m_axis_fifo_41_tlast,
    output m_axis_fifo_41_tvalid,
    output [M_AXIS_FIFO_41_DMWIDTH/8-1:0] m_axis_fifo_41_tkeep,
    output [M_AXIS_FIFO_41_DMWIDTH/8-1:0] m_axis_fifo_41_tstrb,
    output [M_AXIS_FIFO_41_DMWIDTH-1:0] m_axis_fifo_41_tdata,
    input m_axis_fifo_41_tready,
    output ap_fifo_oarg_41_full_n,
    input [M_AXIS_FIFO_41_WIDTH-1:0] ap_fifo_oarg_41_din,
    input ap_fifo_oarg_41_write,
    //output FIFO to AXI-Stream interface 42
    input m_axis_fifo_42_aclk,
    input m_axis_fifo_42_aresetn,
    output m_axis_fifo_42_tlast,
    output m_axis_fifo_42_tvalid,
    output [M_AXIS_FIFO_42_DMWIDTH/8-1:0] m_axis_fifo_42_tkeep,
    output [M_AXIS_FIFO_42_DMWIDTH/8-1:0] m_axis_fifo_42_tstrb,
    output [M_AXIS_FIFO_42_DMWIDTH-1:0] m_axis_fifo_42_tdata,
    input m_axis_fifo_42_tready,
    output ap_fifo_oarg_42_full_n,
    input [M_AXIS_FIFO_42_WIDTH-1:0] ap_fifo_oarg_42_din,
    input ap_fifo_oarg_42_write,
    //output FIFO to AXI-Stream interface 43
    input m_axis_fifo_43_aclk,
    input m_axis_fifo_43_aresetn,
    output m_axis_fifo_43_tlast,
    output m_axis_fifo_43_tvalid,
    output [M_AXIS_FIFO_43_DMWIDTH/8-1:0] m_axis_fifo_43_tkeep,
    output [M_AXIS_FIFO_43_DMWIDTH/8-1:0] m_axis_fifo_43_tstrb,
    output [M_AXIS_FIFO_43_DMWIDTH-1:0] m_axis_fifo_43_tdata,
    input m_axis_fifo_43_tready,
    output ap_fifo_oarg_43_full_n,
    input [M_AXIS_FIFO_43_WIDTH-1:0] ap_fifo_oarg_43_din,
    input ap_fifo_oarg_43_write,
    //output FIFO to AXI-Stream interface 44
    input m_axis_fifo_44_aclk,
    input m_axis_fifo_44_aresetn,
    output m_axis_fifo_44_tlast,
    output m_axis_fifo_44_tvalid,
    output [M_AXIS_FIFO_44_DMWIDTH/8-1:0] m_axis_fifo_44_tkeep,
    output [M_AXIS_FIFO_44_DMWIDTH/8-1:0] m_axis_fifo_44_tstrb,
    output [M_AXIS_FIFO_44_DMWIDTH-1:0] m_axis_fifo_44_tdata,
    input m_axis_fifo_44_tready,
    output ap_fifo_oarg_44_full_n,
    input [M_AXIS_FIFO_44_WIDTH-1:0] ap_fifo_oarg_44_din,
    input ap_fifo_oarg_44_write,
    //output FIFO to AXI-Stream interface 45
    input m_axis_fifo_45_aclk,
    input m_axis_fifo_45_aresetn,
    output m_axis_fifo_45_tlast,
    output m_axis_fifo_45_tvalid,
    output [M_AXIS_FIFO_45_DMWIDTH/8-1:0] m_axis_fifo_45_tkeep,
    output [M_AXIS_FIFO_45_DMWIDTH/8-1:0] m_axis_fifo_45_tstrb,
    output [M_AXIS_FIFO_45_DMWIDTH-1:0] m_axis_fifo_45_tdata,
    input m_axis_fifo_45_tready,
    output ap_fifo_oarg_45_full_n,
    input [M_AXIS_FIFO_45_WIDTH-1:0] ap_fifo_oarg_45_din,
    input ap_fifo_oarg_45_write,
    //output FIFO to AXI-Stream interface 46
    input m_axis_fifo_46_aclk,
    input m_axis_fifo_46_aresetn,
    output m_axis_fifo_46_tlast,
    output m_axis_fifo_46_tvalid,
    output [M_AXIS_FIFO_46_DMWIDTH/8-1:0] m_axis_fifo_46_tkeep,
    output [M_AXIS_FIFO_46_DMWIDTH/8-1:0] m_axis_fifo_46_tstrb,
    output [M_AXIS_FIFO_46_DMWIDTH-1:0] m_axis_fifo_46_tdata,
    input m_axis_fifo_46_tready,
    output ap_fifo_oarg_46_full_n,
    input [M_AXIS_FIFO_46_WIDTH-1:0] ap_fifo_oarg_46_din,
    input ap_fifo_oarg_46_write,
    //output FIFO to AXI-Stream interface 47
    input m_axis_fifo_47_aclk,
    input m_axis_fifo_47_aresetn,
    output m_axis_fifo_47_tlast,
    output m_axis_fifo_47_tvalid,
    output [M_AXIS_FIFO_47_DMWIDTH/8-1:0] m_axis_fifo_47_tkeep,
    output [M_AXIS_FIFO_47_DMWIDTH/8-1:0] m_axis_fifo_47_tstrb,
    output [M_AXIS_FIFO_47_DMWIDTH-1:0] m_axis_fifo_47_tdata,
    input m_axis_fifo_47_tready,
    output ap_fifo_oarg_47_full_n,
    input [M_AXIS_FIFO_47_WIDTH-1:0] ap_fifo_oarg_47_din,
    input ap_fifo_oarg_47_write,
    //output FIFO to AXI-Stream interface 48
    input m_axis_fifo_48_aclk,
    input m_axis_fifo_48_aresetn,
    output m_axis_fifo_48_tlast,
    output m_axis_fifo_48_tvalid,
    output [M_AXIS_FIFO_48_DMWIDTH/8-1:0] m_axis_fifo_48_tkeep,
    output [M_AXIS_FIFO_48_DMWIDTH/8-1:0] m_axis_fifo_48_tstrb,
    output [M_AXIS_FIFO_48_DMWIDTH-1:0] m_axis_fifo_48_tdata,
    input m_axis_fifo_48_tready,
    output ap_fifo_oarg_48_full_n,
    input [M_AXIS_FIFO_48_WIDTH-1:0] ap_fifo_oarg_48_din,
    input ap_fifo_oarg_48_write,
    //output FIFO to AXI-Stream interface 49
    input m_axis_fifo_49_aclk,
    input m_axis_fifo_49_aresetn,
    output m_axis_fifo_49_tlast,
    output m_axis_fifo_49_tvalid,
    output [M_AXIS_FIFO_49_DMWIDTH/8-1:0] m_axis_fifo_49_tkeep,
    output [M_AXIS_FIFO_49_DMWIDTH/8-1:0] m_axis_fifo_49_tstrb,
    output [M_AXIS_FIFO_49_DMWIDTH-1:0] m_axis_fifo_49_tdata,
    input m_axis_fifo_49_tready,
    output ap_fifo_oarg_49_full_n,
    input [M_AXIS_FIFO_49_WIDTH-1:0] ap_fifo_oarg_49_din,
    input ap_fifo_oarg_49_write,
    //output FIFO to AXI-Stream interface 50
    input m_axis_fifo_50_aclk,
    input m_axis_fifo_50_aresetn,
    output m_axis_fifo_50_tlast,
    output m_axis_fifo_50_tvalid,
    output [M_AXIS_FIFO_50_DMWIDTH/8-1:0] m_axis_fifo_50_tkeep,
    output [M_AXIS_FIFO_50_DMWIDTH/8-1:0] m_axis_fifo_50_tstrb,
    output [M_AXIS_FIFO_50_DMWIDTH-1:0] m_axis_fifo_50_tdata,
    input m_axis_fifo_50_tready,
    output ap_fifo_oarg_50_full_n,
    input [M_AXIS_FIFO_50_WIDTH-1:0] ap_fifo_oarg_50_din,
    input ap_fifo_oarg_50_write,
    //output FIFO to AXI-Stream interface 51
    input m_axis_fifo_51_aclk,
    input m_axis_fifo_51_aresetn,
    output m_axis_fifo_51_tlast,
    output m_axis_fifo_51_tvalid,
    output [M_AXIS_FIFO_51_DMWIDTH/8-1:0] m_axis_fifo_51_tkeep,
    output [M_AXIS_FIFO_51_DMWIDTH/8-1:0] m_axis_fifo_51_tstrb,
    output [M_AXIS_FIFO_51_DMWIDTH-1:0] m_axis_fifo_51_tdata,
    input m_axis_fifo_51_tready,
    output ap_fifo_oarg_51_full_n,
    input [M_AXIS_FIFO_51_WIDTH-1:0] ap_fifo_oarg_51_din,
    input ap_fifo_oarg_51_write,
    //output FIFO to AXI-Stream interface 52
    input m_axis_fifo_52_aclk,
    input m_axis_fifo_52_aresetn,
    output m_axis_fifo_52_tlast,
    output m_axis_fifo_52_tvalid,
    output [M_AXIS_FIFO_52_DMWIDTH/8-1:0] m_axis_fifo_52_tkeep,
    output [M_AXIS_FIFO_52_DMWIDTH/8-1:0] m_axis_fifo_52_tstrb,
    output [M_AXIS_FIFO_52_DMWIDTH-1:0] m_axis_fifo_52_tdata,
    input m_axis_fifo_52_tready,
    output ap_fifo_oarg_52_full_n,
    input [M_AXIS_FIFO_52_WIDTH-1:0] ap_fifo_oarg_52_din,
    input ap_fifo_oarg_52_write,
    //output FIFO to AXI-Stream interface 53
    input m_axis_fifo_53_aclk,
    input m_axis_fifo_53_aresetn,
    output m_axis_fifo_53_tlast,
    output m_axis_fifo_53_tvalid,
    output [M_AXIS_FIFO_53_DMWIDTH/8-1:0] m_axis_fifo_53_tkeep,
    output [M_AXIS_FIFO_53_DMWIDTH/8-1:0] m_axis_fifo_53_tstrb,
    output [M_AXIS_FIFO_53_DMWIDTH-1:0] m_axis_fifo_53_tdata,
    input m_axis_fifo_53_tready,
    output ap_fifo_oarg_53_full_n,
    input [M_AXIS_FIFO_53_WIDTH-1:0] ap_fifo_oarg_53_din,
    input ap_fifo_oarg_53_write,
    //output FIFO to AXI-Stream interface 54
    input m_axis_fifo_54_aclk,
    input m_axis_fifo_54_aresetn,
    output m_axis_fifo_54_tlast,
    output m_axis_fifo_54_tvalid,
    output [M_AXIS_FIFO_54_DMWIDTH/8-1:0] m_axis_fifo_54_tkeep,
    output [M_AXIS_FIFO_54_DMWIDTH/8-1:0] m_axis_fifo_54_tstrb,
    output [M_AXIS_FIFO_54_DMWIDTH-1:0] m_axis_fifo_54_tdata,
    input m_axis_fifo_54_tready,
    output ap_fifo_oarg_54_full_n,
    input [M_AXIS_FIFO_54_WIDTH-1:0] ap_fifo_oarg_54_din,
    input ap_fifo_oarg_54_write,
    //output FIFO to AXI-Stream interface 55
    input m_axis_fifo_55_aclk,
    input m_axis_fifo_55_aresetn,
    output m_axis_fifo_55_tlast,
    output m_axis_fifo_55_tvalid,
    output [M_AXIS_FIFO_55_DMWIDTH/8-1:0] m_axis_fifo_55_tkeep,
    output [M_AXIS_FIFO_55_DMWIDTH/8-1:0] m_axis_fifo_55_tstrb,
    output [M_AXIS_FIFO_55_DMWIDTH-1:0] m_axis_fifo_55_tdata,
    input m_axis_fifo_55_tready,
    output ap_fifo_oarg_55_full_n,
    input [M_AXIS_FIFO_55_WIDTH-1:0] ap_fifo_oarg_55_din,
    input ap_fifo_oarg_55_write,
    //output FIFO to AXI-Stream interface 56
    input m_axis_fifo_56_aclk,
    input m_axis_fifo_56_aresetn,
    output m_axis_fifo_56_tlast,
    output m_axis_fifo_56_tvalid,
    output [M_AXIS_FIFO_56_DMWIDTH/8-1:0] m_axis_fifo_56_tkeep,
    output [M_AXIS_FIFO_56_DMWIDTH/8-1:0] m_axis_fifo_56_tstrb,
    output [M_AXIS_FIFO_56_DMWIDTH-1:0] m_axis_fifo_56_tdata,
    input m_axis_fifo_56_tready,
    output ap_fifo_oarg_56_full_n,
    input [M_AXIS_FIFO_56_WIDTH-1:0] ap_fifo_oarg_56_din,
    input ap_fifo_oarg_56_write,
    //output FIFO to AXI-Stream interface 57
    input m_axis_fifo_57_aclk,
    input m_axis_fifo_57_aresetn,
    output m_axis_fifo_57_tlast,
    output m_axis_fifo_57_tvalid,
    output [M_AXIS_FIFO_57_DMWIDTH/8-1:0] m_axis_fifo_57_tkeep,
    output [M_AXIS_FIFO_57_DMWIDTH/8-1:0] m_axis_fifo_57_tstrb,
    output [M_AXIS_FIFO_57_DMWIDTH-1:0] m_axis_fifo_57_tdata,
    input m_axis_fifo_57_tready,
    output ap_fifo_oarg_57_full_n,
    input [M_AXIS_FIFO_57_WIDTH-1:0] ap_fifo_oarg_57_din,
    input ap_fifo_oarg_57_write,
    //output FIFO to AXI-Stream interface 58
    input m_axis_fifo_58_aclk,
    input m_axis_fifo_58_aresetn,
    output m_axis_fifo_58_tlast,
    output m_axis_fifo_58_tvalid,
    output [M_AXIS_FIFO_58_DMWIDTH/8-1:0] m_axis_fifo_58_tkeep,
    output [M_AXIS_FIFO_58_DMWIDTH/8-1:0] m_axis_fifo_58_tstrb,
    output [M_AXIS_FIFO_58_DMWIDTH-1:0] m_axis_fifo_58_tdata,
    input m_axis_fifo_58_tready,
    output ap_fifo_oarg_58_full_n,
    input [M_AXIS_FIFO_58_WIDTH-1:0] ap_fifo_oarg_58_din,
    input ap_fifo_oarg_58_write,
    //output FIFO to AXI-Stream interface 59
    input m_axis_fifo_59_aclk,
    input m_axis_fifo_59_aresetn,
    output m_axis_fifo_59_tlast,
    output m_axis_fifo_59_tvalid,
    output [M_AXIS_FIFO_59_DMWIDTH/8-1:0] m_axis_fifo_59_tkeep,
    output [M_AXIS_FIFO_59_DMWIDTH/8-1:0] m_axis_fifo_59_tstrb,
    output [M_AXIS_FIFO_59_DMWIDTH-1:0] m_axis_fifo_59_tdata,
    input m_axis_fifo_59_tready,
    output ap_fifo_oarg_59_full_n,
    input [M_AXIS_FIFO_59_WIDTH-1:0] ap_fifo_oarg_59_din,
    input ap_fifo_oarg_59_write,
    //output FIFO to AXI-Stream interface 60
    input m_axis_fifo_60_aclk,
    input m_axis_fifo_60_aresetn,
    output m_axis_fifo_60_tlast,
    output m_axis_fifo_60_tvalid,
    output [M_AXIS_FIFO_60_DMWIDTH/8-1:0] m_axis_fifo_60_tkeep,
    output [M_AXIS_FIFO_60_DMWIDTH/8-1:0] m_axis_fifo_60_tstrb,
    output [M_AXIS_FIFO_60_DMWIDTH-1:0] m_axis_fifo_60_tdata,
    input m_axis_fifo_60_tready,
    output ap_fifo_oarg_60_full_n,
    input [M_AXIS_FIFO_60_WIDTH-1:0] ap_fifo_oarg_60_din,
    input ap_fifo_oarg_60_write,
    //output FIFO to AXI-Stream interface 61
    input m_axis_fifo_61_aclk,
    input m_axis_fifo_61_aresetn,
    output m_axis_fifo_61_tlast,
    output m_axis_fifo_61_tvalid,
    output [M_AXIS_FIFO_61_DMWIDTH/8-1:0] m_axis_fifo_61_tkeep,
    output [M_AXIS_FIFO_61_DMWIDTH/8-1:0] m_axis_fifo_61_tstrb,
    output [M_AXIS_FIFO_61_DMWIDTH-1:0] m_axis_fifo_61_tdata,
    input m_axis_fifo_61_tready,
    output ap_fifo_oarg_61_full_n,
    input [M_AXIS_FIFO_61_WIDTH-1:0] ap_fifo_oarg_61_din,
    input ap_fifo_oarg_61_write,
    //output FIFO to AXI-Stream interface 62
    input m_axis_fifo_62_aclk,
    input m_axis_fifo_62_aresetn,
    output m_axis_fifo_62_tlast,
    output m_axis_fifo_62_tvalid,
    output [M_AXIS_FIFO_62_DMWIDTH/8-1:0] m_axis_fifo_62_tkeep,
    output [M_AXIS_FIFO_62_DMWIDTH/8-1:0] m_axis_fifo_62_tstrb,
    output [M_AXIS_FIFO_62_DMWIDTH-1:0] m_axis_fifo_62_tdata,
    input m_axis_fifo_62_tready,
    output ap_fifo_oarg_62_full_n,
    input [M_AXIS_FIFO_62_WIDTH-1:0] ap_fifo_oarg_62_din,
    input ap_fifo_oarg_62_write,
    //output FIFO to AXI-Stream interface 63
    input m_axis_fifo_63_aclk,
    input m_axis_fifo_63_aresetn,
    output m_axis_fifo_63_tlast,
    output m_axis_fifo_63_tvalid,
    output [M_AXIS_FIFO_63_DMWIDTH/8-1:0] m_axis_fifo_63_tkeep,
    output [M_AXIS_FIFO_63_DMWIDTH/8-1:0] m_axis_fifo_63_tstrb,
    output [M_AXIS_FIFO_63_DMWIDTH-1:0] m_axis_fifo_63_tdata,
    input m_axis_fifo_63_tready,
    output ap_fifo_oarg_63_full_n,
    input [M_AXIS_FIFO_63_WIDTH-1:0] ap_fifo_oarg_63_din,
    input ap_fifo_oarg_63_write,
    //output FIFO to AXI-Stream interface 64
    input m_axis_fifo_64_aclk,
    input m_axis_fifo_64_aresetn,
    output m_axis_fifo_64_tlast,
    output m_axis_fifo_64_tvalid,
    output [M_AXIS_FIFO_64_DMWIDTH/8-1:0] m_axis_fifo_64_tkeep,
    output [M_AXIS_FIFO_64_DMWIDTH/8-1:0] m_axis_fifo_64_tstrb,
    output [M_AXIS_FIFO_64_DMWIDTH-1:0] m_axis_fifo_64_tdata,
    input m_axis_fifo_64_tready,
    output ap_fifo_oarg_64_full_n,
    input [M_AXIS_FIFO_64_WIDTH-1:0] ap_fifo_oarg_64_din,
    input ap_fifo_oarg_64_write,
    //output FIFO to AXI-Stream interface 65
    input m_axis_fifo_65_aclk,
    input m_axis_fifo_65_aresetn,
    output m_axis_fifo_65_tlast,
    output m_axis_fifo_65_tvalid,
    output [M_AXIS_FIFO_65_DMWIDTH/8-1:0] m_axis_fifo_65_tkeep,
    output [M_AXIS_FIFO_65_DMWIDTH/8-1:0] m_axis_fifo_65_tstrb,
    output [M_AXIS_FIFO_65_DMWIDTH-1:0] m_axis_fifo_65_tdata,
    input m_axis_fifo_65_tready,
    output ap_fifo_oarg_65_full_n,
    input [M_AXIS_FIFO_65_WIDTH-1:0] ap_fifo_oarg_65_din,
    input ap_fifo_oarg_65_write,
    //output FIFO to AXI-Stream interface 66
    input m_axis_fifo_66_aclk,
    input m_axis_fifo_66_aresetn,
    output m_axis_fifo_66_tlast,
    output m_axis_fifo_66_tvalid,
    output [M_AXIS_FIFO_66_DMWIDTH/8-1:0] m_axis_fifo_66_tkeep,
    output [M_AXIS_FIFO_66_DMWIDTH/8-1:0] m_axis_fifo_66_tstrb,
    output [M_AXIS_FIFO_66_DMWIDTH-1:0] m_axis_fifo_66_tdata,
    input m_axis_fifo_66_tready,
    output ap_fifo_oarg_66_full_n,
    input [M_AXIS_FIFO_66_WIDTH-1:0] ap_fifo_oarg_66_din,
    input ap_fifo_oarg_66_write,
    //output FIFO to AXI-Stream interface 67
    input m_axis_fifo_67_aclk,
    input m_axis_fifo_67_aresetn,
    output m_axis_fifo_67_tlast,
    output m_axis_fifo_67_tvalid,
    output [M_AXIS_FIFO_67_DMWIDTH/8-1:0] m_axis_fifo_67_tkeep,
    output [M_AXIS_FIFO_67_DMWIDTH/8-1:0] m_axis_fifo_67_tstrb,
    output [M_AXIS_FIFO_67_DMWIDTH-1:0] m_axis_fifo_67_tdata,
    input m_axis_fifo_67_tready,
    output ap_fifo_oarg_67_full_n,
    input [M_AXIS_FIFO_67_WIDTH-1:0] ap_fifo_oarg_67_din,
    input ap_fifo_oarg_67_write,
    //output FIFO to AXI-Stream interface 68
    input m_axis_fifo_68_aclk,
    input m_axis_fifo_68_aresetn,
    output m_axis_fifo_68_tlast,
    output m_axis_fifo_68_tvalid,
    output [M_AXIS_FIFO_68_DMWIDTH/8-1:0] m_axis_fifo_68_tkeep,
    output [M_AXIS_FIFO_68_DMWIDTH/8-1:0] m_axis_fifo_68_tstrb,
    output [M_AXIS_FIFO_68_DMWIDTH-1:0] m_axis_fifo_68_tdata,
    input m_axis_fifo_68_tready,
    output ap_fifo_oarg_68_full_n,
    input [M_AXIS_FIFO_68_WIDTH-1:0] ap_fifo_oarg_68_din,
    input ap_fifo_oarg_68_write,
    //output FIFO to AXI-Stream interface 69
    input m_axis_fifo_69_aclk,
    input m_axis_fifo_69_aresetn,
    output m_axis_fifo_69_tlast,
    output m_axis_fifo_69_tvalid,
    output [M_AXIS_FIFO_69_DMWIDTH/8-1:0] m_axis_fifo_69_tkeep,
    output [M_AXIS_FIFO_69_DMWIDTH/8-1:0] m_axis_fifo_69_tstrb,
    output [M_AXIS_FIFO_69_DMWIDTH-1:0] m_axis_fifo_69_tdata,
    input m_axis_fifo_69_tready,
    output ap_fifo_oarg_69_full_n,
    input [M_AXIS_FIFO_69_WIDTH-1:0] ap_fifo_oarg_69_din,
    input ap_fifo_oarg_69_write,
    //output FIFO to AXI-Stream interface 70
    input m_axis_fifo_70_aclk,
    input m_axis_fifo_70_aresetn,
    output m_axis_fifo_70_tlast,
    output m_axis_fifo_70_tvalid,
    output [M_AXIS_FIFO_70_DMWIDTH/8-1:0] m_axis_fifo_70_tkeep,
    output [M_AXIS_FIFO_70_DMWIDTH/8-1:0] m_axis_fifo_70_tstrb,
    output [M_AXIS_FIFO_70_DMWIDTH-1:0] m_axis_fifo_70_tdata,
    input m_axis_fifo_70_tready,
    output ap_fifo_oarg_70_full_n,
    input [M_AXIS_FIFO_70_WIDTH-1:0] ap_fifo_oarg_70_din,
    input ap_fifo_oarg_70_write,
    //output FIFO to AXI-Stream interface 71
    input m_axis_fifo_71_aclk,
    input m_axis_fifo_71_aresetn,
    output m_axis_fifo_71_tlast,
    output m_axis_fifo_71_tvalid,
    output [M_AXIS_FIFO_71_DMWIDTH/8-1:0] m_axis_fifo_71_tkeep,
    output [M_AXIS_FIFO_71_DMWIDTH/8-1:0] m_axis_fifo_71_tstrb,
    output [M_AXIS_FIFO_71_DMWIDTH-1:0] m_axis_fifo_71_tdata,
    input m_axis_fifo_71_tready,
    output ap_fifo_oarg_71_full_n,
    input [M_AXIS_FIFO_71_WIDTH-1:0] ap_fifo_oarg_71_din,
    input ap_fifo_oarg_71_write,
    //output FIFO to AXI-Stream interface 72
    input m_axis_fifo_72_aclk,
    input m_axis_fifo_72_aresetn,
    output m_axis_fifo_72_tlast,
    output m_axis_fifo_72_tvalid,
    output [M_AXIS_FIFO_72_DMWIDTH/8-1:0] m_axis_fifo_72_tkeep,
    output [M_AXIS_FIFO_72_DMWIDTH/8-1:0] m_axis_fifo_72_tstrb,
    output [M_AXIS_FIFO_72_DMWIDTH-1:0] m_axis_fifo_72_tdata,
    input m_axis_fifo_72_tready,
    output ap_fifo_oarg_72_full_n,
    input [M_AXIS_FIFO_72_WIDTH-1:0] ap_fifo_oarg_72_din,
    input ap_fifo_oarg_72_write,
    //output FIFO to AXI-Stream interface 73
    input m_axis_fifo_73_aclk,
    input m_axis_fifo_73_aresetn,
    output m_axis_fifo_73_tlast,
    output m_axis_fifo_73_tvalid,
    output [M_AXIS_FIFO_73_DMWIDTH/8-1:0] m_axis_fifo_73_tkeep,
    output [M_AXIS_FIFO_73_DMWIDTH/8-1:0] m_axis_fifo_73_tstrb,
    output [M_AXIS_FIFO_73_DMWIDTH-1:0] m_axis_fifo_73_tdata,
    input m_axis_fifo_73_tready,
    output ap_fifo_oarg_73_full_n,
    input [M_AXIS_FIFO_73_WIDTH-1:0] ap_fifo_oarg_73_din,
    input ap_fifo_oarg_73_write,
    //output FIFO to AXI-Stream interface 74
    input m_axis_fifo_74_aclk,
    input m_axis_fifo_74_aresetn,
    output m_axis_fifo_74_tlast,
    output m_axis_fifo_74_tvalid,
    output [M_AXIS_FIFO_74_DMWIDTH/8-1:0] m_axis_fifo_74_tkeep,
    output [M_AXIS_FIFO_74_DMWIDTH/8-1:0] m_axis_fifo_74_tstrb,
    output [M_AXIS_FIFO_74_DMWIDTH-1:0] m_axis_fifo_74_tdata,
    input m_axis_fifo_74_tready,
    output ap_fifo_oarg_74_full_n,
    input [M_AXIS_FIFO_74_WIDTH-1:0] ap_fifo_oarg_74_din,
    input ap_fifo_oarg_74_write,
    //output FIFO to AXI-Stream interface 75
    input m_axis_fifo_75_aclk,
    input m_axis_fifo_75_aresetn,
    output m_axis_fifo_75_tlast,
    output m_axis_fifo_75_tvalid,
    output [M_AXIS_FIFO_75_DMWIDTH/8-1:0] m_axis_fifo_75_tkeep,
    output [M_AXIS_FIFO_75_DMWIDTH/8-1:0] m_axis_fifo_75_tstrb,
    output [M_AXIS_FIFO_75_DMWIDTH-1:0] m_axis_fifo_75_tdata,
    input m_axis_fifo_75_tready,
    output ap_fifo_oarg_75_full_n,
    input [M_AXIS_FIFO_75_WIDTH-1:0] ap_fifo_oarg_75_din,
    input ap_fifo_oarg_75_write,
    //output FIFO to AXI-Stream interface 76
    input m_axis_fifo_76_aclk,
    input m_axis_fifo_76_aresetn,
    output m_axis_fifo_76_tlast,
    output m_axis_fifo_76_tvalid,
    output [M_AXIS_FIFO_76_DMWIDTH/8-1:0] m_axis_fifo_76_tkeep,
    output [M_AXIS_FIFO_76_DMWIDTH/8-1:0] m_axis_fifo_76_tstrb,
    output [M_AXIS_FIFO_76_DMWIDTH-1:0] m_axis_fifo_76_tdata,
    input m_axis_fifo_76_tready,
    output ap_fifo_oarg_76_full_n,
    input [M_AXIS_FIFO_76_WIDTH-1:0] ap_fifo_oarg_76_din,
    input ap_fifo_oarg_76_write,
    //output FIFO to AXI-Stream interface 77
    input m_axis_fifo_77_aclk,
    input m_axis_fifo_77_aresetn,
    output m_axis_fifo_77_tlast,
    output m_axis_fifo_77_tvalid,
    output [M_AXIS_FIFO_77_DMWIDTH/8-1:0] m_axis_fifo_77_tkeep,
    output [M_AXIS_FIFO_77_DMWIDTH/8-1:0] m_axis_fifo_77_tstrb,
    output [M_AXIS_FIFO_77_DMWIDTH-1:0] m_axis_fifo_77_tdata,
    input m_axis_fifo_77_tready,
    output ap_fifo_oarg_77_full_n,
    input [M_AXIS_FIFO_77_WIDTH-1:0] ap_fifo_oarg_77_din,
    input ap_fifo_oarg_77_write,
    //output FIFO to AXI-Stream interface 78
    input m_axis_fifo_78_aclk,
    input m_axis_fifo_78_aresetn,
    output m_axis_fifo_78_tlast,
    output m_axis_fifo_78_tvalid,
    output [M_AXIS_FIFO_78_DMWIDTH/8-1:0] m_axis_fifo_78_tkeep,
    output [M_AXIS_FIFO_78_DMWIDTH/8-1:0] m_axis_fifo_78_tstrb,
    output [M_AXIS_FIFO_78_DMWIDTH-1:0] m_axis_fifo_78_tdata,
    input m_axis_fifo_78_tready,
    output ap_fifo_oarg_78_full_n,
    input [M_AXIS_FIFO_78_WIDTH-1:0] ap_fifo_oarg_78_din,
    input ap_fifo_oarg_78_write,
    //output FIFO to AXI-Stream interface 79
    input m_axis_fifo_79_aclk,
    input m_axis_fifo_79_aresetn,
    output m_axis_fifo_79_tlast,
    output m_axis_fifo_79_tvalid,
    output [M_AXIS_FIFO_79_DMWIDTH/8-1:0] m_axis_fifo_79_tkeep,
    output [M_AXIS_FIFO_79_DMWIDTH/8-1:0] m_axis_fifo_79_tstrb,
    output [M_AXIS_FIFO_79_DMWIDTH-1:0] m_axis_fifo_79_tdata,
    input m_axis_fifo_79_tready,
    output ap_fifo_oarg_79_full_n,
    input [M_AXIS_FIFO_79_WIDTH-1:0] ap_fifo_oarg_79_din,
    input ap_fifo_oarg_79_write,
    //output FIFO to AXI-Stream interface 80
    input m_axis_fifo_80_aclk,
    input m_axis_fifo_80_aresetn,
    output m_axis_fifo_80_tlast,
    output m_axis_fifo_80_tvalid,
    output [M_AXIS_FIFO_80_DMWIDTH/8-1:0] m_axis_fifo_80_tkeep,
    output [M_AXIS_FIFO_80_DMWIDTH/8-1:0] m_axis_fifo_80_tstrb,
    output [M_AXIS_FIFO_80_DMWIDTH-1:0] m_axis_fifo_80_tdata,
    input m_axis_fifo_80_tready,
    output ap_fifo_oarg_80_full_n,
    input [M_AXIS_FIFO_80_WIDTH-1:0] ap_fifo_oarg_80_din,
    input ap_fifo_oarg_80_write,
    //output FIFO to AXI-Stream interface 81
    input m_axis_fifo_81_aclk,
    input m_axis_fifo_81_aresetn,
    output m_axis_fifo_81_tlast,
    output m_axis_fifo_81_tvalid,
    output [M_AXIS_FIFO_81_DMWIDTH/8-1:0] m_axis_fifo_81_tkeep,
    output [M_AXIS_FIFO_81_DMWIDTH/8-1:0] m_axis_fifo_81_tstrb,
    output [M_AXIS_FIFO_81_DMWIDTH-1:0] m_axis_fifo_81_tdata,
    input m_axis_fifo_81_tready,
    output ap_fifo_oarg_81_full_n,
    input [M_AXIS_FIFO_81_WIDTH-1:0] ap_fifo_oarg_81_din,
    input ap_fifo_oarg_81_write,
    //output FIFO to AXI-Stream interface 82
    input m_axis_fifo_82_aclk,
    input m_axis_fifo_82_aresetn,
    output m_axis_fifo_82_tlast,
    output m_axis_fifo_82_tvalid,
    output [M_AXIS_FIFO_82_DMWIDTH/8-1:0] m_axis_fifo_82_tkeep,
    output [M_AXIS_FIFO_82_DMWIDTH/8-1:0] m_axis_fifo_82_tstrb,
    output [M_AXIS_FIFO_82_DMWIDTH-1:0] m_axis_fifo_82_tdata,
    input m_axis_fifo_82_tready,
    output ap_fifo_oarg_82_full_n,
    input [M_AXIS_FIFO_82_WIDTH-1:0] ap_fifo_oarg_82_din,
    input ap_fifo_oarg_82_write,
    //output FIFO to AXI-Stream interface 83
    input m_axis_fifo_83_aclk,
    input m_axis_fifo_83_aresetn,
    output m_axis_fifo_83_tlast,
    output m_axis_fifo_83_tvalid,
    output [M_AXIS_FIFO_83_DMWIDTH/8-1:0] m_axis_fifo_83_tkeep,
    output [M_AXIS_FIFO_83_DMWIDTH/8-1:0] m_axis_fifo_83_tstrb,
    output [M_AXIS_FIFO_83_DMWIDTH-1:0] m_axis_fifo_83_tdata,
    input m_axis_fifo_83_tready,
    output ap_fifo_oarg_83_full_n,
    input [M_AXIS_FIFO_83_WIDTH-1:0] ap_fifo_oarg_83_din,
    input ap_fifo_oarg_83_write,
    //output FIFO to AXI-Stream interface 84
    input m_axis_fifo_84_aclk,
    input m_axis_fifo_84_aresetn,
    output m_axis_fifo_84_tlast,
    output m_axis_fifo_84_tvalid,
    output [M_AXIS_FIFO_84_DMWIDTH/8-1:0] m_axis_fifo_84_tkeep,
    output [M_AXIS_FIFO_84_DMWIDTH/8-1:0] m_axis_fifo_84_tstrb,
    output [M_AXIS_FIFO_84_DMWIDTH-1:0] m_axis_fifo_84_tdata,
    input m_axis_fifo_84_tready,
    output ap_fifo_oarg_84_full_n,
    input [M_AXIS_FIFO_84_WIDTH-1:0] ap_fifo_oarg_84_din,
    input ap_fifo_oarg_84_write,
    //output FIFO to AXI-Stream interface 85
    input m_axis_fifo_85_aclk,
    input m_axis_fifo_85_aresetn,
    output m_axis_fifo_85_tlast,
    output m_axis_fifo_85_tvalid,
    output [M_AXIS_FIFO_85_DMWIDTH/8-1:0] m_axis_fifo_85_tkeep,
    output [M_AXIS_FIFO_85_DMWIDTH/8-1:0] m_axis_fifo_85_tstrb,
    output [M_AXIS_FIFO_85_DMWIDTH-1:0] m_axis_fifo_85_tdata,
    input m_axis_fifo_85_tready,
    output ap_fifo_oarg_85_full_n,
    input [M_AXIS_FIFO_85_WIDTH-1:0] ap_fifo_oarg_85_din,
    input ap_fifo_oarg_85_write,
    //output FIFO to AXI-Stream interface 86
    input m_axis_fifo_86_aclk,
    input m_axis_fifo_86_aresetn,
    output m_axis_fifo_86_tlast,
    output m_axis_fifo_86_tvalid,
    output [M_AXIS_FIFO_86_DMWIDTH/8-1:0] m_axis_fifo_86_tkeep,
    output [M_AXIS_FIFO_86_DMWIDTH/8-1:0] m_axis_fifo_86_tstrb,
    output [M_AXIS_FIFO_86_DMWIDTH-1:0] m_axis_fifo_86_tdata,
    input m_axis_fifo_86_tready,
    output ap_fifo_oarg_86_full_n,
    input [M_AXIS_FIFO_86_WIDTH-1:0] ap_fifo_oarg_86_din,
    input ap_fifo_oarg_86_write,
    //output FIFO to AXI-Stream interface 87
    input m_axis_fifo_87_aclk,
    input m_axis_fifo_87_aresetn,
    output m_axis_fifo_87_tlast,
    output m_axis_fifo_87_tvalid,
    output [M_AXIS_FIFO_87_DMWIDTH/8-1:0] m_axis_fifo_87_tkeep,
    output [M_AXIS_FIFO_87_DMWIDTH/8-1:0] m_axis_fifo_87_tstrb,
    output [M_AXIS_FIFO_87_DMWIDTH-1:0] m_axis_fifo_87_tdata,
    input m_axis_fifo_87_tready,
    output ap_fifo_oarg_87_full_n,
    input [M_AXIS_FIFO_87_WIDTH-1:0] ap_fifo_oarg_87_din,
    input ap_fifo_oarg_87_write,
    //output FIFO to AXI-Stream interface 88
    input m_axis_fifo_88_aclk,
    input m_axis_fifo_88_aresetn,
    output m_axis_fifo_88_tlast,
    output m_axis_fifo_88_tvalid,
    output [M_AXIS_FIFO_88_DMWIDTH/8-1:0] m_axis_fifo_88_tkeep,
    output [M_AXIS_FIFO_88_DMWIDTH/8-1:0] m_axis_fifo_88_tstrb,
    output [M_AXIS_FIFO_88_DMWIDTH-1:0] m_axis_fifo_88_tdata,
    input m_axis_fifo_88_tready,
    output ap_fifo_oarg_88_full_n,
    input [M_AXIS_FIFO_88_WIDTH-1:0] ap_fifo_oarg_88_din,
    input ap_fifo_oarg_88_write,
    //output FIFO to AXI-Stream interface 89
    input m_axis_fifo_89_aclk,
    input m_axis_fifo_89_aresetn,
    output m_axis_fifo_89_tlast,
    output m_axis_fifo_89_tvalid,
    output [M_AXIS_FIFO_89_DMWIDTH/8-1:0] m_axis_fifo_89_tkeep,
    output [M_AXIS_FIFO_89_DMWIDTH/8-1:0] m_axis_fifo_89_tstrb,
    output [M_AXIS_FIFO_89_DMWIDTH-1:0] m_axis_fifo_89_tdata,
    input m_axis_fifo_89_tready,
    output ap_fifo_oarg_89_full_n,
    input [M_AXIS_FIFO_89_WIDTH-1:0] ap_fifo_oarg_89_din,
    input ap_fifo_oarg_89_write,
    //output FIFO to AXI-Stream interface 90
    input m_axis_fifo_90_aclk,
    input m_axis_fifo_90_aresetn,
    output m_axis_fifo_90_tlast,
    output m_axis_fifo_90_tvalid,
    output [M_AXIS_FIFO_90_DMWIDTH/8-1:0] m_axis_fifo_90_tkeep,
    output [M_AXIS_FIFO_90_DMWIDTH/8-1:0] m_axis_fifo_90_tstrb,
    output [M_AXIS_FIFO_90_DMWIDTH-1:0] m_axis_fifo_90_tdata,
    input m_axis_fifo_90_tready,
    output ap_fifo_oarg_90_full_n,
    input [M_AXIS_FIFO_90_WIDTH-1:0] ap_fifo_oarg_90_din,
    input ap_fifo_oarg_90_write,
    //output FIFO to AXI-Stream interface 91
    input m_axis_fifo_91_aclk,
    input m_axis_fifo_91_aresetn,
    output m_axis_fifo_91_tlast,
    output m_axis_fifo_91_tvalid,
    output [M_AXIS_FIFO_91_DMWIDTH/8-1:0] m_axis_fifo_91_tkeep,
    output [M_AXIS_FIFO_91_DMWIDTH/8-1:0] m_axis_fifo_91_tstrb,
    output [M_AXIS_FIFO_91_DMWIDTH-1:0] m_axis_fifo_91_tdata,
    input m_axis_fifo_91_tready,
    output ap_fifo_oarg_91_full_n,
    input [M_AXIS_FIFO_91_WIDTH-1:0] ap_fifo_oarg_91_din,
    input ap_fifo_oarg_91_write,
    //output FIFO to AXI-Stream interface 92
    input m_axis_fifo_92_aclk,
    input m_axis_fifo_92_aresetn,
    output m_axis_fifo_92_tlast,
    output m_axis_fifo_92_tvalid,
    output [M_AXIS_FIFO_92_DMWIDTH/8-1:0] m_axis_fifo_92_tkeep,
    output [M_AXIS_FIFO_92_DMWIDTH/8-1:0] m_axis_fifo_92_tstrb,
    output [M_AXIS_FIFO_92_DMWIDTH-1:0] m_axis_fifo_92_tdata,
    input m_axis_fifo_92_tready,
    output ap_fifo_oarg_92_full_n,
    input [M_AXIS_FIFO_92_WIDTH-1:0] ap_fifo_oarg_92_din,
    input ap_fifo_oarg_92_write,
    //output FIFO to AXI-Stream interface 93
    input m_axis_fifo_93_aclk,
    input m_axis_fifo_93_aresetn,
    output m_axis_fifo_93_tlast,
    output m_axis_fifo_93_tvalid,
    output [M_AXIS_FIFO_93_DMWIDTH/8-1:0] m_axis_fifo_93_tkeep,
    output [M_AXIS_FIFO_93_DMWIDTH/8-1:0] m_axis_fifo_93_tstrb,
    output [M_AXIS_FIFO_93_DMWIDTH-1:0] m_axis_fifo_93_tdata,
    input m_axis_fifo_93_tready,
    output ap_fifo_oarg_93_full_n,
    input [M_AXIS_FIFO_93_WIDTH-1:0] ap_fifo_oarg_93_din,
    input ap_fifo_oarg_93_write,
    //output FIFO to AXI-Stream interface 94
    input m_axis_fifo_94_aclk,
    input m_axis_fifo_94_aresetn,
    output m_axis_fifo_94_tlast,
    output m_axis_fifo_94_tvalid,
    output [M_AXIS_FIFO_94_DMWIDTH/8-1:0] m_axis_fifo_94_tkeep,
    output [M_AXIS_FIFO_94_DMWIDTH/8-1:0] m_axis_fifo_94_tstrb,
    output [M_AXIS_FIFO_94_DMWIDTH-1:0] m_axis_fifo_94_tdata,
    input m_axis_fifo_94_tready,
    output ap_fifo_oarg_94_full_n,
    input [M_AXIS_FIFO_94_WIDTH-1:0] ap_fifo_oarg_94_din,
    input ap_fifo_oarg_94_write,
    //output FIFO to AXI-Stream interface 95
    input m_axis_fifo_95_aclk,
    input m_axis_fifo_95_aresetn,
    output m_axis_fifo_95_tlast,
    output m_axis_fifo_95_tvalid,
    output [M_AXIS_FIFO_95_DMWIDTH/8-1:0] m_axis_fifo_95_tkeep,
    output [M_AXIS_FIFO_95_DMWIDTH/8-1:0] m_axis_fifo_95_tstrb,
    output [M_AXIS_FIFO_95_DMWIDTH-1:0] m_axis_fifo_95_tdata,
    input m_axis_fifo_95_tready,
    output ap_fifo_oarg_95_full_n,
    input [M_AXIS_FIFO_95_WIDTH-1:0] ap_fifo_oarg_95_din,
    input ap_fifo_oarg_95_write,
    //output FIFO to AXI-Stream interface 96
    input m_axis_fifo_96_aclk,
    input m_axis_fifo_96_aresetn,
    output m_axis_fifo_96_tlast,
    output m_axis_fifo_96_tvalid,
    output [M_AXIS_FIFO_96_DMWIDTH/8-1:0] m_axis_fifo_96_tkeep,
    output [M_AXIS_FIFO_96_DMWIDTH/8-1:0] m_axis_fifo_96_tstrb,
    output [M_AXIS_FIFO_96_DMWIDTH-1:0] m_axis_fifo_96_tdata,
    input m_axis_fifo_96_tready,
    output ap_fifo_oarg_96_full_n,
    input [M_AXIS_FIFO_96_WIDTH-1:0] ap_fifo_oarg_96_din,
    input ap_fifo_oarg_96_write,
    //output FIFO to AXI-Stream interface 97
    input m_axis_fifo_97_aclk,
    input m_axis_fifo_97_aresetn,
    output m_axis_fifo_97_tlast,
    output m_axis_fifo_97_tvalid,
    output [M_AXIS_FIFO_97_DMWIDTH/8-1:0] m_axis_fifo_97_tkeep,
    output [M_AXIS_FIFO_97_DMWIDTH/8-1:0] m_axis_fifo_97_tstrb,
    output [M_AXIS_FIFO_97_DMWIDTH-1:0] m_axis_fifo_97_tdata,
    input m_axis_fifo_97_tready,
    output ap_fifo_oarg_97_full_n,
    input [M_AXIS_FIFO_97_WIDTH-1:0] ap_fifo_oarg_97_din,
    input ap_fifo_oarg_97_write,
    //output FIFO to AXI-Stream interface 98
    input m_axis_fifo_98_aclk,
    input m_axis_fifo_98_aresetn,
    output m_axis_fifo_98_tlast,
    output m_axis_fifo_98_tvalid,
    output [M_AXIS_FIFO_98_DMWIDTH/8-1:0] m_axis_fifo_98_tkeep,
    output [M_AXIS_FIFO_98_DMWIDTH/8-1:0] m_axis_fifo_98_tstrb,
    output [M_AXIS_FIFO_98_DMWIDTH-1:0] m_axis_fifo_98_tdata,
    input m_axis_fifo_98_tready,
    output ap_fifo_oarg_98_full_n,
    input [M_AXIS_FIFO_98_WIDTH-1:0] ap_fifo_oarg_98_din,
    input ap_fifo_oarg_98_write,
    //output FIFO to AXI-Stream interface 99
    input m_axis_fifo_99_aclk,
    input m_axis_fifo_99_aresetn,
    output m_axis_fifo_99_tlast,
    output m_axis_fifo_99_tvalid,
    output [M_AXIS_FIFO_99_DMWIDTH/8-1:0] m_axis_fifo_99_tkeep,
    output [M_AXIS_FIFO_99_DMWIDTH/8-1:0] m_axis_fifo_99_tstrb,
    output [M_AXIS_FIFO_99_DMWIDTH-1:0] m_axis_fifo_99_tdata,
    input m_axis_fifo_99_tready,
    output ap_fifo_oarg_99_full_n,
    input [M_AXIS_FIFO_99_WIDTH-1:0] ap_fifo_oarg_99_din,
    input ap_fifo_oarg_99_write,
    //output FIFO to AXI-Stream interface 100
    input m_axis_fifo_100_aclk,
    input m_axis_fifo_100_aresetn,
    output m_axis_fifo_100_tlast,
    output m_axis_fifo_100_tvalid,
    output [M_AXIS_FIFO_100_DMWIDTH/8-1:0] m_axis_fifo_100_tkeep,
    output [M_AXIS_FIFO_100_DMWIDTH/8-1:0] m_axis_fifo_100_tstrb,
    output [M_AXIS_FIFO_100_DMWIDTH-1:0] m_axis_fifo_100_tdata,
    input m_axis_fifo_100_tready,
    output ap_fifo_oarg_100_full_n,
    input [M_AXIS_FIFO_100_WIDTH-1:0] ap_fifo_oarg_100_din,
    input ap_fifo_oarg_100_write,
    //output FIFO to AXI-Stream interface 101
    input m_axis_fifo_101_aclk,
    input m_axis_fifo_101_aresetn,
    output m_axis_fifo_101_tlast,
    output m_axis_fifo_101_tvalid,
    output [M_AXIS_FIFO_101_DMWIDTH/8-1:0] m_axis_fifo_101_tkeep,
    output [M_AXIS_FIFO_101_DMWIDTH/8-1:0] m_axis_fifo_101_tstrb,
    output [M_AXIS_FIFO_101_DMWIDTH-1:0] m_axis_fifo_101_tdata,
    input m_axis_fifo_101_tready,
    output ap_fifo_oarg_101_full_n,
    input [M_AXIS_FIFO_101_WIDTH-1:0] ap_fifo_oarg_101_din,
    input ap_fifo_oarg_101_write,
    //output FIFO to AXI-Stream interface 102
    input m_axis_fifo_102_aclk,
    input m_axis_fifo_102_aresetn,
    output m_axis_fifo_102_tlast,
    output m_axis_fifo_102_tvalid,
    output [M_AXIS_FIFO_102_DMWIDTH/8-1:0] m_axis_fifo_102_tkeep,
    output [M_AXIS_FIFO_102_DMWIDTH/8-1:0] m_axis_fifo_102_tstrb,
    output [M_AXIS_FIFO_102_DMWIDTH-1:0] m_axis_fifo_102_tdata,
    input m_axis_fifo_102_tready,
    output ap_fifo_oarg_102_full_n,
    input [M_AXIS_FIFO_102_WIDTH-1:0] ap_fifo_oarg_102_din,
    input ap_fifo_oarg_102_write,
    //output FIFO to AXI-Stream interface 103
    input m_axis_fifo_103_aclk,
    input m_axis_fifo_103_aresetn,
    output m_axis_fifo_103_tlast,
    output m_axis_fifo_103_tvalid,
    output [M_AXIS_FIFO_103_DMWIDTH/8-1:0] m_axis_fifo_103_tkeep,
    output [M_AXIS_FIFO_103_DMWIDTH/8-1:0] m_axis_fifo_103_tstrb,
    output [M_AXIS_FIFO_103_DMWIDTH-1:0] m_axis_fifo_103_tdata,
    input m_axis_fifo_103_tready,
    output ap_fifo_oarg_103_full_n,
    input [M_AXIS_FIFO_103_WIDTH-1:0] ap_fifo_oarg_103_din,
    input ap_fifo_oarg_103_write,
    //output FIFO to AXI-Stream interface 104
    input m_axis_fifo_104_aclk,
    input m_axis_fifo_104_aresetn,
    output m_axis_fifo_104_tlast,
    output m_axis_fifo_104_tvalid,
    output [M_AXIS_FIFO_104_DMWIDTH/8-1:0] m_axis_fifo_104_tkeep,
    output [M_AXIS_FIFO_104_DMWIDTH/8-1:0] m_axis_fifo_104_tstrb,
    output [M_AXIS_FIFO_104_DMWIDTH-1:0] m_axis_fifo_104_tdata,
    input m_axis_fifo_104_tready,
    output ap_fifo_oarg_104_full_n,
    input [M_AXIS_FIFO_104_WIDTH-1:0] ap_fifo_oarg_104_din,
    input ap_fifo_oarg_104_write,
    //output FIFO to AXI-Stream interface 105
    input m_axis_fifo_105_aclk,
    input m_axis_fifo_105_aresetn,
    output m_axis_fifo_105_tlast,
    output m_axis_fifo_105_tvalid,
    output [M_AXIS_FIFO_105_DMWIDTH/8-1:0] m_axis_fifo_105_tkeep,
    output [M_AXIS_FIFO_105_DMWIDTH/8-1:0] m_axis_fifo_105_tstrb,
    output [M_AXIS_FIFO_105_DMWIDTH-1:0] m_axis_fifo_105_tdata,
    input m_axis_fifo_105_tready,
    output ap_fifo_oarg_105_full_n,
    input [M_AXIS_FIFO_105_WIDTH-1:0] ap_fifo_oarg_105_din,
    input ap_fifo_oarg_105_write,
    //output FIFO to AXI-Stream interface 106
    input m_axis_fifo_106_aclk,
    input m_axis_fifo_106_aresetn,
    output m_axis_fifo_106_tlast,
    output m_axis_fifo_106_tvalid,
    output [M_AXIS_FIFO_106_DMWIDTH/8-1:0] m_axis_fifo_106_tkeep,
    output [M_AXIS_FIFO_106_DMWIDTH/8-1:0] m_axis_fifo_106_tstrb,
    output [M_AXIS_FIFO_106_DMWIDTH-1:0] m_axis_fifo_106_tdata,
    input m_axis_fifo_106_tready,
    output ap_fifo_oarg_106_full_n,
    input [M_AXIS_FIFO_106_WIDTH-1:0] ap_fifo_oarg_106_din,
    input ap_fifo_oarg_106_write,
    //output FIFO to AXI-Stream interface 107
    input m_axis_fifo_107_aclk,
    input m_axis_fifo_107_aresetn,
    output m_axis_fifo_107_tlast,
    output m_axis_fifo_107_tvalid,
    output [M_AXIS_FIFO_107_DMWIDTH/8-1:0] m_axis_fifo_107_tkeep,
    output [M_AXIS_FIFO_107_DMWIDTH/8-1:0] m_axis_fifo_107_tstrb,
    output [M_AXIS_FIFO_107_DMWIDTH-1:0] m_axis_fifo_107_tdata,
    input m_axis_fifo_107_tready,
    output ap_fifo_oarg_107_full_n,
    input [M_AXIS_FIFO_107_WIDTH-1:0] ap_fifo_oarg_107_din,
    input ap_fifo_oarg_107_write,
    //output FIFO to AXI-Stream interface 108
    input m_axis_fifo_108_aclk,
    input m_axis_fifo_108_aresetn,
    output m_axis_fifo_108_tlast,
    output m_axis_fifo_108_tvalid,
    output [M_AXIS_FIFO_108_DMWIDTH/8-1:0] m_axis_fifo_108_tkeep,
    output [M_AXIS_FIFO_108_DMWIDTH/8-1:0] m_axis_fifo_108_tstrb,
    output [M_AXIS_FIFO_108_DMWIDTH-1:0] m_axis_fifo_108_tdata,
    input m_axis_fifo_108_tready,
    output ap_fifo_oarg_108_full_n,
    input [M_AXIS_FIFO_108_WIDTH-1:0] ap_fifo_oarg_108_din,
    input ap_fifo_oarg_108_write,
    //output FIFO to AXI-Stream interface 109
    input m_axis_fifo_109_aclk,
    input m_axis_fifo_109_aresetn,
    output m_axis_fifo_109_tlast,
    output m_axis_fifo_109_tvalid,
    output [M_AXIS_FIFO_109_DMWIDTH/8-1:0] m_axis_fifo_109_tkeep,
    output [M_AXIS_FIFO_109_DMWIDTH/8-1:0] m_axis_fifo_109_tstrb,
    output [M_AXIS_FIFO_109_DMWIDTH-1:0] m_axis_fifo_109_tdata,
    input m_axis_fifo_109_tready,
    output ap_fifo_oarg_109_full_n,
    input [M_AXIS_FIFO_109_WIDTH-1:0] ap_fifo_oarg_109_din,
    input ap_fifo_oarg_109_write,
    //output FIFO to AXI-Stream interface 110
    input m_axis_fifo_110_aclk,
    input m_axis_fifo_110_aresetn,
    output m_axis_fifo_110_tlast,
    output m_axis_fifo_110_tvalid,
    output [M_AXIS_FIFO_110_DMWIDTH/8-1:0] m_axis_fifo_110_tkeep,
    output [M_AXIS_FIFO_110_DMWIDTH/8-1:0] m_axis_fifo_110_tstrb,
    output [M_AXIS_FIFO_110_DMWIDTH-1:0] m_axis_fifo_110_tdata,
    input m_axis_fifo_110_tready,
    output ap_fifo_oarg_110_full_n,
    input [M_AXIS_FIFO_110_WIDTH-1:0] ap_fifo_oarg_110_din,
    input ap_fifo_oarg_110_write,
    //output FIFO to AXI-Stream interface 111
    input m_axis_fifo_111_aclk,
    input m_axis_fifo_111_aresetn,
    output m_axis_fifo_111_tlast,
    output m_axis_fifo_111_tvalid,
    output [M_AXIS_FIFO_111_DMWIDTH/8-1:0] m_axis_fifo_111_tkeep,
    output [M_AXIS_FIFO_111_DMWIDTH/8-1:0] m_axis_fifo_111_tstrb,
    output [M_AXIS_FIFO_111_DMWIDTH-1:0] m_axis_fifo_111_tdata,
    input m_axis_fifo_111_tready,
    output ap_fifo_oarg_111_full_n,
    input [M_AXIS_FIFO_111_WIDTH-1:0] ap_fifo_oarg_111_din,
    input ap_fifo_oarg_111_write,
    //output FIFO to AXI-Stream interface 112
    input m_axis_fifo_112_aclk,
    input m_axis_fifo_112_aresetn,
    output m_axis_fifo_112_tlast,
    output m_axis_fifo_112_tvalid,
    output [M_AXIS_FIFO_112_DMWIDTH/8-1:0] m_axis_fifo_112_tkeep,
    output [M_AXIS_FIFO_112_DMWIDTH/8-1:0] m_axis_fifo_112_tstrb,
    output [M_AXIS_FIFO_112_DMWIDTH-1:0] m_axis_fifo_112_tdata,
    input m_axis_fifo_112_tready,
    output ap_fifo_oarg_112_full_n,
    input [M_AXIS_FIFO_112_WIDTH-1:0] ap_fifo_oarg_112_din,
    input ap_fifo_oarg_112_write,
    //output FIFO to AXI-Stream interface 113
    input m_axis_fifo_113_aclk,
    input m_axis_fifo_113_aresetn,
    output m_axis_fifo_113_tlast,
    output m_axis_fifo_113_tvalid,
    output [M_AXIS_FIFO_113_DMWIDTH/8-1:0] m_axis_fifo_113_tkeep,
    output [M_AXIS_FIFO_113_DMWIDTH/8-1:0] m_axis_fifo_113_tstrb,
    output [M_AXIS_FIFO_113_DMWIDTH-1:0] m_axis_fifo_113_tdata,
    input m_axis_fifo_113_tready,
    output ap_fifo_oarg_113_full_n,
    input [M_AXIS_FIFO_113_WIDTH-1:0] ap_fifo_oarg_113_din,
    input ap_fifo_oarg_113_write,
    //output FIFO to AXI-Stream interface 114
    input m_axis_fifo_114_aclk,
    input m_axis_fifo_114_aresetn,
    output m_axis_fifo_114_tlast,
    output m_axis_fifo_114_tvalid,
    output [M_AXIS_FIFO_114_DMWIDTH/8-1:0] m_axis_fifo_114_tkeep,
    output [M_AXIS_FIFO_114_DMWIDTH/8-1:0] m_axis_fifo_114_tstrb,
    output [M_AXIS_FIFO_114_DMWIDTH-1:0] m_axis_fifo_114_tdata,
    input m_axis_fifo_114_tready,
    output ap_fifo_oarg_114_full_n,
    input [M_AXIS_FIFO_114_WIDTH-1:0] ap_fifo_oarg_114_din,
    input ap_fifo_oarg_114_write,
    //output FIFO to AXI-Stream interface 115
    input m_axis_fifo_115_aclk,
    input m_axis_fifo_115_aresetn,
    output m_axis_fifo_115_tlast,
    output m_axis_fifo_115_tvalid,
    output [M_AXIS_FIFO_115_DMWIDTH/8-1:0] m_axis_fifo_115_tkeep,
    output [M_AXIS_FIFO_115_DMWIDTH/8-1:0] m_axis_fifo_115_tstrb,
    output [M_AXIS_FIFO_115_DMWIDTH-1:0] m_axis_fifo_115_tdata,
    input m_axis_fifo_115_tready,
    output ap_fifo_oarg_115_full_n,
    input [M_AXIS_FIFO_115_WIDTH-1:0] ap_fifo_oarg_115_din,
    input ap_fifo_oarg_115_write,
    //output FIFO to AXI-Stream interface 116
    input m_axis_fifo_116_aclk,
    input m_axis_fifo_116_aresetn,
    output m_axis_fifo_116_tlast,
    output m_axis_fifo_116_tvalid,
    output [M_AXIS_FIFO_116_DMWIDTH/8-1:0] m_axis_fifo_116_tkeep,
    output [M_AXIS_FIFO_116_DMWIDTH/8-1:0] m_axis_fifo_116_tstrb,
    output [M_AXIS_FIFO_116_DMWIDTH-1:0] m_axis_fifo_116_tdata,
    input m_axis_fifo_116_tready,
    output ap_fifo_oarg_116_full_n,
    input [M_AXIS_FIFO_116_WIDTH-1:0] ap_fifo_oarg_116_din,
    input ap_fifo_oarg_116_write,
    //output FIFO to AXI-Stream interface 117
    input m_axis_fifo_117_aclk,
    input m_axis_fifo_117_aresetn,
    output m_axis_fifo_117_tlast,
    output m_axis_fifo_117_tvalid,
    output [M_AXIS_FIFO_117_DMWIDTH/8-1:0] m_axis_fifo_117_tkeep,
    output [M_AXIS_FIFO_117_DMWIDTH/8-1:0] m_axis_fifo_117_tstrb,
    output [M_AXIS_FIFO_117_DMWIDTH-1:0] m_axis_fifo_117_tdata,
    input m_axis_fifo_117_tready,
    output ap_fifo_oarg_117_full_n,
    input [M_AXIS_FIFO_117_WIDTH-1:0] ap_fifo_oarg_117_din,
    input ap_fifo_oarg_117_write,
    //output FIFO to AXI-Stream interface 118
    input m_axis_fifo_118_aclk,
    input m_axis_fifo_118_aresetn,
    output m_axis_fifo_118_tlast,
    output m_axis_fifo_118_tvalid,
    output [M_AXIS_FIFO_118_DMWIDTH/8-1:0] m_axis_fifo_118_tkeep,
    output [M_AXIS_FIFO_118_DMWIDTH/8-1:0] m_axis_fifo_118_tstrb,
    output [M_AXIS_FIFO_118_DMWIDTH-1:0] m_axis_fifo_118_tdata,
    input m_axis_fifo_118_tready,
    output ap_fifo_oarg_118_full_n,
    input [M_AXIS_FIFO_118_WIDTH-1:0] ap_fifo_oarg_118_din,
    input ap_fifo_oarg_118_write,
    //output FIFO to AXI-Stream interface 119
    input m_axis_fifo_119_aclk,
    input m_axis_fifo_119_aresetn,
    output m_axis_fifo_119_tlast,
    output m_axis_fifo_119_tvalid,
    output [M_AXIS_FIFO_119_DMWIDTH/8-1:0] m_axis_fifo_119_tkeep,
    output [M_AXIS_FIFO_119_DMWIDTH/8-1:0] m_axis_fifo_119_tstrb,
    output [M_AXIS_FIFO_119_DMWIDTH-1:0] m_axis_fifo_119_tdata,
    input m_axis_fifo_119_tready,
    output ap_fifo_oarg_119_full_n,
    input [M_AXIS_FIFO_119_WIDTH-1:0] ap_fifo_oarg_119_din,
    input ap_fifo_oarg_119_write,
    //output FIFO to AXI-Stream interface 120
    input m_axis_fifo_120_aclk,
    input m_axis_fifo_120_aresetn,
    output m_axis_fifo_120_tlast,
    output m_axis_fifo_120_tvalid,
    output [M_AXIS_FIFO_120_DMWIDTH/8-1:0] m_axis_fifo_120_tkeep,
    output [M_AXIS_FIFO_120_DMWIDTH/8-1:0] m_axis_fifo_120_tstrb,
    output [M_AXIS_FIFO_120_DMWIDTH-1:0] m_axis_fifo_120_tdata,
    input m_axis_fifo_120_tready,
    output ap_fifo_oarg_120_full_n,
    input [M_AXIS_FIFO_120_WIDTH-1:0] ap_fifo_oarg_120_din,
    input ap_fifo_oarg_120_write,
    //output FIFO to AXI-Stream interface 121
    input m_axis_fifo_121_aclk,
    input m_axis_fifo_121_aresetn,
    output m_axis_fifo_121_tlast,
    output m_axis_fifo_121_tvalid,
    output [M_AXIS_FIFO_121_DMWIDTH/8-1:0] m_axis_fifo_121_tkeep,
    output [M_AXIS_FIFO_121_DMWIDTH/8-1:0] m_axis_fifo_121_tstrb,
    output [M_AXIS_FIFO_121_DMWIDTH-1:0] m_axis_fifo_121_tdata,
    input m_axis_fifo_121_tready,
    output ap_fifo_oarg_121_full_n,
    input [M_AXIS_FIFO_121_WIDTH-1:0] ap_fifo_oarg_121_din,
    input ap_fifo_oarg_121_write,
    //output FIFO to AXI-Stream interface 122
    input m_axis_fifo_122_aclk,
    input m_axis_fifo_122_aresetn,
    output m_axis_fifo_122_tlast,
    output m_axis_fifo_122_tvalid,
    output [M_AXIS_FIFO_122_DMWIDTH/8-1:0] m_axis_fifo_122_tkeep,
    output [M_AXIS_FIFO_122_DMWIDTH/8-1:0] m_axis_fifo_122_tstrb,
    output [M_AXIS_FIFO_122_DMWIDTH-1:0] m_axis_fifo_122_tdata,
    input m_axis_fifo_122_tready,
    output ap_fifo_oarg_122_full_n,
    input [M_AXIS_FIFO_122_WIDTH-1:0] ap_fifo_oarg_122_din,
    input ap_fifo_oarg_122_write,
    //output FIFO to AXI-Stream interface 123
    input m_axis_fifo_123_aclk,
    input m_axis_fifo_123_aresetn,
    output m_axis_fifo_123_tlast,
    output m_axis_fifo_123_tvalid,
    output [M_AXIS_FIFO_123_DMWIDTH/8-1:0] m_axis_fifo_123_tkeep,
    output [M_AXIS_FIFO_123_DMWIDTH/8-1:0] m_axis_fifo_123_tstrb,
    output [M_AXIS_FIFO_123_DMWIDTH-1:0] m_axis_fifo_123_tdata,
    input m_axis_fifo_123_tready,
    output ap_fifo_oarg_123_full_n,
    input [M_AXIS_FIFO_123_WIDTH-1:0] ap_fifo_oarg_123_din,
    input ap_fifo_oarg_123_write,
    //output FIFO to AXI-Stream interface 124
    input m_axis_fifo_124_aclk,
    input m_axis_fifo_124_aresetn,
    output m_axis_fifo_124_tlast,
    output m_axis_fifo_124_tvalid,
    output [M_AXIS_FIFO_124_DMWIDTH/8-1:0] m_axis_fifo_124_tkeep,
    output [M_AXIS_FIFO_124_DMWIDTH/8-1:0] m_axis_fifo_124_tstrb,
    output [M_AXIS_FIFO_124_DMWIDTH-1:0] m_axis_fifo_124_tdata,
    input m_axis_fifo_124_tready,
    output ap_fifo_oarg_124_full_n,
    input [M_AXIS_FIFO_124_WIDTH-1:0] ap_fifo_oarg_124_din,
    input ap_fifo_oarg_124_write,
    //output FIFO to AXI-Stream interface 125
    input m_axis_fifo_125_aclk,
    input m_axis_fifo_125_aresetn,
    output m_axis_fifo_125_tlast,
    output m_axis_fifo_125_tvalid,
    output [M_AXIS_FIFO_125_DMWIDTH/8-1:0] m_axis_fifo_125_tkeep,
    output [M_AXIS_FIFO_125_DMWIDTH/8-1:0] m_axis_fifo_125_tstrb,
    output [M_AXIS_FIFO_125_DMWIDTH-1:0] m_axis_fifo_125_tdata,
    input m_axis_fifo_125_tready,
    output ap_fifo_oarg_125_full_n,
    input [M_AXIS_FIFO_125_WIDTH-1:0] ap_fifo_oarg_125_din,
    input ap_fifo_oarg_125_write,
    //output FIFO to AXI-Stream interface 126
    input m_axis_fifo_126_aclk,
    input m_axis_fifo_126_aresetn,
    output m_axis_fifo_126_tlast,
    output m_axis_fifo_126_tvalid,
    output [M_AXIS_FIFO_126_DMWIDTH/8-1:0] m_axis_fifo_126_tkeep,
    output [M_AXIS_FIFO_126_DMWIDTH/8-1:0] m_axis_fifo_126_tstrb,
    output [M_AXIS_FIFO_126_DMWIDTH-1:0] m_axis_fifo_126_tdata,
    input m_axis_fifo_126_tready,
    output ap_fifo_oarg_126_full_n,
    input [M_AXIS_FIFO_126_WIDTH-1:0] ap_fifo_oarg_126_din,
    input ap_fifo_oarg_126_write,
    //output FIFO to AXI-Stream interface 127
    input m_axis_fifo_127_aclk,
    input m_axis_fifo_127_aresetn,
    output m_axis_fifo_127_tlast,
    output m_axis_fifo_127_tvalid,
    output [M_AXIS_FIFO_127_DMWIDTH/8-1:0] m_axis_fifo_127_tkeep,
    output [M_AXIS_FIFO_127_DMWIDTH/8-1:0] m_axis_fifo_127_tstrb,
    output [M_AXIS_FIFO_127_DMWIDTH-1:0] m_axis_fifo_127_tdata,
    input m_axis_fifo_127_tready,
    output ap_fifo_oarg_127_full_n,
    input [M_AXIS_FIFO_127_WIDTH-1:0] ap_fifo_oarg_127_din,
    input ap_fifo_oarg_127_write,
    //-----------------------------------------------------
    //input AXI-Stream to BRAM interface 0
    input s_axis_bram_0_aclk,
    input s_axis_bram_0_aresetn,
    input s_axis_bram_0_tlast,
    input s_axis_bram_0_tvalid,
    input [S_AXIS_BRAM_0_DMWIDTH/8-1:0] s_axis_bram_0_tkeep,
    input [S_AXIS_BRAM_0_DMWIDTH/8-1:0] s_axis_bram_0_tstrb,
    input [S_AXIS_BRAM_0_DMWIDTH-1:0] s_axis_bram_0_tdata,
    output s_axis_bram_0_tready,
    input [S_AXIS_BRAM_0_ADDR_WIDTH-1:0] ap_bram_iarg_0_addr0,
    input [S_AXIS_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_din0,
    output [S_AXIS_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_dout0,
    input ap_bram_iarg_0_clk0,
    input ap_bram_iarg_0_rst0,
    input [S_AXIS_BRAM_0_WIDTH/8-1:0] ap_bram_iarg_0_we0,
    input ap_bram_iarg_0_en0,
    input [S_AXIS_BRAM_0_ADDR_WIDTH-1:0] ap_bram_iarg_0_addr1,
    input [S_AXIS_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_din1,
    output [S_AXIS_BRAM_0_WIDTH-1:0] ap_bram_iarg_0_dout1,
    input ap_bram_iarg_0_clk1,
    input ap_bram_iarg_0_rst1,
    input [S_AXIS_BRAM_0_WIDTH/8-1:0] ap_bram_iarg_0_we1,
    input ap_bram_iarg_0_en1,
    //input AXI-Stream to BRAM interface 1
    input s_axis_bram_1_aclk,
    input s_axis_bram_1_aresetn,
    input s_axis_bram_1_tlast,
    input s_axis_bram_1_tvalid,
    input [S_AXIS_BRAM_1_DMWIDTH/8-1:0] s_axis_bram_1_tkeep,
    input [S_AXIS_BRAM_1_DMWIDTH/8-1:0] s_axis_bram_1_tstrb,
    input [S_AXIS_BRAM_1_DMWIDTH-1:0] s_axis_bram_1_tdata,
    output s_axis_bram_1_tready,
    input [S_AXIS_BRAM_1_ADDR_WIDTH-1:0] ap_bram_iarg_1_addr0,
    input [S_AXIS_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_din0,
    output [S_AXIS_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_dout0,
    input ap_bram_iarg_1_clk0,
    input ap_bram_iarg_1_rst0,
    input [S_AXIS_BRAM_1_WIDTH/8-1:0] ap_bram_iarg_1_we0,
    input ap_bram_iarg_1_en0,
    input [S_AXIS_BRAM_1_ADDR_WIDTH-1:0] ap_bram_iarg_1_addr1,
    input [S_AXIS_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_din1,
    output [S_AXIS_BRAM_1_WIDTH-1:0] ap_bram_iarg_1_dout1,
    input ap_bram_iarg_1_clk1,
    input ap_bram_iarg_1_rst1,
    input [S_AXIS_BRAM_1_WIDTH/8-1:0] ap_bram_iarg_1_we1,
    input ap_bram_iarg_1_en1,
    //input AXI-Stream to BRAM interface 2
    input s_axis_bram_2_aclk,
    input s_axis_bram_2_aresetn,
    input s_axis_bram_2_tlast,
    input s_axis_bram_2_tvalid,
    input [S_AXIS_BRAM_2_DMWIDTH/8-1:0] s_axis_bram_2_tkeep,
    input [S_AXIS_BRAM_2_DMWIDTH/8-1:0] s_axis_bram_2_tstrb,
    input [S_AXIS_BRAM_2_DMWIDTH-1:0] s_axis_bram_2_tdata,
    output s_axis_bram_2_tready,
    input [S_AXIS_BRAM_2_ADDR_WIDTH-1:0] ap_bram_iarg_2_addr0,
    input [S_AXIS_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_din0,
    output [S_AXIS_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_dout0,
    input ap_bram_iarg_2_clk0,
    input ap_bram_iarg_2_rst0,
    input [S_AXIS_BRAM_2_WIDTH/8-1:0] ap_bram_iarg_2_we0,
    input ap_bram_iarg_2_en0,
    input [S_AXIS_BRAM_2_ADDR_WIDTH-1:0] ap_bram_iarg_2_addr1,
    input [S_AXIS_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_din1,
    output [S_AXIS_BRAM_2_WIDTH-1:0] ap_bram_iarg_2_dout1,
    input ap_bram_iarg_2_clk1,
    input ap_bram_iarg_2_rst1,
    input [S_AXIS_BRAM_2_WIDTH/8-1:0] ap_bram_iarg_2_we1,
    input ap_bram_iarg_2_en1,
    //input AXI-Stream to BRAM interface 3
    input s_axis_bram_3_aclk,
    input s_axis_bram_3_aresetn,
    input s_axis_bram_3_tlast,
    input s_axis_bram_3_tvalid,
    input [S_AXIS_BRAM_3_DMWIDTH/8-1:0] s_axis_bram_3_tkeep,
    input [S_AXIS_BRAM_3_DMWIDTH/8-1:0] s_axis_bram_3_tstrb,
    input [S_AXIS_BRAM_3_DMWIDTH-1:0] s_axis_bram_3_tdata,
    output s_axis_bram_3_tready,
    input [S_AXIS_BRAM_3_ADDR_WIDTH-1:0] ap_bram_iarg_3_addr0,
    input [S_AXIS_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_din0,
    output [S_AXIS_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_dout0,
    input ap_bram_iarg_3_clk0,
    input ap_bram_iarg_3_rst0,
    input [S_AXIS_BRAM_3_WIDTH/8-1:0] ap_bram_iarg_3_we0,
    input ap_bram_iarg_3_en0,
    input [S_AXIS_BRAM_3_ADDR_WIDTH-1:0] ap_bram_iarg_3_addr1,
    input [S_AXIS_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_din1,
    output [S_AXIS_BRAM_3_WIDTH-1:0] ap_bram_iarg_3_dout1,
    input ap_bram_iarg_3_clk1,
    input ap_bram_iarg_3_rst1,
    input [S_AXIS_BRAM_3_WIDTH/8-1:0] ap_bram_iarg_3_we1,
    input ap_bram_iarg_3_en1,
    //input AXI-Stream to BRAM interface 4
    input s_axis_bram_4_aclk,
    input s_axis_bram_4_aresetn,
    input s_axis_bram_4_tlast,
    input s_axis_bram_4_tvalid,
    input [S_AXIS_BRAM_4_DMWIDTH/8-1:0] s_axis_bram_4_tkeep,
    input [S_AXIS_BRAM_4_DMWIDTH/8-1:0] s_axis_bram_4_tstrb,
    input [S_AXIS_BRAM_4_DMWIDTH-1:0] s_axis_bram_4_tdata,
    output s_axis_bram_4_tready,
    input [S_AXIS_BRAM_4_ADDR_WIDTH-1:0] ap_bram_iarg_4_addr0,
    input [S_AXIS_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_din0,
    output [S_AXIS_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_dout0,
    input ap_bram_iarg_4_clk0,
    input ap_bram_iarg_4_rst0,
    input [S_AXIS_BRAM_4_WIDTH/8-1:0] ap_bram_iarg_4_we0,
    input ap_bram_iarg_4_en0,
    input [S_AXIS_BRAM_4_ADDR_WIDTH-1:0] ap_bram_iarg_4_addr1,
    input [S_AXIS_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_din1,
    output [S_AXIS_BRAM_4_WIDTH-1:0] ap_bram_iarg_4_dout1,
    input ap_bram_iarg_4_clk1,
    input ap_bram_iarg_4_rst1,
    input [S_AXIS_BRAM_4_WIDTH/8-1:0] ap_bram_iarg_4_we1,
    input ap_bram_iarg_4_en1,
    //input AXI-Stream to BRAM interface 5
    input s_axis_bram_5_aclk,
    input s_axis_bram_5_aresetn,
    input s_axis_bram_5_tlast,
    input s_axis_bram_5_tvalid,
    input [S_AXIS_BRAM_5_DMWIDTH/8-1:0] s_axis_bram_5_tkeep,
    input [S_AXIS_BRAM_5_DMWIDTH/8-1:0] s_axis_bram_5_tstrb,
    input [S_AXIS_BRAM_5_DMWIDTH-1:0] s_axis_bram_5_tdata,
    output s_axis_bram_5_tready,
    input [S_AXIS_BRAM_5_ADDR_WIDTH-1:0] ap_bram_iarg_5_addr0,
    input [S_AXIS_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_din0,
    output [S_AXIS_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_dout0,
    input ap_bram_iarg_5_clk0,
    input ap_bram_iarg_5_rst0,
    input [S_AXIS_BRAM_5_WIDTH/8-1:0] ap_bram_iarg_5_we0,
    input ap_bram_iarg_5_en0,
    input [S_AXIS_BRAM_5_ADDR_WIDTH-1:0] ap_bram_iarg_5_addr1,
    input [S_AXIS_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_din1,
    output [S_AXIS_BRAM_5_WIDTH-1:0] ap_bram_iarg_5_dout1,
    input ap_bram_iarg_5_clk1,
    input ap_bram_iarg_5_rst1,
    input [S_AXIS_BRAM_5_WIDTH/8-1:0] ap_bram_iarg_5_we1,
    input ap_bram_iarg_5_en1,
    //input AXI-Stream to BRAM interface 6
    input s_axis_bram_6_aclk,
    input s_axis_bram_6_aresetn,
    input s_axis_bram_6_tlast,
    input s_axis_bram_6_tvalid,
    input [S_AXIS_BRAM_6_DMWIDTH/8-1:0] s_axis_bram_6_tkeep,
    input [S_AXIS_BRAM_6_DMWIDTH/8-1:0] s_axis_bram_6_tstrb,
    input [S_AXIS_BRAM_6_DMWIDTH-1:0] s_axis_bram_6_tdata,
    output s_axis_bram_6_tready,
    input [S_AXIS_BRAM_6_ADDR_WIDTH-1:0] ap_bram_iarg_6_addr0,
    input [S_AXIS_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_din0,
    output [S_AXIS_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_dout0,
    input ap_bram_iarg_6_clk0,
    input ap_bram_iarg_6_rst0,
    input [S_AXIS_BRAM_6_WIDTH/8-1:0] ap_bram_iarg_6_we0,
    input ap_bram_iarg_6_en0,
    input [S_AXIS_BRAM_6_ADDR_WIDTH-1:0] ap_bram_iarg_6_addr1,
    input [S_AXIS_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_din1,
    output [S_AXIS_BRAM_6_WIDTH-1:0] ap_bram_iarg_6_dout1,
    input ap_bram_iarg_6_clk1,
    input ap_bram_iarg_6_rst1,
    input [S_AXIS_BRAM_6_WIDTH/8-1:0] ap_bram_iarg_6_we1,
    input ap_bram_iarg_6_en1,
    //input AXI-Stream to BRAM interface 7
    input s_axis_bram_7_aclk,
    input s_axis_bram_7_aresetn,
    input s_axis_bram_7_tlast,
    input s_axis_bram_7_tvalid,
    input [S_AXIS_BRAM_7_DMWIDTH/8-1:0] s_axis_bram_7_tkeep,
    input [S_AXIS_BRAM_7_DMWIDTH/8-1:0] s_axis_bram_7_tstrb,
    input [S_AXIS_BRAM_7_DMWIDTH-1:0] s_axis_bram_7_tdata,
    output s_axis_bram_7_tready,
    input [S_AXIS_BRAM_7_ADDR_WIDTH-1:0] ap_bram_iarg_7_addr0,
    input [S_AXIS_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_din0,
    output [S_AXIS_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_dout0,
    input ap_bram_iarg_7_clk0,
    input ap_bram_iarg_7_rst0,
    input [S_AXIS_BRAM_7_WIDTH/8-1:0] ap_bram_iarg_7_we0,
    input ap_bram_iarg_7_en0,
    input [S_AXIS_BRAM_7_ADDR_WIDTH-1:0] ap_bram_iarg_7_addr1,
    input [S_AXIS_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_din1,
    output [S_AXIS_BRAM_7_WIDTH-1:0] ap_bram_iarg_7_dout1,
    input ap_bram_iarg_7_clk1,
    input ap_bram_iarg_7_rst1,
    input [S_AXIS_BRAM_7_WIDTH/8-1:0] ap_bram_iarg_7_we1,
    input ap_bram_iarg_7_en1,
    //input AXI-Stream to BRAM interface 8
    input s_axis_bram_8_aclk,
    input s_axis_bram_8_aresetn,
    input s_axis_bram_8_tlast,
    input s_axis_bram_8_tvalid,
    input [S_AXIS_BRAM_8_DMWIDTH/8-1:0] s_axis_bram_8_tkeep,
    input [S_AXIS_BRAM_8_DMWIDTH/8-1:0] s_axis_bram_8_tstrb,
    input [S_AXIS_BRAM_8_DMWIDTH-1:0] s_axis_bram_8_tdata,
    output s_axis_bram_8_tready,
    input [S_AXIS_BRAM_8_ADDR_WIDTH-1:0] ap_bram_iarg_8_addr0,
    input [S_AXIS_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_din0,
    output [S_AXIS_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_dout0,
    input ap_bram_iarg_8_clk0,
    input ap_bram_iarg_8_rst0,
    input [S_AXIS_BRAM_8_WIDTH/8-1:0] ap_bram_iarg_8_we0,
    input ap_bram_iarg_8_en0,
    input [S_AXIS_BRAM_8_ADDR_WIDTH-1:0] ap_bram_iarg_8_addr1,
    input [S_AXIS_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_din1,
    output [S_AXIS_BRAM_8_WIDTH-1:0] ap_bram_iarg_8_dout1,
    input ap_bram_iarg_8_clk1,
    input ap_bram_iarg_8_rst1,
    input [S_AXIS_BRAM_8_WIDTH/8-1:0] ap_bram_iarg_8_we1,
    input ap_bram_iarg_8_en1,
    //input AXI-Stream to BRAM interface 9
    input s_axis_bram_9_aclk,
    input s_axis_bram_9_aresetn,
    input s_axis_bram_9_tlast,
    input s_axis_bram_9_tvalid,
    input [S_AXIS_BRAM_9_DMWIDTH/8-1:0] s_axis_bram_9_tkeep,
    input [S_AXIS_BRAM_9_DMWIDTH/8-1:0] s_axis_bram_9_tstrb,
    input [S_AXIS_BRAM_9_DMWIDTH-1:0] s_axis_bram_9_tdata,
    output s_axis_bram_9_tready,
    input [S_AXIS_BRAM_9_ADDR_WIDTH-1:0] ap_bram_iarg_9_addr0,
    input [S_AXIS_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_din0,
    output [S_AXIS_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_dout0,
    input ap_bram_iarg_9_clk0,
    input ap_bram_iarg_9_rst0,
    input [S_AXIS_BRAM_9_WIDTH/8-1:0] ap_bram_iarg_9_we0,
    input ap_bram_iarg_9_en0,
    input [S_AXIS_BRAM_9_ADDR_WIDTH-1:0] ap_bram_iarg_9_addr1,
    input [S_AXIS_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_din1,
    output [S_AXIS_BRAM_9_WIDTH-1:0] ap_bram_iarg_9_dout1,
    input ap_bram_iarg_9_clk1,
    input ap_bram_iarg_9_rst1,
    input [S_AXIS_BRAM_9_WIDTH/8-1:0] ap_bram_iarg_9_we1,
    input ap_bram_iarg_9_en1,
    //input AXI-Stream to BRAM interface 10
    input s_axis_bram_10_aclk,
    input s_axis_bram_10_aresetn,
    input s_axis_bram_10_tlast,
    input s_axis_bram_10_tvalid,
    input [S_AXIS_BRAM_10_DMWIDTH/8-1:0] s_axis_bram_10_tkeep,
    input [S_AXIS_BRAM_10_DMWIDTH/8-1:0] s_axis_bram_10_tstrb,
    input [S_AXIS_BRAM_10_DMWIDTH-1:0] s_axis_bram_10_tdata,
    output s_axis_bram_10_tready,
    input [S_AXIS_BRAM_10_ADDR_WIDTH-1:0] ap_bram_iarg_10_addr0,
    input [S_AXIS_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_din0,
    output [S_AXIS_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_dout0,
    input ap_bram_iarg_10_clk0,
    input ap_bram_iarg_10_rst0,
    input [S_AXIS_BRAM_10_WIDTH/8-1:0] ap_bram_iarg_10_we0,
    input ap_bram_iarg_10_en0,
    input [S_AXIS_BRAM_10_ADDR_WIDTH-1:0] ap_bram_iarg_10_addr1,
    input [S_AXIS_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_din1,
    output [S_AXIS_BRAM_10_WIDTH-1:0] ap_bram_iarg_10_dout1,
    input ap_bram_iarg_10_clk1,
    input ap_bram_iarg_10_rst1,
    input [S_AXIS_BRAM_10_WIDTH/8-1:0] ap_bram_iarg_10_we1,
    input ap_bram_iarg_10_en1,
    //input AXI-Stream to BRAM interface 11
    input s_axis_bram_11_aclk,
    input s_axis_bram_11_aresetn,
    input s_axis_bram_11_tlast,
    input s_axis_bram_11_tvalid,
    input [S_AXIS_BRAM_11_DMWIDTH/8-1:0] s_axis_bram_11_tkeep,
    input [S_AXIS_BRAM_11_DMWIDTH/8-1:0] s_axis_bram_11_tstrb,
    input [S_AXIS_BRAM_11_DMWIDTH-1:0] s_axis_bram_11_tdata,
    output s_axis_bram_11_tready,
    input [S_AXIS_BRAM_11_ADDR_WIDTH-1:0] ap_bram_iarg_11_addr0,
    input [S_AXIS_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_din0,
    output [S_AXIS_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_dout0,
    input ap_bram_iarg_11_clk0,
    input ap_bram_iarg_11_rst0,
    input [S_AXIS_BRAM_11_WIDTH/8-1:0] ap_bram_iarg_11_we0,
    input ap_bram_iarg_11_en0,
    input [S_AXIS_BRAM_11_ADDR_WIDTH-1:0] ap_bram_iarg_11_addr1,
    input [S_AXIS_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_din1,
    output [S_AXIS_BRAM_11_WIDTH-1:0] ap_bram_iarg_11_dout1,
    input ap_bram_iarg_11_clk1,
    input ap_bram_iarg_11_rst1,
    input [S_AXIS_BRAM_11_WIDTH/8-1:0] ap_bram_iarg_11_we1,
    input ap_bram_iarg_11_en1,
    //input AXI-Stream to BRAM interface 12
    input s_axis_bram_12_aclk,
    input s_axis_bram_12_aresetn,
    input s_axis_bram_12_tlast,
    input s_axis_bram_12_tvalid,
    input [S_AXIS_BRAM_12_DMWIDTH/8-1:0] s_axis_bram_12_tkeep,
    input [S_AXIS_BRAM_12_DMWIDTH/8-1:0] s_axis_bram_12_tstrb,
    input [S_AXIS_BRAM_12_DMWIDTH-1:0] s_axis_bram_12_tdata,
    output s_axis_bram_12_tready,
    input [S_AXIS_BRAM_12_ADDR_WIDTH-1:0] ap_bram_iarg_12_addr0,
    input [S_AXIS_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_din0,
    output [S_AXIS_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_dout0,
    input ap_bram_iarg_12_clk0,
    input ap_bram_iarg_12_rst0,
    input [S_AXIS_BRAM_12_WIDTH/8-1:0] ap_bram_iarg_12_we0,
    input ap_bram_iarg_12_en0,
    input [S_AXIS_BRAM_12_ADDR_WIDTH-1:0] ap_bram_iarg_12_addr1,
    input [S_AXIS_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_din1,
    output [S_AXIS_BRAM_12_WIDTH-1:0] ap_bram_iarg_12_dout1,
    input ap_bram_iarg_12_clk1,
    input ap_bram_iarg_12_rst1,
    input [S_AXIS_BRAM_12_WIDTH/8-1:0] ap_bram_iarg_12_we1,
    input ap_bram_iarg_12_en1,
    //input AXI-Stream to BRAM interface 13
    input s_axis_bram_13_aclk,
    input s_axis_bram_13_aresetn,
    input s_axis_bram_13_tlast,
    input s_axis_bram_13_tvalid,
    input [S_AXIS_BRAM_13_DMWIDTH/8-1:0] s_axis_bram_13_tkeep,
    input [S_AXIS_BRAM_13_DMWIDTH/8-1:0] s_axis_bram_13_tstrb,
    input [S_AXIS_BRAM_13_DMWIDTH-1:0] s_axis_bram_13_tdata,
    output s_axis_bram_13_tready,
    input [S_AXIS_BRAM_13_ADDR_WIDTH-1:0] ap_bram_iarg_13_addr0,
    input [S_AXIS_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_din0,
    output [S_AXIS_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_dout0,
    input ap_bram_iarg_13_clk0,
    input ap_bram_iarg_13_rst0,
    input [S_AXIS_BRAM_13_WIDTH/8-1:0] ap_bram_iarg_13_we0,
    input ap_bram_iarg_13_en0,
    input [S_AXIS_BRAM_13_ADDR_WIDTH-1:0] ap_bram_iarg_13_addr1,
    input [S_AXIS_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_din1,
    output [S_AXIS_BRAM_13_WIDTH-1:0] ap_bram_iarg_13_dout1,
    input ap_bram_iarg_13_clk1,
    input ap_bram_iarg_13_rst1,
    input [S_AXIS_BRAM_13_WIDTH/8-1:0] ap_bram_iarg_13_we1,
    input ap_bram_iarg_13_en1,
    //input AXI-Stream to BRAM interface 14
    input s_axis_bram_14_aclk,
    input s_axis_bram_14_aresetn,
    input s_axis_bram_14_tlast,
    input s_axis_bram_14_tvalid,
    input [S_AXIS_BRAM_14_DMWIDTH/8-1:0] s_axis_bram_14_tkeep,
    input [S_AXIS_BRAM_14_DMWIDTH/8-1:0] s_axis_bram_14_tstrb,
    input [S_AXIS_BRAM_14_DMWIDTH-1:0] s_axis_bram_14_tdata,
    output s_axis_bram_14_tready,
    input [S_AXIS_BRAM_14_ADDR_WIDTH-1:0] ap_bram_iarg_14_addr0,
    input [S_AXIS_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_din0,
    output [S_AXIS_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_dout0,
    input ap_bram_iarg_14_clk0,
    input ap_bram_iarg_14_rst0,
    input [S_AXIS_BRAM_14_WIDTH/8-1:0] ap_bram_iarg_14_we0,
    input ap_bram_iarg_14_en0,
    input [S_AXIS_BRAM_14_ADDR_WIDTH-1:0] ap_bram_iarg_14_addr1,
    input [S_AXIS_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_din1,
    output [S_AXIS_BRAM_14_WIDTH-1:0] ap_bram_iarg_14_dout1,
    input ap_bram_iarg_14_clk1,
    input ap_bram_iarg_14_rst1,
    input [S_AXIS_BRAM_14_WIDTH/8-1:0] ap_bram_iarg_14_we1,
    input ap_bram_iarg_14_en1,
    //input AXI-Stream to BRAM interface 15
    input s_axis_bram_15_aclk,
    input s_axis_bram_15_aresetn,
    input s_axis_bram_15_tlast,
    input s_axis_bram_15_tvalid,
    input [S_AXIS_BRAM_15_DMWIDTH/8-1:0] s_axis_bram_15_tkeep,
    input [S_AXIS_BRAM_15_DMWIDTH/8-1:0] s_axis_bram_15_tstrb,
    input [S_AXIS_BRAM_15_DMWIDTH-1:0] s_axis_bram_15_tdata,
    output s_axis_bram_15_tready,
    input [S_AXIS_BRAM_15_ADDR_WIDTH-1:0] ap_bram_iarg_15_addr0,
    input [S_AXIS_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_din0,
    output [S_AXIS_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_dout0,
    input ap_bram_iarg_15_clk0,
    input ap_bram_iarg_15_rst0,
    input [S_AXIS_BRAM_15_WIDTH/8-1:0] ap_bram_iarg_15_we0,
    input ap_bram_iarg_15_en0,
    input [S_AXIS_BRAM_15_ADDR_WIDTH-1:0] ap_bram_iarg_15_addr1,
    input [S_AXIS_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_din1,
    output [S_AXIS_BRAM_15_WIDTH-1:0] ap_bram_iarg_15_dout1,
    input ap_bram_iarg_15_clk1,
    input ap_bram_iarg_15_rst1,
    input [S_AXIS_BRAM_15_WIDTH/8-1:0] ap_bram_iarg_15_we1,
    input ap_bram_iarg_15_en1,
    //input AXI-Stream to BRAM interface 16
    input s_axis_bram_16_aclk,
    input s_axis_bram_16_aresetn,
    input s_axis_bram_16_tlast,
    input s_axis_bram_16_tvalid,
    input [S_AXIS_BRAM_16_DMWIDTH/8-1:0] s_axis_bram_16_tkeep,
    input [S_AXIS_BRAM_16_DMWIDTH/8-1:0] s_axis_bram_16_tstrb,
    input [S_AXIS_BRAM_16_DMWIDTH-1:0] s_axis_bram_16_tdata,
    output s_axis_bram_16_tready,
    input [S_AXIS_BRAM_16_ADDR_WIDTH-1:0] ap_bram_iarg_16_addr0,
    input [S_AXIS_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_din0,
    output [S_AXIS_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_dout0,
    input ap_bram_iarg_16_clk0,
    input ap_bram_iarg_16_rst0,
    input [S_AXIS_BRAM_16_WIDTH/8-1:0] ap_bram_iarg_16_we0,
    input ap_bram_iarg_16_en0,
    input [S_AXIS_BRAM_16_ADDR_WIDTH-1:0] ap_bram_iarg_16_addr1,
    input [S_AXIS_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_din1,
    output [S_AXIS_BRAM_16_WIDTH-1:0] ap_bram_iarg_16_dout1,
    input ap_bram_iarg_16_clk1,
    input ap_bram_iarg_16_rst1,
    input [S_AXIS_BRAM_16_WIDTH/8-1:0] ap_bram_iarg_16_we1,
    input ap_bram_iarg_16_en1,
    //input AXI-Stream to BRAM interface 17
    input s_axis_bram_17_aclk,
    input s_axis_bram_17_aresetn,
    input s_axis_bram_17_tlast,
    input s_axis_bram_17_tvalid,
    input [S_AXIS_BRAM_17_DMWIDTH/8-1:0] s_axis_bram_17_tkeep,
    input [S_AXIS_BRAM_17_DMWIDTH/8-1:0] s_axis_bram_17_tstrb,
    input [S_AXIS_BRAM_17_DMWIDTH-1:0] s_axis_bram_17_tdata,
    output s_axis_bram_17_tready,
    input [S_AXIS_BRAM_17_ADDR_WIDTH-1:0] ap_bram_iarg_17_addr0,
    input [S_AXIS_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_din0,
    output [S_AXIS_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_dout0,
    input ap_bram_iarg_17_clk0,
    input ap_bram_iarg_17_rst0,
    input [S_AXIS_BRAM_17_WIDTH/8-1:0] ap_bram_iarg_17_we0,
    input ap_bram_iarg_17_en0,
    input [S_AXIS_BRAM_17_ADDR_WIDTH-1:0] ap_bram_iarg_17_addr1,
    input [S_AXIS_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_din1,
    output [S_AXIS_BRAM_17_WIDTH-1:0] ap_bram_iarg_17_dout1,
    input ap_bram_iarg_17_clk1,
    input ap_bram_iarg_17_rst1,
    input [S_AXIS_BRAM_17_WIDTH/8-1:0] ap_bram_iarg_17_we1,
    input ap_bram_iarg_17_en1,
    //input AXI-Stream to BRAM interface 18
    input s_axis_bram_18_aclk,
    input s_axis_bram_18_aresetn,
    input s_axis_bram_18_tlast,
    input s_axis_bram_18_tvalid,
    input [S_AXIS_BRAM_18_DMWIDTH/8-1:0] s_axis_bram_18_tkeep,
    input [S_AXIS_BRAM_18_DMWIDTH/8-1:0] s_axis_bram_18_tstrb,
    input [S_AXIS_BRAM_18_DMWIDTH-1:0] s_axis_bram_18_tdata,
    output s_axis_bram_18_tready,
    input [S_AXIS_BRAM_18_ADDR_WIDTH-1:0] ap_bram_iarg_18_addr0,
    input [S_AXIS_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_din0,
    output [S_AXIS_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_dout0,
    input ap_bram_iarg_18_clk0,
    input ap_bram_iarg_18_rst0,
    input [S_AXIS_BRAM_18_WIDTH/8-1:0] ap_bram_iarg_18_we0,
    input ap_bram_iarg_18_en0,
    input [S_AXIS_BRAM_18_ADDR_WIDTH-1:0] ap_bram_iarg_18_addr1,
    input [S_AXIS_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_din1,
    output [S_AXIS_BRAM_18_WIDTH-1:0] ap_bram_iarg_18_dout1,
    input ap_bram_iarg_18_clk1,
    input ap_bram_iarg_18_rst1,
    input [S_AXIS_BRAM_18_WIDTH/8-1:0] ap_bram_iarg_18_we1,
    input ap_bram_iarg_18_en1,
    //input AXI-Stream to BRAM interface 19
    input s_axis_bram_19_aclk,
    input s_axis_bram_19_aresetn,
    input s_axis_bram_19_tlast,
    input s_axis_bram_19_tvalid,
    input [S_AXIS_BRAM_19_DMWIDTH/8-1:0] s_axis_bram_19_tkeep,
    input [S_AXIS_BRAM_19_DMWIDTH/8-1:0] s_axis_bram_19_tstrb,
    input [S_AXIS_BRAM_19_DMWIDTH-1:0] s_axis_bram_19_tdata,
    output s_axis_bram_19_tready,
    input [S_AXIS_BRAM_19_ADDR_WIDTH-1:0] ap_bram_iarg_19_addr0,
    input [S_AXIS_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_din0,
    output [S_AXIS_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_dout0,
    input ap_bram_iarg_19_clk0,
    input ap_bram_iarg_19_rst0,
    input [S_AXIS_BRAM_19_WIDTH/8-1:0] ap_bram_iarg_19_we0,
    input ap_bram_iarg_19_en0,
    input [S_AXIS_BRAM_19_ADDR_WIDTH-1:0] ap_bram_iarg_19_addr1,
    input [S_AXIS_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_din1,
    output [S_AXIS_BRAM_19_WIDTH-1:0] ap_bram_iarg_19_dout1,
    input ap_bram_iarg_19_clk1,
    input ap_bram_iarg_19_rst1,
    input [S_AXIS_BRAM_19_WIDTH/8-1:0] ap_bram_iarg_19_we1,
    input ap_bram_iarg_19_en1,
    //input AXI-Stream to BRAM interface 20
    input s_axis_bram_20_aclk,
    input s_axis_bram_20_aresetn,
    input s_axis_bram_20_tlast,
    input s_axis_bram_20_tvalid,
    input [S_AXIS_BRAM_20_DMWIDTH/8-1:0] s_axis_bram_20_tkeep,
    input [S_AXIS_BRAM_20_DMWIDTH/8-1:0] s_axis_bram_20_tstrb,
    input [S_AXIS_BRAM_20_DMWIDTH-1:0] s_axis_bram_20_tdata,
    output s_axis_bram_20_tready,
    input [S_AXIS_BRAM_20_ADDR_WIDTH-1:0] ap_bram_iarg_20_addr0,
    input [S_AXIS_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_din0,
    output [S_AXIS_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_dout0,
    input ap_bram_iarg_20_clk0,
    input ap_bram_iarg_20_rst0,
    input [S_AXIS_BRAM_20_WIDTH/8-1:0] ap_bram_iarg_20_we0,
    input ap_bram_iarg_20_en0,
    input [S_AXIS_BRAM_20_ADDR_WIDTH-1:0] ap_bram_iarg_20_addr1,
    input [S_AXIS_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_din1,
    output [S_AXIS_BRAM_20_WIDTH-1:0] ap_bram_iarg_20_dout1,
    input ap_bram_iarg_20_clk1,
    input ap_bram_iarg_20_rst1,
    input [S_AXIS_BRAM_20_WIDTH/8-1:0] ap_bram_iarg_20_we1,
    input ap_bram_iarg_20_en1,
    //input AXI-Stream to BRAM interface 21
    input s_axis_bram_21_aclk,
    input s_axis_bram_21_aresetn,
    input s_axis_bram_21_tlast,
    input s_axis_bram_21_tvalid,
    input [S_AXIS_BRAM_21_DMWIDTH/8-1:0] s_axis_bram_21_tkeep,
    input [S_AXIS_BRAM_21_DMWIDTH/8-1:0] s_axis_bram_21_tstrb,
    input [S_AXIS_BRAM_21_DMWIDTH-1:0] s_axis_bram_21_tdata,
    output s_axis_bram_21_tready,
    input [S_AXIS_BRAM_21_ADDR_WIDTH-1:0] ap_bram_iarg_21_addr0,
    input [S_AXIS_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_din0,
    output [S_AXIS_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_dout0,
    input ap_bram_iarg_21_clk0,
    input ap_bram_iarg_21_rst0,
    input [S_AXIS_BRAM_21_WIDTH/8-1:0] ap_bram_iarg_21_we0,
    input ap_bram_iarg_21_en0,
    input [S_AXIS_BRAM_21_ADDR_WIDTH-1:0] ap_bram_iarg_21_addr1,
    input [S_AXIS_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_din1,
    output [S_AXIS_BRAM_21_WIDTH-1:0] ap_bram_iarg_21_dout1,
    input ap_bram_iarg_21_clk1,
    input ap_bram_iarg_21_rst1,
    input [S_AXIS_BRAM_21_WIDTH/8-1:0] ap_bram_iarg_21_we1,
    input ap_bram_iarg_21_en1,
    //input AXI-Stream to BRAM interface 22
    input s_axis_bram_22_aclk,
    input s_axis_bram_22_aresetn,
    input s_axis_bram_22_tlast,
    input s_axis_bram_22_tvalid,
    input [S_AXIS_BRAM_22_DMWIDTH/8-1:0] s_axis_bram_22_tkeep,
    input [S_AXIS_BRAM_22_DMWIDTH/8-1:0] s_axis_bram_22_tstrb,
    input [S_AXIS_BRAM_22_DMWIDTH-1:0] s_axis_bram_22_tdata,
    output s_axis_bram_22_tready,
    input [S_AXIS_BRAM_22_ADDR_WIDTH-1:0] ap_bram_iarg_22_addr0,
    input [S_AXIS_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_din0,
    output [S_AXIS_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_dout0,
    input ap_bram_iarg_22_clk0,
    input ap_bram_iarg_22_rst0,
    input [S_AXIS_BRAM_22_WIDTH/8-1:0] ap_bram_iarg_22_we0,
    input ap_bram_iarg_22_en0,
    input [S_AXIS_BRAM_22_ADDR_WIDTH-1:0] ap_bram_iarg_22_addr1,
    input [S_AXIS_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_din1,
    output [S_AXIS_BRAM_22_WIDTH-1:0] ap_bram_iarg_22_dout1,
    input ap_bram_iarg_22_clk1,
    input ap_bram_iarg_22_rst1,
    input [S_AXIS_BRAM_22_WIDTH/8-1:0] ap_bram_iarg_22_we1,
    input ap_bram_iarg_22_en1,
    //input AXI-Stream to BRAM interface 23
    input s_axis_bram_23_aclk,
    input s_axis_bram_23_aresetn,
    input s_axis_bram_23_tlast,
    input s_axis_bram_23_tvalid,
    input [S_AXIS_BRAM_23_DMWIDTH/8-1:0] s_axis_bram_23_tkeep,
    input [S_AXIS_BRAM_23_DMWIDTH/8-1:0] s_axis_bram_23_tstrb,
    input [S_AXIS_BRAM_23_DMWIDTH-1:0] s_axis_bram_23_tdata,
    output s_axis_bram_23_tready,
    input [S_AXIS_BRAM_23_ADDR_WIDTH-1:0] ap_bram_iarg_23_addr0,
    input [S_AXIS_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_din0,
    output [S_AXIS_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_dout0,
    input ap_bram_iarg_23_clk0,
    input ap_bram_iarg_23_rst0,
    input [S_AXIS_BRAM_23_WIDTH/8-1:0] ap_bram_iarg_23_we0,
    input ap_bram_iarg_23_en0,
    input [S_AXIS_BRAM_23_ADDR_WIDTH-1:0] ap_bram_iarg_23_addr1,
    input [S_AXIS_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_din1,
    output [S_AXIS_BRAM_23_WIDTH-1:0] ap_bram_iarg_23_dout1,
    input ap_bram_iarg_23_clk1,
    input ap_bram_iarg_23_rst1,
    input [S_AXIS_BRAM_23_WIDTH/8-1:0] ap_bram_iarg_23_we1,
    input ap_bram_iarg_23_en1,
    //input AXI-Stream to BRAM interface 24
    input s_axis_bram_24_aclk,
    input s_axis_bram_24_aresetn,
    input s_axis_bram_24_tlast,
    input s_axis_bram_24_tvalid,
    input [S_AXIS_BRAM_24_DMWIDTH/8-1:0] s_axis_bram_24_tkeep,
    input [S_AXIS_BRAM_24_DMWIDTH/8-1:0] s_axis_bram_24_tstrb,
    input [S_AXIS_BRAM_24_DMWIDTH-1:0] s_axis_bram_24_tdata,
    output s_axis_bram_24_tready,
    input [S_AXIS_BRAM_24_ADDR_WIDTH-1:0] ap_bram_iarg_24_addr0,
    input [S_AXIS_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_din0,
    output [S_AXIS_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_dout0,
    input ap_bram_iarg_24_clk0,
    input ap_bram_iarg_24_rst0,
    input [S_AXIS_BRAM_24_WIDTH/8-1:0] ap_bram_iarg_24_we0,
    input ap_bram_iarg_24_en0,
    input [S_AXIS_BRAM_24_ADDR_WIDTH-1:0] ap_bram_iarg_24_addr1,
    input [S_AXIS_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_din1,
    output [S_AXIS_BRAM_24_WIDTH-1:0] ap_bram_iarg_24_dout1,
    input ap_bram_iarg_24_clk1,
    input ap_bram_iarg_24_rst1,
    input [S_AXIS_BRAM_24_WIDTH/8-1:0] ap_bram_iarg_24_we1,
    input ap_bram_iarg_24_en1,
    //input AXI-Stream to BRAM interface 25
    input s_axis_bram_25_aclk,
    input s_axis_bram_25_aresetn,
    input s_axis_bram_25_tlast,
    input s_axis_bram_25_tvalid,
    input [S_AXIS_BRAM_25_DMWIDTH/8-1:0] s_axis_bram_25_tkeep,
    input [S_AXIS_BRAM_25_DMWIDTH/8-1:0] s_axis_bram_25_tstrb,
    input [S_AXIS_BRAM_25_DMWIDTH-1:0] s_axis_bram_25_tdata,
    output s_axis_bram_25_tready,
    input [S_AXIS_BRAM_25_ADDR_WIDTH-1:0] ap_bram_iarg_25_addr0,
    input [S_AXIS_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_din0,
    output [S_AXIS_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_dout0,
    input ap_bram_iarg_25_clk0,
    input ap_bram_iarg_25_rst0,
    input [S_AXIS_BRAM_25_WIDTH/8-1:0] ap_bram_iarg_25_we0,
    input ap_bram_iarg_25_en0,
    input [S_AXIS_BRAM_25_ADDR_WIDTH-1:0] ap_bram_iarg_25_addr1,
    input [S_AXIS_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_din1,
    output [S_AXIS_BRAM_25_WIDTH-1:0] ap_bram_iarg_25_dout1,
    input ap_bram_iarg_25_clk1,
    input ap_bram_iarg_25_rst1,
    input [S_AXIS_BRAM_25_WIDTH/8-1:0] ap_bram_iarg_25_we1,
    input ap_bram_iarg_25_en1,
    //input AXI-Stream to BRAM interface 26
    input s_axis_bram_26_aclk,
    input s_axis_bram_26_aresetn,
    input s_axis_bram_26_tlast,
    input s_axis_bram_26_tvalid,
    input [S_AXIS_BRAM_26_DMWIDTH/8-1:0] s_axis_bram_26_tkeep,
    input [S_AXIS_BRAM_26_DMWIDTH/8-1:0] s_axis_bram_26_tstrb,
    input [S_AXIS_BRAM_26_DMWIDTH-1:0] s_axis_bram_26_tdata,
    output s_axis_bram_26_tready,
    input [S_AXIS_BRAM_26_ADDR_WIDTH-1:0] ap_bram_iarg_26_addr0,
    input [S_AXIS_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_din0,
    output [S_AXIS_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_dout0,
    input ap_bram_iarg_26_clk0,
    input ap_bram_iarg_26_rst0,
    input [S_AXIS_BRAM_26_WIDTH/8-1:0] ap_bram_iarg_26_we0,
    input ap_bram_iarg_26_en0,
    input [S_AXIS_BRAM_26_ADDR_WIDTH-1:0] ap_bram_iarg_26_addr1,
    input [S_AXIS_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_din1,
    output [S_AXIS_BRAM_26_WIDTH-1:0] ap_bram_iarg_26_dout1,
    input ap_bram_iarg_26_clk1,
    input ap_bram_iarg_26_rst1,
    input [S_AXIS_BRAM_26_WIDTH/8-1:0] ap_bram_iarg_26_we1,
    input ap_bram_iarg_26_en1,
    //input AXI-Stream to BRAM interface 27
    input s_axis_bram_27_aclk,
    input s_axis_bram_27_aresetn,
    input s_axis_bram_27_tlast,
    input s_axis_bram_27_tvalid,
    input [S_AXIS_BRAM_27_DMWIDTH/8-1:0] s_axis_bram_27_tkeep,
    input [S_AXIS_BRAM_27_DMWIDTH/8-1:0] s_axis_bram_27_tstrb,
    input [S_AXIS_BRAM_27_DMWIDTH-1:0] s_axis_bram_27_tdata,
    output s_axis_bram_27_tready,
    input [S_AXIS_BRAM_27_ADDR_WIDTH-1:0] ap_bram_iarg_27_addr0,
    input [S_AXIS_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_din0,
    output [S_AXIS_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_dout0,
    input ap_bram_iarg_27_clk0,
    input ap_bram_iarg_27_rst0,
    input [S_AXIS_BRAM_27_WIDTH/8-1:0] ap_bram_iarg_27_we0,
    input ap_bram_iarg_27_en0,
    input [S_AXIS_BRAM_27_ADDR_WIDTH-1:0] ap_bram_iarg_27_addr1,
    input [S_AXIS_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_din1,
    output [S_AXIS_BRAM_27_WIDTH-1:0] ap_bram_iarg_27_dout1,
    input ap_bram_iarg_27_clk1,
    input ap_bram_iarg_27_rst1,
    input [S_AXIS_BRAM_27_WIDTH/8-1:0] ap_bram_iarg_27_we1,
    input ap_bram_iarg_27_en1,
    //input AXI-Stream to BRAM interface 28
    input s_axis_bram_28_aclk,
    input s_axis_bram_28_aresetn,
    input s_axis_bram_28_tlast,
    input s_axis_bram_28_tvalid,
    input [S_AXIS_BRAM_28_DMWIDTH/8-1:0] s_axis_bram_28_tkeep,
    input [S_AXIS_BRAM_28_DMWIDTH/8-1:0] s_axis_bram_28_tstrb,
    input [S_AXIS_BRAM_28_DMWIDTH-1:0] s_axis_bram_28_tdata,
    output s_axis_bram_28_tready,
    input [S_AXIS_BRAM_28_ADDR_WIDTH-1:0] ap_bram_iarg_28_addr0,
    input [S_AXIS_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_din0,
    output [S_AXIS_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_dout0,
    input ap_bram_iarg_28_clk0,
    input ap_bram_iarg_28_rst0,
    input [S_AXIS_BRAM_28_WIDTH/8-1:0] ap_bram_iarg_28_we0,
    input ap_bram_iarg_28_en0,
    input [S_AXIS_BRAM_28_ADDR_WIDTH-1:0] ap_bram_iarg_28_addr1,
    input [S_AXIS_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_din1,
    output [S_AXIS_BRAM_28_WIDTH-1:0] ap_bram_iarg_28_dout1,
    input ap_bram_iarg_28_clk1,
    input ap_bram_iarg_28_rst1,
    input [S_AXIS_BRAM_28_WIDTH/8-1:0] ap_bram_iarg_28_we1,
    input ap_bram_iarg_28_en1,
    //input AXI-Stream to BRAM interface 29
    input s_axis_bram_29_aclk,
    input s_axis_bram_29_aresetn,
    input s_axis_bram_29_tlast,
    input s_axis_bram_29_tvalid,
    input [S_AXIS_BRAM_29_DMWIDTH/8-1:0] s_axis_bram_29_tkeep,
    input [S_AXIS_BRAM_29_DMWIDTH/8-1:0] s_axis_bram_29_tstrb,
    input [S_AXIS_BRAM_29_DMWIDTH-1:0] s_axis_bram_29_tdata,
    output s_axis_bram_29_tready,
    input [S_AXIS_BRAM_29_ADDR_WIDTH-1:0] ap_bram_iarg_29_addr0,
    input [S_AXIS_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_din0,
    output [S_AXIS_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_dout0,
    input ap_bram_iarg_29_clk0,
    input ap_bram_iarg_29_rst0,
    input [S_AXIS_BRAM_29_WIDTH/8-1:0] ap_bram_iarg_29_we0,
    input ap_bram_iarg_29_en0,
    input [S_AXIS_BRAM_29_ADDR_WIDTH-1:0] ap_bram_iarg_29_addr1,
    input [S_AXIS_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_din1,
    output [S_AXIS_BRAM_29_WIDTH-1:0] ap_bram_iarg_29_dout1,
    input ap_bram_iarg_29_clk1,
    input ap_bram_iarg_29_rst1,
    input [S_AXIS_BRAM_29_WIDTH/8-1:0] ap_bram_iarg_29_we1,
    input ap_bram_iarg_29_en1,
    //input AXI-Stream to BRAM interface 30
    input s_axis_bram_30_aclk,
    input s_axis_bram_30_aresetn,
    input s_axis_bram_30_tlast,
    input s_axis_bram_30_tvalid,
    input [S_AXIS_BRAM_30_DMWIDTH/8-1:0] s_axis_bram_30_tkeep,
    input [S_AXIS_BRAM_30_DMWIDTH/8-1:0] s_axis_bram_30_tstrb,
    input [S_AXIS_BRAM_30_DMWIDTH-1:0] s_axis_bram_30_tdata,
    output s_axis_bram_30_tready,
    input [S_AXIS_BRAM_30_ADDR_WIDTH-1:0] ap_bram_iarg_30_addr0,
    input [S_AXIS_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_din0,
    output [S_AXIS_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_dout0,
    input ap_bram_iarg_30_clk0,
    input ap_bram_iarg_30_rst0,
    input [S_AXIS_BRAM_30_WIDTH/8-1:0] ap_bram_iarg_30_we0,
    input ap_bram_iarg_30_en0,
    input [S_AXIS_BRAM_30_ADDR_WIDTH-1:0] ap_bram_iarg_30_addr1,
    input [S_AXIS_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_din1,
    output [S_AXIS_BRAM_30_WIDTH-1:0] ap_bram_iarg_30_dout1,
    input ap_bram_iarg_30_clk1,
    input ap_bram_iarg_30_rst1,
    input [S_AXIS_BRAM_30_WIDTH/8-1:0] ap_bram_iarg_30_we1,
    input ap_bram_iarg_30_en1,
    //input AXI-Stream to BRAM interface 31
    input s_axis_bram_31_aclk,
    input s_axis_bram_31_aresetn,
    input s_axis_bram_31_tlast,
    input s_axis_bram_31_tvalid,
    input [S_AXIS_BRAM_31_DMWIDTH/8-1:0] s_axis_bram_31_tkeep,
    input [S_AXIS_BRAM_31_DMWIDTH/8-1:0] s_axis_bram_31_tstrb,
    input [S_AXIS_BRAM_31_DMWIDTH-1:0] s_axis_bram_31_tdata,
    output s_axis_bram_31_tready,
    input [S_AXIS_BRAM_31_ADDR_WIDTH-1:0] ap_bram_iarg_31_addr0,
    input [S_AXIS_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_din0,
    output [S_AXIS_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_dout0,
    input ap_bram_iarg_31_clk0,
    input ap_bram_iarg_31_rst0,
    input [S_AXIS_BRAM_31_WIDTH/8-1:0] ap_bram_iarg_31_we0,
    input ap_bram_iarg_31_en0,
    input [S_AXIS_BRAM_31_ADDR_WIDTH-1:0] ap_bram_iarg_31_addr1,
    input [S_AXIS_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_din1,
    output [S_AXIS_BRAM_31_WIDTH-1:0] ap_bram_iarg_31_dout1,
    input ap_bram_iarg_31_clk1,
    input ap_bram_iarg_31_rst1,
    input [S_AXIS_BRAM_31_WIDTH/8-1:0] ap_bram_iarg_31_we1,
    input ap_bram_iarg_31_en1,
    //input AXI-Stream to BRAM interface 32
    input s_axis_bram_32_aclk,
    input s_axis_bram_32_aresetn,
    input s_axis_bram_32_tlast,
    input s_axis_bram_32_tvalid,
    input [S_AXIS_BRAM_32_DMWIDTH/8-1:0] s_axis_bram_32_tkeep,
    input [S_AXIS_BRAM_32_DMWIDTH/8-1:0] s_axis_bram_32_tstrb,
    input [S_AXIS_BRAM_32_DMWIDTH-1:0] s_axis_bram_32_tdata,
    output s_axis_bram_32_tready,
    input [S_AXIS_BRAM_32_ADDR_WIDTH-1:0] ap_bram_iarg_32_addr0,
    input [S_AXIS_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_din0,
    output [S_AXIS_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_dout0,
    input ap_bram_iarg_32_clk0,
    input ap_bram_iarg_32_rst0,
    input [S_AXIS_BRAM_32_WIDTH/8-1:0] ap_bram_iarg_32_we0,
    input ap_bram_iarg_32_en0,
    input [S_AXIS_BRAM_32_ADDR_WIDTH-1:0] ap_bram_iarg_32_addr1,
    input [S_AXIS_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_din1,
    output [S_AXIS_BRAM_32_WIDTH-1:0] ap_bram_iarg_32_dout1,
    input ap_bram_iarg_32_clk1,
    input ap_bram_iarg_32_rst1,
    input [S_AXIS_BRAM_32_WIDTH/8-1:0] ap_bram_iarg_32_we1,
    input ap_bram_iarg_32_en1,
    //input AXI-Stream to BRAM interface 33
    input s_axis_bram_33_aclk,
    input s_axis_bram_33_aresetn,
    input s_axis_bram_33_tlast,
    input s_axis_bram_33_tvalid,
    input [S_AXIS_BRAM_33_DMWIDTH/8-1:0] s_axis_bram_33_tkeep,
    input [S_AXIS_BRAM_33_DMWIDTH/8-1:0] s_axis_bram_33_tstrb,
    input [S_AXIS_BRAM_33_DMWIDTH-1:0] s_axis_bram_33_tdata,
    output s_axis_bram_33_tready,
    input [S_AXIS_BRAM_33_ADDR_WIDTH-1:0] ap_bram_iarg_33_addr0,
    input [S_AXIS_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_din0,
    output [S_AXIS_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_dout0,
    input ap_bram_iarg_33_clk0,
    input ap_bram_iarg_33_rst0,
    input [S_AXIS_BRAM_33_WIDTH/8-1:0] ap_bram_iarg_33_we0,
    input ap_bram_iarg_33_en0,
    input [S_AXIS_BRAM_33_ADDR_WIDTH-1:0] ap_bram_iarg_33_addr1,
    input [S_AXIS_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_din1,
    output [S_AXIS_BRAM_33_WIDTH-1:0] ap_bram_iarg_33_dout1,
    input ap_bram_iarg_33_clk1,
    input ap_bram_iarg_33_rst1,
    input [S_AXIS_BRAM_33_WIDTH/8-1:0] ap_bram_iarg_33_we1,
    input ap_bram_iarg_33_en1,
    //input AXI-Stream to BRAM interface 34
    input s_axis_bram_34_aclk,
    input s_axis_bram_34_aresetn,
    input s_axis_bram_34_tlast,
    input s_axis_bram_34_tvalid,
    input [S_AXIS_BRAM_34_DMWIDTH/8-1:0] s_axis_bram_34_tkeep,
    input [S_AXIS_BRAM_34_DMWIDTH/8-1:0] s_axis_bram_34_tstrb,
    input [S_AXIS_BRAM_34_DMWIDTH-1:0] s_axis_bram_34_tdata,
    output s_axis_bram_34_tready,
    input [S_AXIS_BRAM_34_ADDR_WIDTH-1:0] ap_bram_iarg_34_addr0,
    input [S_AXIS_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_din0,
    output [S_AXIS_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_dout0,
    input ap_bram_iarg_34_clk0,
    input ap_bram_iarg_34_rst0,
    input [S_AXIS_BRAM_34_WIDTH/8-1:0] ap_bram_iarg_34_we0,
    input ap_bram_iarg_34_en0,
    input [S_AXIS_BRAM_34_ADDR_WIDTH-1:0] ap_bram_iarg_34_addr1,
    input [S_AXIS_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_din1,
    output [S_AXIS_BRAM_34_WIDTH-1:0] ap_bram_iarg_34_dout1,
    input ap_bram_iarg_34_clk1,
    input ap_bram_iarg_34_rst1,
    input [S_AXIS_BRAM_34_WIDTH/8-1:0] ap_bram_iarg_34_we1,
    input ap_bram_iarg_34_en1,
    //input AXI-Stream to BRAM interface 35
    input s_axis_bram_35_aclk,
    input s_axis_bram_35_aresetn,
    input s_axis_bram_35_tlast,
    input s_axis_bram_35_tvalid,
    input [S_AXIS_BRAM_35_DMWIDTH/8-1:0] s_axis_bram_35_tkeep,
    input [S_AXIS_BRAM_35_DMWIDTH/8-1:0] s_axis_bram_35_tstrb,
    input [S_AXIS_BRAM_35_DMWIDTH-1:0] s_axis_bram_35_tdata,
    output s_axis_bram_35_tready,
    input [S_AXIS_BRAM_35_ADDR_WIDTH-1:0] ap_bram_iarg_35_addr0,
    input [S_AXIS_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_din0,
    output [S_AXIS_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_dout0,
    input ap_bram_iarg_35_clk0,
    input ap_bram_iarg_35_rst0,
    input [S_AXIS_BRAM_35_WIDTH/8-1:0] ap_bram_iarg_35_we0,
    input ap_bram_iarg_35_en0,
    input [S_AXIS_BRAM_35_ADDR_WIDTH-1:0] ap_bram_iarg_35_addr1,
    input [S_AXIS_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_din1,
    output [S_AXIS_BRAM_35_WIDTH-1:0] ap_bram_iarg_35_dout1,
    input ap_bram_iarg_35_clk1,
    input ap_bram_iarg_35_rst1,
    input [S_AXIS_BRAM_35_WIDTH/8-1:0] ap_bram_iarg_35_we1,
    input ap_bram_iarg_35_en1,
    //input AXI-Stream to BRAM interface 36
    input s_axis_bram_36_aclk,
    input s_axis_bram_36_aresetn,
    input s_axis_bram_36_tlast,
    input s_axis_bram_36_tvalid,
    input [S_AXIS_BRAM_36_DMWIDTH/8-1:0] s_axis_bram_36_tkeep,
    input [S_AXIS_BRAM_36_DMWIDTH/8-1:0] s_axis_bram_36_tstrb,
    input [S_AXIS_BRAM_36_DMWIDTH-1:0] s_axis_bram_36_tdata,
    output s_axis_bram_36_tready,
    input [S_AXIS_BRAM_36_ADDR_WIDTH-1:0] ap_bram_iarg_36_addr0,
    input [S_AXIS_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_din0,
    output [S_AXIS_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_dout0,
    input ap_bram_iarg_36_clk0,
    input ap_bram_iarg_36_rst0,
    input [S_AXIS_BRAM_36_WIDTH/8-1:0] ap_bram_iarg_36_we0,
    input ap_bram_iarg_36_en0,
    input [S_AXIS_BRAM_36_ADDR_WIDTH-1:0] ap_bram_iarg_36_addr1,
    input [S_AXIS_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_din1,
    output [S_AXIS_BRAM_36_WIDTH-1:0] ap_bram_iarg_36_dout1,
    input ap_bram_iarg_36_clk1,
    input ap_bram_iarg_36_rst1,
    input [S_AXIS_BRAM_36_WIDTH/8-1:0] ap_bram_iarg_36_we1,
    input ap_bram_iarg_36_en1,
    //input AXI-Stream to BRAM interface 37
    input s_axis_bram_37_aclk,
    input s_axis_bram_37_aresetn,
    input s_axis_bram_37_tlast,
    input s_axis_bram_37_tvalid,
    input [S_AXIS_BRAM_37_DMWIDTH/8-1:0] s_axis_bram_37_tkeep,
    input [S_AXIS_BRAM_37_DMWIDTH/8-1:0] s_axis_bram_37_tstrb,
    input [S_AXIS_BRAM_37_DMWIDTH-1:0] s_axis_bram_37_tdata,
    output s_axis_bram_37_tready,
    input [S_AXIS_BRAM_37_ADDR_WIDTH-1:0] ap_bram_iarg_37_addr0,
    input [S_AXIS_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_din0,
    output [S_AXIS_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_dout0,
    input ap_bram_iarg_37_clk0,
    input ap_bram_iarg_37_rst0,
    input [S_AXIS_BRAM_37_WIDTH/8-1:0] ap_bram_iarg_37_we0,
    input ap_bram_iarg_37_en0,
    input [S_AXIS_BRAM_37_ADDR_WIDTH-1:0] ap_bram_iarg_37_addr1,
    input [S_AXIS_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_din1,
    output [S_AXIS_BRAM_37_WIDTH-1:0] ap_bram_iarg_37_dout1,
    input ap_bram_iarg_37_clk1,
    input ap_bram_iarg_37_rst1,
    input [S_AXIS_BRAM_37_WIDTH/8-1:0] ap_bram_iarg_37_we1,
    input ap_bram_iarg_37_en1,
    //input AXI-Stream to BRAM interface 38
    input s_axis_bram_38_aclk,
    input s_axis_bram_38_aresetn,
    input s_axis_bram_38_tlast,
    input s_axis_bram_38_tvalid,
    input [S_AXIS_BRAM_38_DMWIDTH/8-1:0] s_axis_bram_38_tkeep,
    input [S_AXIS_BRAM_38_DMWIDTH/8-1:0] s_axis_bram_38_tstrb,
    input [S_AXIS_BRAM_38_DMWIDTH-1:0] s_axis_bram_38_tdata,
    output s_axis_bram_38_tready,
    input [S_AXIS_BRAM_38_ADDR_WIDTH-1:0] ap_bram_iarg_38_addr0,
    input [S_AXIS_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_din0,
    output [S_AXIS_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_dout0,
    input ap_bram_iarg_38_clk0,
    input ap_bram_iarg_38_rst0,
    input [S_AXIS_BRAM_38_WIDTH/8-1:0] ap_bram_iarg_38_we0,
    input ap_bram_iarg_38_en0,
    input [S_AXIS_BRAM_38_ADDR_WIDTH-1:0] ap_bram_iarg_38_addr1,
    input [S_AXIS_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_din1,
    output [S_AXIS_BRAM_38_WIDTH-1:0] ap_bram_iarg_38_dout1,
    input ap_bram_iarg_38_clk1,
    input ap_bram_iarg_38_rst1,
    input [S_AXIS_BRAM_38_WIDTH/8-1:0] ap_bram_iarg_38_we1,
    input ap_bram_iarg_38_en1,
    //input AXI-Stream to BRAM interface 39
    input s_axis_bram_39_aclk,
    input s_axis_bram_39_aresetn,
    input s_axis_bram_39_tlast,
    input s_axis_bram_39_tvalid,
    input [S_AXIS_BRAM_39_DMWIDTH/8-1:0] s_axis_bram_39_tkeep,
    input [S_AXIS_BRAM_39_DMWIDTH/8-1:0] s_axis_bram_39_tstrb,
    input [S_AXIS_BRAM_39_DMWIDTH-1:0] s_axis_bram_39_tdata,
    output s_axis_bram_39_tready,
    input [S_AXIS_BRAM_39_ADDR_WIDTH-1:0] ap_bram_iarg_39_addr0,
    input [S_AXIS_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_din0,
    output [S_AXIS_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_dout0,
    input ap_bram_iarg_39_clk0,
    input ap_bram_iarg_39_rst0,
    input [S_AXIS_BRAM_39_WIDTH/8-1:0] ap_bram_iarg_39_we0,
    input ap_bram_iarg_39_en0,
    input [S_AXIS_BRAM_39_ADDR_WIDTH-1:0] ap_bram_iarg_39_addr1,
    input [S_AXIS_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_din1,
    output [S_AXIS_BRAM_39_WIDTH-1:0] ap_bram_iarg_39_dout1,
    input ap_bram_iarg_39_clk1,
    input ap_bram_iarg_39_rst1,
    input [S_AXIS_BRAM_39_WIDTH/8-1:0] ap_bram_iarg_39_we1,
    input ap_bram_iarg_39_en1,
    //input AXI-Stream to BRAM interface 40
    input s_axis_bram_40_aclk,
    input s_axis_bram_40_aresetn,
    input s_axis_bram_40_tlast,
    input s_axis_bram_40_tvalid,
    input [S_AXIS_BRAM_40_DMWIDTH/8-1:0] s_axis_bram_40_tkeep,
    input [S_AXIS_BRAM_40_DMWIDTH/8-1:0] s_axis_bram_40_tstrb,
    input [S_AXIS_BRAM_40_DMWIDTH-1:0] s_axis_bram_40_tdata,
    output s_axis_bram_40_tready,
    input [S_AXIS_BRAM_40_ADDR_WIDTH-1:0] ap_bram_iarg_40_addr0,
    input [S_AXIS_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_din0,
    output [S_AXIS_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_dout0,
    input ap_bram_iarg_40_clk0,
    input ap_bram_iarg_40_rst0,
    input [S_AXIS_BRAM_40_WIDTH/8-1:0] ap_bram_iarg_40_we0,
    input ap_bram_iarg_40_en0,
    input [S_AXIS_BRAM_40_ADDR_WIDTH-1:0] ap_bram_iarg_40_addr1,
    input [S_AXIS_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_din1,
    output [S_AXIS_BRAM_40_WIDTH-1:0] ap_bram_iarg_40_dout1,
    input ap_bram_iarg_40_clk1,
    input ap_bram_iarg_40_rst1,
    input [S_AXIS_BRAM_40_WIDTH/8-1:0] ap_bram_iarg_40_we1,
    input ap_bram_iarg_40_en1,
    //input AXI-Stream to BRAM interface 41
    input s_axis_bram_41_aclk,
    input s_axis_bram_41_aresetn,
    input s_axis_bram_41_tlast,
    input s_axis_bram_41_tvalid,
    input [S_AXIS_BRAM_41_DMWIDTH/8-1:0] s_axis_bram_41_tkeep,
    input [S_AXIS_BRAM_41_DMWIDTH/8-1:0] s_axis_bram_41_tstrb,
    input [S_AXIS_BRAM_41_DMWIDTH-1:0] s_axis_bram_41_tdata,
    output s_axis_bram_41_tready,
    input [S_AXIS_BRAM_41_ADDR_WIDTH-1:0] ap_bram_iarg_41_addr0,
    input [S_AXIS_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_din0,
    output [S_AXIS_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_dout0,
    input ap_bram_iarg_41_clk0,
    input ap_bram_iarg_41_rst0,
    input [S_AXIS_BRAM_41_WIDTH/8-1:0] ap_bram_iarg_41_we0,
    input ap_bram_iarg_41_en0,
    input [S_AXIS_BRAM_41_ADDR_WIDTH-1:0] ap_bram_iarg_41_addr1,
    input [S_AXIS_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_din1,
    output [S_AXIS_BRAM_41_WIDTH-1:0] ap_bram_iarg_41_dout1,
    input ap_bram_iarg_41_clk1,
    input ap_bram_iarg_41_rst1,
    input [S_AXIS_BRAM_41_WIDTH/8-1:0] ap_bram_iarg_41_we1,
    input ap_bram_iarg_41_en1,
    //input AXI-Stream to BRAM interface 42
    input s_axis_bram_42_aclk,
    input s_axis_bram_42_aresetn,
    input s_axis_bram_42_tlast,
    input s_axis_bram_42_tvalid,
    input [S_AXIS_BRAM_42_DMWIDTH/8-1:0] s_axis_bram_42_tkeep,
    input [S_AXIS_BRAM_42_DMWIDTH/8-1:0] s_axis_bram_42_tstrb,
    input [S_AXIS_BRAM_42_DMWIDTH-1:0] s_axis_bram_42_tdata,
    output s_axis_bram_42_tready,
    input [S_AXIS_BRAM_42_ADDR_WIDTH-1:0] ap_bram_iarg_42_addr0,
    input [S_AXIS_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_din0,
    output [S_AXIS_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_dout0,
    input ap_bram_iarg_42_clk0,
    input ap_bram_iarg_42_rst0,
    input [S_AXIS_BRAM_42_WIDTH/8-1:0] ap_bram_iarg_42_we0,
    input ap_bram_iarg_42_en0,
    input [S_AXIS_BRAM_42_ADDR_WIDTH-1:0] ap_bram_iarg_42_addr1,
    input [S_AXIS_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_din1,
    output [S_AXIS_BRAM_42_WIDTH-1:0] ap_bram_iarg_42_dout1,
    input ap_bram_iarg_42_clk1,
    input ap_bram_iarg_42_rst1,
    input [S_AXIS_BRAM_42_WIDTH/8-1:0] ap_bram_iarg_42_we1,
    input ap_bram_iarg_42_en1,
    //input AXI-Stream to BRAM interface 43
    input s_axis_bram_43_aclk,
    input s_axis_bram_43_aresetn,
    input s_axis_bram_43_tlast,
    input s_axis_bram_43_tvalid,
    input [S_AXIS_BRAM_43_DMWIDTH/8-1:0] s_axis_bram_43_tkeep,
    input [S_AXIS_BRAM_43_DMWIDTH/8-1:0] s_axis_bram_43_tstrb,
    input [S_AXIS_BRAM_43_DMWIDTH-1:0] s_axis_bram_43_tdata,
    output s_axis_bram_43_tready,
    input [S_AXIS_BRAM_43_ADDR_WIDTH-1:0] ap_bram_iarg_43_addr0,
    input [S_AXIS_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_din0,
    output [S_AXIS_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_dout0,
    input ap_bram_iarg_43_clk0,
    input ap_bram_iarg_43_rst0,
    input [S_AXIS_BRAM_43_WIDTH/8-1:0] ap_bram_iarg_43_we0,
    input ap_bram_iarg_43_en0,
    input [S_AXIS_BRAM_43_ADDR_WIDTH-1:0] ap_bram_iarg_43_addr1,
    input [S_AXIS_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_din1,
    output [S_AXIS_BRAM_43_WIDTH-1:0] ap_bram_iarg_43_dout1,
    input ap_bram_iarg_43_clk1,
    input ap_bram_iarg_43_rst1,
    input [S_AXIS_BRAM_43_WIDTH/8-1:0] ap_bram_iarg_43_we1,
    input ap_bram_iarg_43_en1,
    //input AXI-Stream to BRAM interface 44
    input s_axis_bram_44_aclk,
    input s_axis_bram_44_aresetn,
    input s_axis_bram_44_tlast,
    input s_axis_bram_44_tvalid,
    input [S_AXIS_BRAM_44_DMWIDTH/8-1:0] s_axis_bram_44_tkeep,
    input [S_AXIS_BRAM_44_DMWIDTH/8-1:0] s_axis_bram_44_tstrb,
    input [S_AXIS_BRAM_44_DMWIDTH-1:0] s_axis_bram_44_tdata,
    output s_axis_bram_44_tready,
    input [S_AXIS_BRAM_44_ADDR_WIDTH-1:0] ap_bram_iarg_44_addr0,
    input [S_AXIS_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_din0,
    output [S_AXIS_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_dout0,
    input ap_bram_iarg_44_clk0,
    input ap_bram_iarg_44_rst0,
    input [S_AXIS_BRAM_44_WIDTH/8-1:0] ap_bram_iarg_44_we0,
    input ap_bram_iarg_44_en0,
    input [S_AXIS_BRAM_44_ADDR_WIDTH-1:0] ap_bram_iarg_44_addr1,
    input [S_AXIS_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_din1,
    output [S_AXIS_BRAM_44_WIDTH-1:0] ap_bram_iarg_44_dout1,
    input ap_bram_iarg_44_clk1,
    input ap_bram_iarg_44_rst1,
    input [S_AXIS_BRAM_44_WIDTH/8-1:0] ap_bram_iarg_44_we1,
    input ap_bram_iarg_44_en1,
    //input AXI-Stream to BRAM interface 45
    input s_axis_bram_45_aclk,
    input s_axis_bram_45_aresetn,
    input s_axis_bram_45_tlast,
    input s_axis_bram_45_tvalid,
    input [S_AXIS_BRAM_45_DMWIDTH/8-1:0] s_axis_bram_45_tkeep,
    input [S_AXIS_BRAM_45_DMWIDTH/8-1:0] s_axis_bram_45_tstrb,
    input [S_AXIS_BRAM_45_DMWIDTH-1:0] s_axis_bram_45_tdata,
    output s_axis_bram_45_tready,
    input [S_AXIS_BRAM_45_ADDR_WIDTH-1:0] ap_bram_iarg_45_addr0,
    input [S_AXIS_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_din0,
    output [S_AXIS_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_dout0,
    input ap_bram_iarg_45_clk0,
    input ap_bram_iarg_45_rst0,
    input [S_AXIS_BRAM_45_WIDTH/8-1:0] ap_bram_iarg_45_we0,
    input ap_bram_iarg_45_en0,
    input [S_AXIS_BRAM_45_ADDR_WIDTH-1:0] ap_bram_iarg_45_addr1,
    input [S_AXIS_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_din1,
    output [S_AXIS_BRAM_45_WIDTH-1:0] ap_bram_iarg_45_dout1,
    input ap_bram_iarg_45_clk1,
    input ap_bram_iarg_45_rst1,
    input [S_AXIS_BRAM_45_WIDTH/8-1:0] ap_bram_iarg_45_we1,
    input ap_bram_iarg_45_en1,
    //input AXI-Stream to BRAM interface 46
    input s_axis_bram_46_aclk,
    input s_axis_bram_46_aresetn,
    input s_axis_bram_46_tlast,
    input s_axis_bram_46_tvalid,
    input [S_AXIS_BRAM_46_DMWIDTH/8-1:0] s_axis_bram_46_tkeep,
    input [S_AXIS_BRAM_46_DMWIDTH/8-1:0] s_axis_bram_46_tstrb,
    input [S_AXIS_BRAM_46_DMWIDTH-1:0] s_axis_bram_46_tdata,
    output s_axis_bram_46_tready,
    input [S_AXIS_BRAM_46_ADDR_WIDTH-1:0] ap_bram_iarg_46_addr0,
    input [S_AXIS_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_din0,
    output [S_AXIS_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_dout0,
    input ap_bram_iarg_46_clk0,
    input ap_bram_iarg_46_rst0,
    input [S_AXIS_BRAM_46_WIDTH/8-1:0] ap_bram_iarg_46_we0,
    input ap_bram_iarg_46_en0,
    input [S_AXIS_BRAM_46_ADDR_WIDTH-1:0] ap_bram_iarg_46_addr1,
    input [S_AXIS_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_din1,
    output [S_AXIS_BRAM_46_WIDTH-1:0] ap_bram_iarg_46_dout1,
    input ap_bram_iarg_46_clk1,
    input ap_bram_iarg_46_rst1,
    input [S_AXIS_BRAM_46_WIDTH/8-1:0] ap_bram_iarg_46_we1,
    input ap_bram_iarg_46_en1,
    //input AXI-Stream to BRAM interface 47
    input s_axis_bram_47_aclk,
    input s_axis_bram_47_aresetn,
    input s_axis_bram_47_tlast,
    input s_axis_bram_47_tvalid,
    input [S_AXIS_BRAM_47_DMWIDTH/8-1:0] s_axis_bram_47_tkeep,
    input [S_AXIS_BRAM_47_DMWIDTH/8-1:0] s_axis_bram_47_tstrb,
    input [S_AXIS_BRAM_47_DMWIDTH-1:0] s_axis_bram_47_tdata,
    output s_axis_bram_47_tready,
    input [S_AXIS_BRAM_47_ADDR_WIDTH-1:0] ap_bram_iarg_47_addr0,
    input [S_AXIS_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_din0,
    output [S_AXIS_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_dout0,
    input ap_bram_iarg_47_clk0,
    input ap_bram_iarg_47_rst0,
    input [S_AXIS_BRAM_47_WIDTH/8-1:0] ap_bram_iarg_47_we0,
    input ap_bram_iarg_47_en0,
    input [S_AXIS_BRAM_47_ADDR_WIDTH-1:0] ap_bram_iarg_47_addr1,
    input [S_AXIS_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_din1,
    output [S_AXIS_BRAM_47_WIDTH-1:0] ap_bram_iarg_47_dout1,
    input ap_bram_iarg_47_clk1,
    input ap_bram_iarg_47_rst1,
    input [S_AXIS_BRAM_47_WIDTH/8-1:0] ap_bram_iarg_47_we1,
    input ap_bram_iarg_47_en1,
    //input AXI-Stream to BRAM interface 48
    input s_axis_bram_48_aclk,
    input s_axis_bram_48_aresetn,
    input s_axis_bram_48_tlast,
    input s_axis_bram_48_tvalid,
    input [S_AXIS_BRAM_48_DMWIDTH/8-1:0] s_axis_bram_48_tkeep,
    input [S_AXIS_BRAM_48_DMWIDTH/8-1:0] s_axis_bram_48_tstrb,
    input [S_AXIS_BRAM_48_DMWIDTH-1:0] s_axis_bram_48_tdata,
    output s_axis_bram_48_tready,
    input [S_AXIS_BRAM_48_ADDR_WIDTH-1:0] ap_bram_iarg_48_addr0,
    input [S_AXIS_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_din0,
    output [S_AXIS_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_dout0,
    input ap_bram_iarg_48_clk0,
    input ap_bram_iarg_48_rst0,
    input [S_AXIS_BRAM_48_WIDTH/8-1:0] ap_bram_iarg_48_we0,
    input ap_bram_iarg_48_en0,
    input [S_AXIS_BRAM_48_ADDR_WIDTH-1:0] ap_bram_iarg_48_addr1,
    input [S_AXIS_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_din1,
    output [S_AXIS_BRAM_48_WIDTH-1:0] ap_bram_iarg_48_dout1,
    input ap_bram_iarg_48_clk1,
    input ap_bram_iarg_48_rst1,
    input [S_AXIS_BRAM_48_WIDTH/8-1:0] ap_bram_iarg_48_we1,
    input ap_bram_iarg_48_en1,
    //input AXI-Stream to BRAM interface 49
    input s_axis_bram_49_aclk,
    input s_axis_bram_49_aresetn,
    input s_axis_bram_49_tlast,
    input s_axis_bram_49_tvalid,
    input [S_AXIS_BRAM_49_DMWIDTH/8-1:0] s_axis_bram_49_tkeep,
    input [S_AXIS_BRAM_49_DMWIDTH/8-1:0] s_axis_bram_49_tstrb,
    input [S_AXIS_BRAM_49_DMWIDTH-1:0] s_axis_bram_49_tdata,
    output s_axis_bram_49_tready,
    input [S_AXIS_BRAM_49_ADDR_WIDTH-1:0] ap_bram_iarg_49_addr0,
    input [S_AXIS_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_din0,
    output [S_AXIS_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_dout0,
    input ap_bram_iarg_49_clk0,
    input ap_bram_iarg_49_rst0,
    input [S_AXIS_BRAM_49_WIDTH/8-1:0] ap_bram_iarg_49_we0,
    input ap_bram_iarg_49_en0,
    input [S_AXIS_BRAM_49_ADDR_WIDTH-1:0] ap_bram_iarg_49_addr1,
    input [S_AXIS_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_din1,
    output [S_AXIS_BRAM_49_WIDTH-1:0] ap_bram_iarg_49_dout1,
    input ap_bram_iarg_49_clk1,
    input ap_bram_iarg_49_rst1,
    input [S_AXIS_BRAM_49_WIDTH/8-1:0] ap_bram_iarg_49_we1,
    input ap_bram_iarg_49_en1,
    //input AXI-Stream to BRAM interface 50
    input s_axis_bram_50_aclk,
    input s_axis_bram_50_aresetn,
    input s_axis_bram_50_tlast,
    input s_axis_bram_50_tvalid,
    input [S_AXIS_BRAM_50_DMWIDTH/8-1:0] s_axis_bram_50_tkeep,
    input [S_AXIS_BRAM_50_DMWIDTH/8-1:0] s_axis_bram_50_tstrb,
    input [S_AXIS_BRAM_50_DMWIDTH-1:0] s_axis_bram_50_tdata,
    output s_axis_bram_50_tready,
    input [S_AXIS_BRAM_50_ADDR_WIDTH-1:0] ap_bram_iarg_50_addr0,
    input [S_AXIS_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_din0,
    output [S_AXIS_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_dout0,
    input ap_bram_iarg_50_clk0,
    input ap_bram_iarg_50_rst0,
    input [S_AXIS_BRAM_50_WIDTH/8-1:0] ap_bram_iarg_50_we0,
    input ap_bram_iarg_50_en0,
    input [S_AXIS_BRAM_50_ADDR_WIDTH-1:0] ap_bram_iarg_50_addr1,
    input [S_AXIS_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_din1,
    output [S_AXIS_BRAM_50_WIDTH-1:0] ap_bram_iarg_50_dout1,
    input ap_bram_iarg_50_clk1,
    input ap_bram_iarg_50_rst1,
    input [S_AXIS_BRAM_50_WIDTH/8-1:0] ap_bram_iarg_50_we1,
    input ap_bram_iarg_50_en1,
    //input AXI-Stream to BRAM interface 51
    input s_axis_bram_51_aclk,
    input s_axis_bram_51_aresetn,
    input s_axis_bram_51_tlast,
    input s_axis_bram_51_tvalid,
    input [S_AXIS_BRAM_51_DMWIDTH/8-1:0] s_axis_bram_51_tkeep,
    input [S_AXIS_BRAM_51_DMWIDTH/8-1:0] s_axis_bram_51_tstrb,
    input [S_AXIS_BRAM_51_DMWIDTH-1:0] s_axis_bram_51_tdata,
    output s_axis_bram_51_tready,
    input [S_AXIS_BRAM_51_ADDR_WIDTH-1:0] ap_bram_iarg_51_addr0,
    input [S_AXIS_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_din0,
    output [S_AXIS_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_dout0,
    input ap_bram_iarg_51_clk0,
    input ap_bram_iarg_51_rst0,
    input [S_AXIS_BRAM_51_WIDTH/8-1:0] ap_bram_iarg_51_we0,
    input ap_bram_iarg_51_en0,
    input [S_AXIS_BRAM_51_ADDR_WIDTH-1:0] ap_bram_iarg_51_addr1,
    input [S_AXIS_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_din1,
    output [S_AXIS_BRAM_51_WIDTH-1:0] ap_bram_iarg_51_dout1,
    input ap_bram_iarg_51_clk1,
    input ap_bram_iarg_51_rst1,
    input [S_AXIS_BRAM_51_WIDTH/8-1:0] ap_bram_iarg_51_we1,
    input ap_bram_iarg_51_en1,
    //input AXI-Stream to BRAM interface 52
    input s_axis_bram_52_aclk,
    input s_axis_bram_52_aresetn,
    input s_axis_bram_52_tlast,
    input s_axis_bram_52_tvalid,
    input [S_AXIS_BRAM_52_DMWIDTH/8-1:0] s_axis_bram_52_tkeep,
    input [S_AXIS_BRAM_52_DMWIDTH/8-1:0] s_axis_bram_52_tstrb,
    input [S_AXIS_BRAM_52_DMWIDTH-1:0] s_axis_bram_52_tdata,
    output s_axis_bram_52_tready,
    input [S_AXIS_BRAM_52_ADDR_WIDTH-1:0] ap_bram_iarg_52_addr0,
    input [S_AXIS_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_din0,
    output [S_AXIS_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_dout0,
    input ap_bram_iarg_52_clk0,
    input ap_bram_iarg_52_rst0,
    input [S_AXIS_BRAM_52_WIDTH/8-1:0] ap_bram_iarg_52_we0,
    input ap_bram_iarg_52_en0,
    input [S_AXIS_BRAM_52_ADDR_WIDTH-1:0] ap_bram_iarg_52_addr1,
    input [S_AXIS_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_din1,
    output [S_AXIS_BRAM_52_WIDTH-1:0] ap_bram_iarg_52_dout1,
    input ap_bram_iarg_52_clk1,
    input ap_bram_iarg_52_rst1,
    input [S_AXIS_BRAM_52_WIDTH/8-1:0] ap_bram_iarg_52_we1,
    input ap_bram_iarg_52_en1,
    //input AXI-Stream to BRAM interface 53
    input s_axis_bram_53_aclk,
    input s_axis_bram_53_aresetn,
    input s_axis_bram_53_tlast,
    input s_axis_bram_53_tvalid,
    input [S_AXIS_BRAM_53_DMWIDTH/8-1:0] s_axis_bram_53_tkeep,
    input [S_AXIS_BRAM_53_DMWIDTH/8-1:0] s_axis_bram_53_tstrb,
    input [S_AXIS_BRAM_53_DMWIDTH-1:0] s_axis_bram_53_tdata,
    output s_axis_bram_53_tready,
    input [S_AXIS_BRAM_53_ADDR_WIDTH-1:0] ap_bram_iarg_53_addr0,
    input [S_AXIS_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_din0,
    output [S_AXIS_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_dout0,
    input ap_bram_iarg_53_clk0,
    input ap_bram_iarg_53_rst0,
    input [S_AXIS_BRAM_53_WIDTH/8-1:0] ap_bram_iarg_53_we0,
    input ap_bram_iarg_53_en0,
    input [S_AXIS_BRAM_53_ADDR_WIDTH-1:0] ap_bram_iarg_53_addr1,
    input [S_AXIS_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_din1,
    output [S_AXIS_BRAM_53_WIDTH-1:0] ap_bram_iarg_53_dout1,
    input ap_bram_iarg_53_clk1,
    input ap_bram_iarg_53_rst1,
    input [S_AXIS_BRAM_53_WIDTH/8-1:0] ap_bram_iarg_53_we1,
    input ap_bram_iarg_53_en1,
    //input AXI-Stream to BRAM interface 54
    input s_axis_bram_54_aclk,
    input s_axis_bram_54_aresetn,
    input s_axis_bram_54_tlast,
    input s_axis_bram_54_tvalid,
    input [S_AXIS_BRAM_54_DMWIDTH/8-1:0] s_axis_bram_54_tkeep,
    input [S_AXIS_BRAM_54_DMWIDTH/8-1:0] s_axis_bram_54_tstrb,
    input [S_AXIS_BRAM_54_DMWIDTH-1:0] s_axis_bram_54_tdata,
    output s_axis_bram_54_tready,
    input [S_AXIS_BRAM_54_ADDR_WIDTH-1:0] ap_bram_iarg_54_addr0,
    input [S_AXIS_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_din0,
    output [S_AXIS_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_dout0,
    input ap_bram_iarg_54_clk0,
    input ap_bram_iarg_54_rst0,
    input [S_AXIS_BRAM_54_WIDTH/8-1:0] ap_bram_iarg_54_we0,
    input ap_bram_iarg_54_en0,
    input [S_AXIS_BRAM_54_ADDR_WIDTH-1:0] ap_bram_iarg_54_addr1,
    input [S_AXIS_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_din1,
    output [S_AXIS_BRAM_54_WIDTH-1:0] ap_bram_iarg_54_dout1,
    input ap_bram_iarg_54_clk1,
    input ap_bram_iarg_54_rst1,
    input [S_AXIS_BRAM_54_WIDTH/8-1:0] ap_bram_iarg_54_we1,
    input ap_bram_iarg_54_en1,
    //input AXI-Stream to BRAM interface 55
    input s_axis_bram_55_aclk,
    input s_axis_bram_55_aresetn,
    input s_axis_bram_55_tlast,
    input s_axis_bram_55_tvalid,
    input [S_AXIS_BRAM_55_DMWIDTH/8-1:0] s_axis_bram_55_tkeep,
    input [S_AXIS_BRAM_55_DMWIDTH/8-1:0] s_axis_bram_55_tstrb,
    input [S_AXIS_BRAM_55_DMWIDTH-1:0] s_axis_bram_55_tdata,
    output s_axis_bram_55_tready,
    input [S_AXIS_BRAM_55_ADDR_WIDTH-1:0] ap_bram_iarg_55_addr0,
    input [S_AXIS_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_din0,
    output [S_AXIS_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_dout0,
    input ap_bram_iarg_55_clk0,
    input ap_bram_iarg_55_rst0,
    input [S_AXIS_BRAM_55_WIDTH/8-1:0] ap_bram_iarg_55_we0,
    input ap_bram_iarg_55_en0,
    input [S_AXIS_BRAM_55_ADDR_WIDTH-1:0] ap_bram_iarg_55_addr1,
    input [S_AXIS_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_din1,
    output [S_AXIS_BRAM_55_WIDTH-1:0] ap_bram_iarg_55_dout1,
    input ap_bram_iarg_55_clk1,
    input ap_bram_iarg_55_rst1,
    input [S_AXIS_BRAM_55_WIDTH/8-1:0] ap_bram_iarg_55_we1,
    input ap_bram_iarg_55_en1,
    //input AXI-Stream to BRAM interface 56
    input s_axis_bram_56_aclk,
    input s_axis_bram_56_aresetn,
    input s_axis_bram_56_tlast,
    input s_axis_bram_56_tvalid,
    input [S_AXIS_BRAM_56_DMWIDTH/8-1:0] s_axis_bram_56_tkeep,
    input [S_AXIS_BRAM_56_DMWIDTH/8-1:0] s_axis_bram_56_tstrb,
    input [S_AXIS_BRAM_56_DMWIDTH-1:0] s_axis_bram_56_tdata,
    output s_axis_bram_56_tready,
    input [S_AXIS_BRAM_56_ADDR_WIDTH-1:0] ap_bram_iarg_56_addr0,
    input [S_AXIS_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_din0,
    output [S_AXIS_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_dout0,
    input ap_bram_iarg_56_clk0,
    input ap_bram_iarg_56_rst0,
    input [S_AXIS_BRAM_56_WIDTH/8-1:0] ap_bram_iarg_56_we0,
    input ap_bram_iarg_56_en0,
    input [S_AXIS_BRAM_56_ADDR_WIDTH-1:0] ap_bram_iarg_56_addr1,
    input [S_AXIS_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_din1,
    output [S_AXIS_BRAM_56_WIDTH-1:0] ap_bram_iarg_56_dout1,
    input ap_bram_iarg_56_clk1,
    input ap_bram_iarg_56_rst1,
    input [S_AXIS_BRAM_56_WIDTH/8-1:0] ap_bram_iarg_56_we1,
    input ap_bram_iarg_56_en1,
    //input AXI-Stream to BRAM interface 57
    input s_axis_bram_57_aclk,
    input s_axis_bram_57_aresetn,
    input s_axis_bram_57_tlast,
    input s_axis_bram_57_tvalid,
    input [S_AXIS_BRAM_57_DMWIDTH/8-1:0] s_axis_bram_57_tkeep,
    input [S_AXIS_BRAM_57_DMWIDTH/8-1:0] s_axis_bram_57_tstrb,
    input [S_AXIS_BRAM_57_DMWIDTH-1:0] s_axis_bram_57_tdata,
    output s_axis_bram_57_tready,
    input [S_AXIS_BRAM_57_ADDR_WIDTH-1:0] ap_bram_iarg_57_addr0,
    input [S_AXIS_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_din0,
    output [S_AXIS_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_dout0,
    input ap_bram_iarg_57_clk0,
    input ap_bram_iarg_57_rst0,
    input [S_AXIS_BRAM_57_WIDTH/8-1:0] ap_bram_iarg_57_we0,
    input ap_bram_iarg_57_en0,
    input [S_AXIS_BRAM_57_ADDR_WIDTH-1:0] ap_bram_iarg_57_addr1,
    input [S_AXIS_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_din1,
    output [S_AXIS_BRAM_57_WIDTH-1:0] ap_bram_iarg_57_dout1,
    input ap_bram_iarg_57_clk1,
    input ap_bram_iarg_57_rst1,
    input [S_AXIS_BRAM_57_WIDTH/8-1:0] ap_bram_iarg_57_we1,
    input ap_bram_iarg_57_en1,
    //input AXI-Stream to BRAM interface 58
    input s_axis_bram_58_aclk,
    input s_axis_bram_58_aresetn,
    input s_axis_bram_58_tlast,
    input s_axis_bram_58_tvalid,
    input [S_AXIS_BRAM_58_DMWIDTH/8-1:0] s_axis_bram_58_tkeep,
    input [S_AXIS_BRAM_58_DMWIDTH/8-1:0] s_axis_bram_58_tstrb,
    input [S_AXIS_BRAM_58_DMWIDTH-1:0] s_axis_bram_58_tdata,
    output s_axis_bram_58_tready,
    input [S_AXIS_BRAM_58_ADDR_WIDTH-1:0] ap_bram_iarg_58_addr0,
    input [S_AXIS_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_din0,
    output [S_AXIS_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_dout0,
    input ap_bram_iarg_58_clk0,
    input ap_bram_iarg_58_rst0,
    input [S_AXIS_BRAM_58_WIDTH/8-1:0] ap_bram_iarg_58_we0,
    input ap_bram_iarg_58_en0,
    input [S_AXIS_BRAM_58_ADDR_WIDTH-1:0] ap_bram_iarg_58_addr1,
    input [S_AXIS_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_din1,
    output [S_AXIS_BRAM_58_WIDTH-1:0] ap_bram_iarg_58_dout1,
    input ap_bram_iarg_58_clk1,
    input ap_bram_iarg_58_rst1,
    input [S_AXIS_BRAM_58_WIDTH/8-1:0] ap_bram_iarg_58_we1,
    input ap_bram_iarg_58_en1,
    //input AXI-Stream to BRAM interface 59
    input s_axis_bram_59_aclk,
    input s_axis_bram_59_aresetn,
    input s_axis_bram_59_tlast,
    input s_axis_bram_59_tvalid,
    input [S_AXIS_BRAM_59_DMWIDTH/8-1:0] s_axis_bram_59_tkeep,
    input [S_AXIS_BRAM_59_DMWIDTH/8-1:0] s_axis_bram_59_tstrb,
    input [S_AXIS_BRAM_59_DMWIDTH-1:0] s_axis_bram_59_tdata,
    output s_axis_bram_59_tready,
    input [S_AXIS_BRAM_59_ADDR_WIDTH-1:0] ap_bram_iarg_59_addr0,
    input [S_AXIS_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_din0,
    output [S_AXIS_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_dout0,
    input ap_bram_iarg_59_clk0,
    input ap_bram_iarg_59_rst0,
    input [S_AXIS_BRAM_59_WIDTH/8-1:0] ap_bram_iarg_59_we0,
    input ap_bram_iarg_59_en0,
    input [S_AXIS_BRAM_59_ADDR_WIDTH-1:0] ap_bram_iarg_59_addr1,
    input [S_AXIS_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_din1,
    output [S_AXIS_BRAM_59_WIDTH-1:0] ap_bram_iarg_59_dout1,
    input ap_bram_iarg_59_clk1,
    input ap_bram_iarg_59_rst1,
    input [S_AXIS_BRAM_59_WIDTH/8-1:0] ap_bram_iarg_59_we1,
    input ap_bram_iarg_59_en1,
    //input AXI-Stream to BRAM interface 60
    input s_axis_bram_60_aclk,
    input s_axis_bram_60_aresetn,
    input s_axis_bram_60_tlast,
    input s_axis_bram_60_tvalid,
    input [S_AXIS_BRAM_60_DMWIDTH/8-1:0] s_axis_bram_60_tkeep,
    input [S_AXIS_BRAM_60_DMWIDTH/8-1:0] s_axis_bram_60_tstrb,
    input [S_AXIS_BRAM_60_DMWIDTH-1:0] s_axis_bram_60_tdata,
    output s_axis_bram_60_tready,
    input [S_AXIS_BRAM_60_ADDR_WIDTH-1:0] ap_bram_iarg_60_addr0,
    input [S_AXIS_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_din0,
    output [S_AXIS_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_dout0,
    input ap_bram_iarg_60_clk0,
    input ap_bram_iarg_60_rst0,
    input [S_AXIS_BRAM_60_WIDTH/8-1:0] ap_bram_iarg_60_we0,
    input ap_bram_iarg_60_en0,
    input [S_AXIS_BRAM_60_ADDR_WIDTH-1:0] ap_bram_iarg_60_addr1,
    input [S_AXIS_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_din1,
    output [S_AXIS_BRAM_60_WIDTH-1:0] ap_bram_iarg_60_dout1,
    input ap_bram_iarg_60_clk1,
    input ap_bram_iarg_60_rst1,
    input [S_AXIS_BRAM_60_WIDTH/8-1:0] ap_bram_iarg_60_we1,
    input ap_bram_iarg_60_en1,
    //input AXI-Stream to BRAM interface 61
    input s_axis_bram_61_aclk,
    input s_axis_bram_61_aresetn,
    input s_axis_bram_61_tlast,
    input s_axis_bram_61_tvalid,
    input [S_AXIS_BRAM_61_DMWIDTH/8-1:0] s_axis_bram_61_tkeep,
    input [S_AXIS_BRAM_61_DMWIDTH/8-1:0] s_axis_bram_61_tstrb,
    input [S_AXIS_BRAM_61_DMWIDTH-1:0] s_axis_bram_61_tdata,
    output s_axis_bram_61_tready,
    input [S_AXIS_BRAM_61_ADDR_WIDTH-1:0] ap_bram_iarg_61_addr0,
    input [S_AXIS_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_din0,
    output [S_AXIS_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_dout0,
    input ap_bram_iarg_61_clk0,
    input ap_bram_iarg_61_rst0,
    input [S_AXIS_BRAM_61_WIDTH/8-1:0] ap_bram_iarg_61_we0,
    input ap_bram_iarg_61_en0,
    input [S_AXIS_BRAM_61_ADDR_WIDTH-1:0] ap_bram_iarg_61_addr1,
    input [S_AXIS_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_din1,
    output [S_AXIS_BRAM_61_WIDTH-1:0] ap_bram_iarg_61_dout1,
    input ap_bram_iarg_61_clk1,
    input ap_bram_iarg_61_rst1,
    input [S_AXIS_BRAM_61_WIDTH/8-1:0] ap_bram_iarg_61_we1,
    input ap_bram_iarg_61_en1,
    //input AXI-Stream to BRAM interface 62
    input s_axis_bram_62_aclk,
    input s_axis_bram_62_aresetn,
    input s_axis_bram_62_tlast,
    input s_axis_bram_62_tvalid,
    input [S_AXIS_BRAM_62_DMWIDTH/8-1:0] s_axis_bram_62_tkeep,
    input [S_AXIS_BRAM_62_DMWIDTH/8-1:0] s_axis_bram_62_tstrb,
    input [S_AXIS_BRAM_62_DMWIDTH-1:0] s_axis_bram_62_tdata,
    output s_axis_bram_62_tready,
    input [S_AXIS_BRAM_62_ADDR_WIDTH-1:0] ap_bram_iarg_62_addr0,
    input [S_AXIS_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_din0,
    output [S_AXIS_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_dout0,
    input ap_bram_iarg_62_clk0,
    input ap_bram_iarg_62_rst0,
    input [S_AXIS_BRAM_62_WIDTH/8-1:0] ap_bram_iarg_62_we0,
    input ap_bram_iarg_62_en0,
    input [S_AXIS_BRAM_62_ADDR_WIDTH-1:0] ap_bram_iarg_62_addr1,
    input [S_AXIS_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_din1,
    output [S_AXIS_BRAM_62_WIDTH-1:0] ap_bram_iarg_62_dout1,
    input ap_bram_iarg_62_clk1,
    input ap_bram_iarg_62_rst1,
    input [S_AXIS_BRAM_62_WIDTH/8-1:0] ap_bram_iarg_62_we1,
    input ap_bram_iarg_62_en1,
    //input AXI-Stream to BRAM interface 63
    input s_axis_bram_63_aclk,
    input s_axis_bram_63_aresetn,
    input s_axis_bram_63_tlast,
    input s_axis_bram_63_tvalid,
    input [S_AXIS_BRAM_63_DMWIDTH/8-1:0] s_axis_bram_63_tkeep,
    input [S_AXIS_BRAM_63_DMWIDTH/8-1:0] s_axis_bram_63_tstrb,
    input [S_AXIS_BRAM_63_DMWIDTH-1:0] s_axis_bram_63_tdata,
    output s_axis_bram_63_tready,
    input [S_AXIS_BRAM_63_ADDR_WIDTH-1:0] ap_bram_iarg_63_addr0,
    input [S_AXIS_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_din0,
    output [S_AXIS_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_dout0,
    input ap_bram_iarg_63_clk0,
    input ap_bram_iarg_63_rst0,
    input [S_AXIS_BRAM_63_WIDTH/8-1:0] ap_bram_iarg_63_we0,
    input ap_bram_iarg_63_en0,
    input [S_AXIS_BRAM_63_ADDR_WIDTH-1:0] ap_bram_iarg_63_addr1,
    input [S_AXIS_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_din1,
    output [S_AXIS_BRAM_63_WIDTH-1:0] ap_bram_iarg_63_dout1,
    input ap_bram_iarg_63_clk1,
    input ap_bram_iarg_63_rst1,
    input [S_AXIS_BRAM_63_WIDTH/8-1:0] ap_bram_iarg_63_we1,
    input ap_bram_iarg_63_en1,
    //input AXI-Stream to BRAM interface 64
    input s_axis_bram_64_aclk,
    input s_axis_bram_64_aresetn,
    input s_axis_bram_64_tlast,
    input s_axis_bram_64_tvalid,
    input [S_AXIS_BRAM_64_DMWIDTH/8-1:0] s_axis_bram_64_tkeep,
    input [S_AXIS_BRAM_64_DMWIDTH/8-1:0] s_axis_bram_64_tstrb,
    input [S_AXIS_BRAM_64_DMWIDTH-1:0] s_axis_bram_64_tdata,
    output s_axis_bram_64_tready,
    input [S_AXIS_BRAM_64_ADDR_WIDTH-1:0] ap_bram_iarg_64_addr0,
    input [S_AXIS_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_din0,
    output [S_AXIS_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_dout0,
    input ap_bram_iarg_64_clk0,
    input ap_bram_iarg_64_rst0,
    input [S_AXIS_BRAM_64_WIDTH/8-1:0] ap_bram_iarg_64_we0,
    input ap_bram_iarg_64_en0,
    input [S_AXIS_BRAM_64_ADDR_WIDTH-1:0] ap_bram_iarg_64_addr1,
    input [S_AXIS_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_din1,
    output [S_AXIS_BRAM_64_WIDTH-1:0] ap_bram_iarg_64_dout1,
    input ap_bram_iarg_64_clk1,
    input ap_bram_iarg_64_rst1,
    input [S_AXIS_BRAM_64_WIDTH/8-1:0] ap_bram_iarg_64_we1,
    input ap_bram_iarg_64_en1,
    //input AXI-Stream to BRAM interface 65
    input s_axis_bram_65_aclk,
    input s_axis_bram_65_aresetn,
    input s_axis_bram_65_tlast,
    input s_axis_bram_65_tvalid,
    input [S_AXIS_BRAM_65_DMWIDTH/8-1:0] s_axis_bram_65_tkeep,
    input [S_AXIS_BRAM_65_DMWIDTH/8-1:0] s_axis_bram_65_tstrb,
    input [S_AXIS_BRAM_65_DMWIDTH-1:0] s_axis_bram_65_tdata,
    output s_axis_bram_65_tready,
    input [S_AXIS_BRAM_65_ADDR_WIDTH-1:0] ap_bram_iarg_65_addr0,
    input [S_AXIS_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_din0,
    output [S_AXIS_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_dout0,
    input ap_bram_iarg_65_clk0,
    input ap_bram_iarg_65_rst0,
    input [S_AXIS_BRAM_65_WIDTH/8-1:0] ap_bram_iarg_65_we0,
    input ap_bram_iarg_65_en0,
    input [S_AXIS_BRAM_65_ADDR_WIDTH-1:0] ap_bram_iarg_65_addr1,
    input [S_AXIS_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_din1,
    output [S_AXIS_BRAM_65_WIDTH-1:0] ap_bram_iarg_65_dout1,
    input ap_bram_iarg_65_clk1,
    input ap_bram_iarg_65_rst1,
    input [S_AXIS_BRAM_65_WIDTH/8-1:0] ap_bram_iarg_65_we1,
    input ap_bram_iarg_65_en1,
    //input AXI-Stream to BRAM interface 66
    input s_axis_bram_66_aclk,
    input s_axis_bram_66_aresetn,
    input s_axis_bram_66_tlast,
    input s_axis_bram_66_tvalid,
    input [S_AXIS_BRAM_66_DMWIDTH/8-1:0] s_axis_bram_66_tkeep,
    input [S_AXIS_BRAM_66_DMWIDTH/8-1:0] s_axis_bram_66_tstrb,
    input [S_AXIS_BRAM_66_DMWIDTH-1:0] s_axis_bram_66_tdata,
    output s_axis_bram_66_tready,
    input [S_AXIS_BRAM_66_ADDR_WIDTH-1:0] ap_bram_iarg_66_addr0,
    input [S_AXIS_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_din0,
    output [S_AXIS_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_dout0,
    input ap_bram_iarg_66_clk0,
    input ap_bram_iarg_66_rst0,
    input [S_AXIS_BRAM_66_WIDTH/8-1:0] ap_bram_iarg_66_we0,
    input ap_bram_iarg_66_en0,
    input [S_AXIS_BRAM_66_ADDR_WIDTH-1:0] ap_bram_iarg_66_addr1,
    input [S_AXIS_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_din1,
    output [S_AXIS_BRAM_66_WIDTH-1:0] ap_bram_iarg_66_dout1,
    input ap_bram_iarg_66_clk1,
    input ap_bram_iarg_66_rst1,
    input [S_AXIS_BRAM_66_WIDTH/8-1:0] ap_bram_iarg_66_we1,
    input ap_bram_iarg_66_en1,
    //input AXI-Stream to BRAM interface 67
    input s_axis_bram_67_aclk,
    input s_axis_bram_67_aresetn,
    input s_axis_bram_67_tlast,
    input s_axis_bram_67_tvalid,
    input [S_AXIS_BRAM_67_DMWIDTH/8-1:0] s_axis_bram_67_tkeep,
    input [S_AXIS_BRAM_67_DMWIDTH/8-1:0] s_axis_bram_67_tstrb,
    input [S_AXIS_BRAM_67_DMWIDTH-1:0] s_axis_bram_67_tdata,
    output s_axis_bram_67_tready,
    input [S_AXIS_BRAM_67_ADDR_WIDTH-1:0] ap_bram_iarg_67_addr0,
    input [S_AXIS_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_din0,
    output [S_AXIS_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_dout0,
    input ap_bram_iarg_67_clk0,
    input ap_bram_iarg_67_rst0,
    input [S_AXIS_BRAM_67_WIDTH/8-1:0] ap_bram_iarg_67_we0,
    input ap_bram_iarg_67_en0,
    input [S_AXIS_BRAM_67_ADDR_WIDTH-1:0] ap_bram_iarg_67_addr1,
    input [S_AXIS_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_din1,
    output [S_AXIS_BRAM_67_WIDTH-1:0] ap_bram_iarg_67_dout1,
    input ap_bram_iarg_67_clk1,
    input ap_bram_iarg_67_rst1,
    input [S_AXIS_BRAM_67_WIDTH/8-1:0] ap_bram_iarg_67_we1,
    input ap_bram_iarg_67_en1,
    //input AXI-Stream to BRAM interface 68
    input s_axis_bram_68_aclk,
    input s_axis_bram_68_aresetn,
    input s_axis_bram_68_tlast,
    input s_axis_bram_68_tvalid,
    input [S_AXIS_BRAM_68_DMWIDTH/8-1:0] s_axis_bram_68_tkeep,
    input [S_AXIS_BRAM_68_DMWIDTH/8-1:0] s_axis_bram_68_tstrb,
    input [S_AXIS_BRAM_68_DMWIDTH-1:0] s_axis_bram_68_tdata,
    output s_axis_bram_68_tready,
    input [S_AXIS_BRAM_68_ADDR_WIDTH-1:0] ap_bram_iarg_68_addr0,
    input [S_AXIS_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_din0,
    output [S_AXIS_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_dout0,
    input ap_bram_iarg_68_clk0,
    input ap_bram_iarg_68_rst0,
    input [S_AXIS_BRAM_68_WIDTH/8-1:0] ap_bram_iarg_68_we0,
    input ap_bram_iarg_68_en0,
    input [S_AXIS_BRAM_68_ADDR_WIDTH-1:0] ap_bram_iarg_68_addr1,
    input [S_AXIS_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_din1,
    output [S_AXIS_BRAM_68_WIDTH-1:0] ap_bram_iarg_68_dout1,
    input ap_bram_iarg_68_clk1,
    input ap_bram_iarg_68_rst1,
    input [S_AXIS_BRAM_68_WIDTH/8-1:0] ap_bram_iarg_68_we1,
    input ap_bram_iarg_68_en1,
    //input AXI-Stream to BRAM interface 69
    input s_axis_bram_69_aclk,
    input s_axis_bram_69_aresetn,
    input s_axis_bram_69_tlast,
    input s_axis_bram_69_tvalid,
    input [S_AXIS_BRAM_69_DMWIDTH/8-1:0] s_axis_bram_69_tkeep,
    input [S_AXIS_BRAM_69_DMWIDTH/8-1:0] s_axis_bram_69_tstrb,
    input [S_AXIS_BRAM_69_DMWIDTH-1:0] s_axis_bram_69_tdata,
    output s_axis_bram_69_tready,
    input [S_AXIS_BRAM_69_ADDR_WIDTH-1:0] ap_bram_iarg_69_addr0,
    input [S_AXIS_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_din0,
    output [S_AXIS_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_dout0,
    input ap_bram_iarg_69_clk0,
    input ap_bram_iarg_69_rst0,
    input [S_AXIS_BRAM_69_WIDTH/8-1:0] ap_bram_iarg_69_we0,
    input ap_bram_iarg_69_en0,
    input [S_AXIS_BRAM_69_ADDR_WIDTH-1:0] ap_bram_iarg_69_addr1,
    input [S_AXIS_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_din1,
    output [S_AXIS_BRAM_69_WIDTH-1:0] ap_bram_iarg_69_dout1,
    input ap_bram_iarg_69_clk1,
    input ap_bram_iarg_69_rst1,
    input [S_AXIS_BRAM_69_WIDTH/8-1:0] ap_bram_iarg_69_we1,
    input ap_bram_iarg_69_en1,
    //input AXI-Stream to BRAM interface 70
    input s_axis_bram_70_aclk,
    input s_axis_bram_70_aresetn,
    input s_axis_bram_70_tlast,
    input s_axis_bram_70_tvalid,
    input [S_AXIS_BRAM_70_DMWIDTH/8-1:0] s_axis_bram_70_tkeep,
    input [S_AXIS_BRAM_70_DMWIDTH/8-1:0] s_axis_bram_70_tstrb,
    input [S_AXIS_BRAM_70_DMWIDTH-1:0] s_axis_bram_70_tdata,
    output s_axis_bram_70_tready,
    input [S_AXIS_BRAM_70_ADDR_WIDTH-1:0] ap_bram_iarg_70_addr0,
    input [S_AXIS_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_din0,
    output [S_AXIS_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_dout0,
    input ap_bram_iarg_70_clk0,
    input ap_bram_iarg_70_rst0,
    input [S_AXIS_BRAM_70_WIDTH/8-1:0] ap_bram_iarg_70_we0,
    input ap_bram_iarg_70_en0,
    input [S_AXIS_BRAM_70_ADDR_WIDTH-1:0] ap_bram_iarg_70_addr1,
    input [S_AXIS_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_din1,
    output [S_AXIS_BRAM_70_WIDTH-1:0] ap_bram_iarg_70_dout1,
    input ap_bram_iarg_70_clk1,
    input ap_bram_iarg_70_rst1,
    input [S_AXIS_BRAM_70_WIDTH/8-1:0] ap_bram_iarg_70_we1,
    input ap_bram_iarg_70_en1,
    //input AXI-Stream to BRAM interface 71
    input s_axis_bram_71_aclk,
    input s_axis_bram_71_aresetn,
    input s_axis_bram_71_tlast,
    input s_axis_bram_71_tvalid,
    input [S_AXIS_BRAM_71_DMWIDTH/8-1:0] s_axis_bram_71_tkeep,
    input [S_AXIS_BRAM_71_DMWIDTH/8-1:0] s_axis_bram_71_tstrb,
    input [S_AXIS_BRAM_71_DMWIDTH-1:0] s_axis_bram_71_tdata,
    output s_axis_bram_71_tready,
    input [S_AXIS_BRAM_71_ADDR_WIDTH-1:0] ap_bram_iarg_71_addr0,
    input [S_AXIS_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_din0,
    output [S_AXIS_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_dout0,
    input ap_bram_iarg_71_clk0,
    input ap_bram_iarg_71_rst0,
    input [S_AXIS_BRAM_71_WIDTH/8-1:0] ap_bram_iarg_71_we0,
    input ap_bram_iarg_71_en0,
    input [S_AXIS_BRAM_71_ADDR_WIDTH-1:0] ap_bram_iarg_71_addr1,
    input [S_AXIS_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_din1,
    output [S_AXIS_BRAM_71_WIDTH-1:0] ap_bram_iarg_71_dout1,
    input ap_bram_iarg_71_clk1,
    input ap_bram_iarg_71_rst1,
    input [S_AXIS_BRAM_71_WIDTH/8-1:0] ap_bram_iarg_71_we1,
    input ap_bram_iarg_71_en1,
    //input AXI-Stream to BRAM interface 72
    input s_axis_bram_72_aclk,
    input s_axis_bram_72_aresetn,
    input s_axis_bram_72_tlast,
    input s_axis_bram_72_tvalid,
    input [S_AXIS_BRAM_72_DMWIDTH/8-1:0] s_axis_bram_72_tkeep,
    input [S_AXIS_BRAM_72_DMWIDTH/8-1:0] s_axis_bram_72_tstrb,
    input [S_AXIS_BRAM_72_DMWIDTH-1:0] s_axis_bram_72_tdata,
    output s_axis_bram_72_tready,
    input [S_AXIS_BRAM_72_ADDR_WIDTH-1:0] ap_bram_iarg_72_addr0,
    input [S_AXIS_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_din0,
    output [S_AXIS_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_dout0,
    input ap_bram_iarg_72_clk0,
    input ap_bram_iarg_72_rst0,
    input [S_AXIS_BRAM_72_WIDTH/8-1:0] ap_bram_iarg_72_we0,
    input ap_bram_iarg_72_en0,
    input [S_AXIS_BRAM_72_ADDR_WIDTH-1:0] ap_bram_iarg_72_addr1,
    input [S_AXIS_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_din1,
    output [S_AXIS_BRAM_72_WIDTH-1:0] ap_bram_iarg_72_dout1,
    input ap_bram_iarg_72_clk1,
    input ap_bram_iarg_72_rst1,
    input [S_AXIS_BRAM_72_WIDTH/8-1:0] ap_bram_iarg_72_we1,
    input ap_bram_iarg_72_en1,
    //input AXI-Stream to BRAM interface 73
    input s_axis_bram_73_aclk,
    input s_axis_bram_73_aresetn,
    input s_axis_bram_73_tlast,
    input s_axis_bram_73_tvalid,
    input [S_AXIS_BRAM_73_DMWIDTH/8-1:0] s_axis_bram_73_tkeep,
    input [S_AXIS_BRAM_73_DMWIDTH/8-1:0] s_axis_bram_73_tstrb,
    input [S_AXIS_BRAM_73_DMWIDTH-1:0] s_axis_bram_73_tdata,
    output s_axis_bram_73_tready,
    input [S_AXIS_BRAM_73_ADDR_WIDTH-1:0] ap_bram_iarg_73_addr0,
    input [S_AXIS_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_din0,
    output [S_AXIS_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_dout0,
    input ap_bram_iarg_73_clk0,
    input ap_bram_iarg_73_rst0,
    input [S_AXIS_BRAM_73_WIDTH/8-1:0] ap_bram_iarg_73_we0,
    input ap_bram_iarg_73_en0,
    input [S_AXIS_BRAM_73_ADDR_WIDTH-1:0] ap_bram_iarg_73_addr1,
    input [S_AXIS_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_din1,
    output [S_AXIS_BRAM_73_WIDTH-1:0] ap_bram_iarg_73_dout1,
    input ap_bram_iarg_73_clk1,
    input ap_bram_iarg_73_rst1,
    input [S_AXIS_BRAM_73_WIDTH/8-1:0] ap_bram_iarg_73_we1,
    input ap_bram_iarg_73_en1,
    //input AXI-Stream to BRAM interface 74
    input s_axis_bram_74_aclk,
    input s_axis_bram_74_aresetn,
    input s_axis_bram_74_tlast,
    input s_axis_bram_74_tvalid,
    input [S_AXIS_BRAM_74_DMWIDTH/8-1:0] s_axis_bram_74_tkeep,
    input [S_AXIS_BRAM_74_DMWIDTH/8-1:0] s_axis_bram_74_tstrb,
    input [S_AXIS_BRAM_74_DMWIDTH-1:0] s_axis_bram_74_tdata,
    output s_axis_bram_74_tready,
    input [S_AXIS_BRAM_74_ADDR_WIDTH-1:0] ap_bram_iarg_74_addr0,
    input [S_AXIS_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_din0,
    output [S_AXIS_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_dout0,
    input ap_bram_iarg_74_clk0,
    input ap_bram_iarg_74_rst0,
    input [S_AXIS_BRAM_74_WIDTH/8-1:0] ap_bram_iarg_74_we0,
    input ap_bram_iarg_74_en0,
    input [S_AXIS_BRAM_74_ADDR_WIDTH-1:0] ap_bram_iarg_74_addr1,
    input [S_AXIS_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_din1,
    output [S_AXIS_BRAM_74_WIDTH-1:0] ap_bram_iarg_74_dout1,
    input ap_bram_iarg_74_clk1,
    input ap_bram_iarg_74_rst1,
    input [S_AXIS_BRAM_74_WIDTH/8-1:0] ap_bram_iarg_74_we1,
    input ap_bram_iarg_74_en1,
    //input AXI-Stream to BRAM interface 75
    input s_axis_bram_75_aclk,
    input s_axis_bram_75_aresetn,
    input s_axis_bram_75_tlast,
    input s_axis_bram_75_tvalid,
    input [S_AXIS_BRAM_75_DMWIDTH/8-1:0] s_axis_bram_75_tkeep,
    input [S_AXIS_BRAM_75_DMWIDTH/8-1:0] s_axis_bram_75_tstrb,
    input [S_AXIS_BRAM_75_DMWIDTH-1:0] s_axis_bram_75_tdata,
    output s_axis_bram_75_tready,
    input [S_AXIS_BRAM_75_ADDR_WIDTH-1:0] ap_bram_iarg_75_addr0,
    input [S_AXIS_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_din0,
    output [S_AXIS_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_dout0,
    input ap_bram_iarg_75_clk0,
    input ap_bram_iarg_75_rst0,
    input [S_AXIS_BRAM_75_WIDTH/8-1:0] ap_bram_iarg_75_we0,
    input ap_bram_iarg_75_en0,
    input [S_AXIS_BRAM_75_ADDR_WIDTH-1:0] ap_bram_iarg_75_addr1,
    input [S_AXIS_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_din1,
    output [S_AXIS_BRAM_75_WIDTH-1:0] ap_bram_iarg_75_dout1,
    input ap_bram_iarg_75_clk1,
    input ap_bram_iarg_75_rst1,
    input [S_AXIS_BRAM_75_WIDTH/8-1:0] ap_bram_iarg_75_we1,
    input ap_bram_iarg_75_en1,
    //input AXI-Stream to BRAM interface 76
    input s_axis_bram_76_aclk,
    input s_axis_bram_76_aresetn,
    input s_axis_bram_76_tlast,
    input s_axis_bram_76_tvalid,
    input [S_AXIS_BRAM_76_DMWIDTH/8-1:0] s_axis_bram_76_tkeep,
    input [S_AXIS_BRAM_76_DMWIDTH/8-1:0] s_axis_bram_76_tstrb,
    input [S_AXIS_BRAM_76_DMWIDTH-1:0] s_axis_bram_76_tdata,
    output s_axis_bram_76_tready,
    input [S_AXIS_BRAM_76_ADDR_WIDTH-1:0] ap_bram_iarg_76_addr0,
    input [S_AXIS_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_din0,
    output [S_AXIS_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_dout0,
    input ap_bram_iarg_76_clk0,
    input ap_bram_iarg_76_rst0,
    input [S_AXIS_BRAM_76_WIDTH/8-1:0] ap_bram_iarg_76_we0,
    input ap_bram_iarg_76_en0,
    input [S_AXIS_BRAM_76_ADDR_WIDTH-1:0] ap_bram_iarg_76_addr1,
    input [S_AXIS_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_din1,
    output [S_AXIS_BRAM_76_WIDTH-1:0] ap_bram_iarg_76_dout1,
    input ap_bram_iarg_76_clk1,
    input ap_bram_iarg_76_rst1,
    input [S_AXIS_BRAM_76_WIDTH/8-1:0] ap_bram_iarg_76_we1,
    input ap_bram_iarg_76_en1,
    //input AXI-Stream to BRAM interface 77
    input s_axis_bram_77_aclk,
    input s_axis_bram_77_aresetn,
    input s_axis_bram_77_tlast,
    input s_axis_bram_77_tvalid,
    input [S_AXIS_BRAM_77_DMWIDTH/8-1:0] s_axis_bram_77_tkeep,
    input [S_AXIS_BRAM_77_DMWIDTH/8-1:0] s_axis_bram_77_tstrb,
    input [S_AXIS_BRAM_77_DMWIDTH-1:0] s_axis_bram_77_tdata,
    output s_axis_bram_77_tready,
    input [S_AXIS_BRAM_77_ADDR_WIDTH-1:0] ap_bram_iarg_77_addr0,
    input [S_AXIS_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_din0,
    output [S_AXIS_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_dout0,
    input ap_bram_iarg_77_clk0,
    input ap_bram_iarg_77_rst0,
    input [S_AXIS_BRAM_77_WIDTH/8-1:0] ap_bram_iarg_77_we0,
    input ap_bram_iarg_77_en0,
    input [S_AXIS_BRAM_77_ADDR_WIDTH-1:0] ap_bram_iarg_77_addr1,
    input [S_AXIS_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_din1,
    output [S_AXIS_BRAM_77_WIDTH-1:0] ap_bram_iarg_77_dout1,
    input ap_bram_iarg_77_clk1,
    input ap_bram_iarg_77_rst1,
    input [S_AXIS_BRAM_77_WIDTH/8-1:0] ap_bram_iarg_77_we1,
    input ap_bram_iarg_77_en1,
    //input AXI-Stream to BRAM interface 78
    input s_axis_bram_78_aclk,
    input s_axis_bram_78_aresetn,
    input s_axis_bram_78_tlast,
    input s_axis_bram_78_tvalid,
    input [S_AXIS_BRAM_78_DMWIDTH/8-1:0] s_axis_bram_78_tkeep,
    input [S_AXIS_BRAM_78_DMWIDTH/8-1:0] s_axis_bram_78_tstrb,
    input [S_AXIS_BRAM_78_DMWIDTH-1:0] s_axis_bram_78_tdata,
    output s_axis_bram_78_tready,
    input [S_AXIS_BRAM_78_ADDR_WIDTH-1:0] ap_bram_iarg_78_addr0,
    input [S_AXIS_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_din0,
    output [S_AXIS_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_dout0,
    input ap_bram_iarg_78_clk0,
    input ap_bram_iarg_78_rst0,
    input [S_AXIS_BRAM_78_WIDTH/8-1:0] ap_bram_iarg_78_we0,
    input ap_bram_iarg_78_en0,
    input [S_AXIS_BRAM_78_ADDR_WIDTH-1:0] ap_bram_iarg_78_addr1,
    input [S_AXIS_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_din1,
    output [S_AXIS_BRAM_78_WIDTH-1:0] ap_bram_iarg_78_dout1,
    input ap_bram_iarg_78_clk1,
    input ap_bram_iarg_78_rst1,
    input [S_AXIS_BRAM_78_WIDTH/8-1:0] ap_bram_iarg_78_we1,
    input ap_bram_iarg_78_en1,
    //input AXI-Stream to BRAM interface 79
    input s_axis_bram_79_aclk,
    input s_axis_bram_79_aresetn,
    input s_axis_bram_79_tlast,
    input s_axis_bram_79_tvalid,
    input [S_AXIS_BRAM_79_DMWIDTH/8-1:0] s_axis_bram_79_tkeep,
    input [S_AXIS_BRAM_79_DMWIDTH/8-1:0] s_axis_bram_79_tstrb,
    input [S_AXIS_BRAM_79_DMWIDTH-1:0] s_axis_bram_79_tdata,
    output s_axis_bram_79_tready,
    input [S_AXIS_BRAM_79_ADDR_WIDTH-1:0] ap_bram_iarg_79_addr0,
    input [S_AXIS_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_din0,
    output [S_AXIS_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_dout0,
    input ap_bram_iarg_79_clk0,
    input ap_bram_iarg_79_rst0,
    input [S_AXIS_BRAM_79_WIDTH/8-1:0] ap_bram_iarg_79_we0,
    input ap_bram_iarg_79_en0,
    input [S_AXIS_BRAM_79_ADDR_WIDTH-1:0] ap_bram_iarg_79_addr1,
    input [S_AXIS_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_din1,
    output [S_AXIS_BRAM_79_WIDTH-1:0] ap_bram_iarg_79_dout1,
    input ap_bram_iarg_79_clk1,
    input ap_bram_iarg_79_rst1,
    input [S_AXIS_BRAM_79_WIDTH/8-1:0] ap_bram_iarg_79_we1,
    input ap_bram_iarg_79_en1,
    //input AXI-Stream to BRAM interface 80
    input s_axis_bram_80_aclk,
    input s_axis_bram_80_aresetn,
    input s_axis_bram_80_tlast,
    input s_axis_bram_80_tvalid,
    input [S_AXIS_BRAM_80_DMWIDTH/8-1:0] s_axis_bram_80_tkeep,
    input [S_AXIS_BRAM_80_DMWIDTH/8-1:0] s_axis_bram_80_tstrb,
    input [S_AXIS_BRAM_80_DMWIDTH-1:0] s_axis_bram_80_tdata,
    output s_axis_bram_80_tready,
    input [S_AXIS_BRAM_80_ADDR_WIDTH-1:0] ap_bram_iarg_80_addr0,
    input [S_AXIS_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_din0,
    output [S_AXIS_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_dout0,
    input ap_bram_iarg_80_clk0,
    input ap_bram_iarg_80_rst0,
    input [S_AXIS_BRAM_80_WIDTH/8-1:0] ap_bram_iarg_80_we0,
    input ap_bram_iarg_80_en0,
    input [S_AXIS_BRAM_80_ADDR_WIDTH-1:0] ap_bram_iarg_80_addr1,
    input [S_AXIS_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_din1,
    output [S_AXIS_BRAM_80_WIDTH-1:0] ap_bram_iarg_80_dout1,
    input ap_bram_iarg_80_clk1,
    input ap_bram_iarg_80_rst1,
    input [S_AXIS_BRAM_80_WIDTH/8-1:0] ap_bram_iarg_80_we1,
    input ap_bram_iarg_80_en1,
    //input AXI-Stream to BRAM interface 81
    input s_axis_bram_81_aclk,
    input s_axis_bram_81_aresetn,
    input s_axis_bram_81_tlast,
    input s_axis_bram_81_tvalid,
    input [S_AXIS_BRAM_81_DMWIDTH/8-1:0] s_axis_bram_81_tkeep,
    input [S_AXIS_BRAM_81_DMWIDTH/8-1:0] s_axis_bram_81_tstrb,
    input [S_AXIS_BRAM_81_DMWIDTH-1:0] s_axis_bram_81_tdata,
    output s_axis_bram_81_tready,
    input [S_AXIS_BRAM_81_ADDR_WIDTH-1:0] ap_bram_iarg_81_addr0,
    input [S_AXIS_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_din0,
    output [S_AXIS_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_dout0,
    input ap_bram_iarg_81_clk0,
    input ap_bram_iarg_81_rst0,
    input [S_AXIS_BRAM_81_WIDTH/8-1:0] ap_bram_iarg_81_we0,
    input ap_bram_iarg_81_en0,
    input [S_AXIS_BRAM_81_ADDR_WIDTH-1:0] ap_bram_iarg_81_addr1,
    input [S_AXIS_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_din1,
    output [S_AXIS_BRAM_81_WIDTH-1:0] ap_bram_iarg_81_dout1,
    input ap_bram_iarg_81_clk1,
    input ap_bram_iarg_81_rst1,
    input [S_AXIS_BRAM_81_WIDTH/8-1:0] ap_bram_iarg_81_we1,
    input ap_bram_iarg_81_en1,
    //input AXI-Stream to BRAM interface 82
    input s_axis_bram_82_aclk,
    input s_axis_bram_82_aresetn,
    input s_axis_bram_82_tlast,
    input s_axis_bram_82_tvalid,
    input [S_AXIS_BRAM_82_DMWIDTH/8-1:0] s_axis_bram_82_tkeep,
    input [S_AXIS_BRAM_82_DMWIDTH/8-1:0] s_axis_bram_82_tstrb,
    input [S_AXIS_BRAM_82_DMWIDTH-1:0] s_axis_bram_82_tdata,
    output s_axis_bram_82_tready,
    input [S_AXIS_BRAM_82_ADDR_WIDTH-1:0] ap_bram_iarg_82_addr0,
    input [S_AXIS_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_din0,
    output [S_AXIS_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_dout0,
    input ap_bram_iarg_82_clk0,
    input ap_bram_iarg_82_rst0,
    input [S_AXIS_BRAM_82_WIDTH/8-1:0] ap_bram_iarg_82_we0,
    input ap_bram_iarg_82_en0,
    input [S_AXIS_BRAM_82_ADDR_WIDTH-1:0] ap_bram_iarg_82_addr1,
    input [S_AXIS_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_din1,
    output [S_AXIS_BRAM_82_WIDTH-1:0] ap_bram_iarg_82_dout1,
    input ap_bram_iarg_82_clk1,
    input ap_bram_iarg_82_rst1,
    input [S_AXIS_BRAM_82_WIDTH/8-1:0] ap_bram_iarg_82_we1,
    input ap_bram_iarg_82_en1,
    //input AXI-Stream to BRAM interface 83
    input s_axis_bram_83_aclk,
    input s_axis_bram_83_aresetn,
    input s_axis_bram_83_tlast,
    input s_axis_bram_83_tvalid,
    input [S_AXIS_BRAM_83_DMWIDTH/8-1:0] s_axis_bram_83_tkeep,
    input [S_AXIS_BRAM_83_DMWIDTH/8-1:0] s_axis_bram_83_tstrb,
    input [S_AXIS_BRAM_83_DMWIDTH-1:0] s_axis_bram_83_tdata,
    output s_axis_bram_83_tready,
    input [S_AXIS_BRAM_83_ADDR_WIDTH-1:0] ap_bram_iarg_83_addr0,
    input [S_AXIS_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_din0,
    output [S_AXIS_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_dout0,
    input ap_bram_iarg_83_clk0,
    input ap_bram_iarg_83_rst0,
    input [S_AXIS_BRAM_83_WIDTH/8-1:0] ap_bram_iarg_83_we0,
    input ap_bram_iarg_83_en0,
    input [S_AXIS_BRAM_83_ADDR_WIDTH-1:0] ap_bram_iarg_83_addr1,
    input [S_AXIS_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_din1,
    output [S_AXIS_BRAM_83_WIDTH-1:0] ap_bram_iarg_83_dout1,
    input ap_bram_iarg_83_clk1,
    input ap_bram_iarg_83_rst1,
    input [S_AXIS_BRAM_83_WIDTH/8-1:0] ap_bram_iarg_83_we1,
    input ap_bram_iarg_83_en1,
    //input AXI-Stream to BRAM interface 84
    input s_axis_bram_84_aclk,
    input s_axis_bram_84_aresetn,
    input s_axis_bram_84_tlast,
    input s_axis_bram_84_tvalid,
    input [S_AXIS_BRAM_84_DMWIDTH/8-1:0] s_axis_bram_84_tkeep,
    input [S_AXIS_BRAM_84_DMWIDTH/8-1:0] s_axis_bram_84_tstrb,
    input [S_AXIS_BRAM_84_DMWIDTH-1:0] s_axis_bram_84_tdata,
    output s_axis_bram_84_tready,
    input [S_AXIS_BRAM_84_ADDR_WIDTH-1:0] ap_bram_iarg_84_addr0,
    input [S_AXIS_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_din0,
    output [S_AXIS_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_dout0,
    input ap_bram_iarg_84_clk0,
    input ap_bram_iarg_84_rst0,
    input [S_AXIS_BRAM_84_WIDTH/8-1:0] ap_bram_iarg_84_we0,
    input ap_bram_iarg_84_en0,
    input [S_AXIS_BRAM_84_ADDR_WIDTH-1:0] ap_bram_iarg_84_addr1,
    input [S_AXIS_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_din1,
    output [S_AXIS_BRAM_84_WIDTH-1:0] ap_bram_iarg_84_dout1,
    input ap_bram_iarg_84_clk1,
    input ap_bram_iarg_84_rst1,
    input [S_AXIS_BRAM_84_WIDTH/8-1:0] ap_bram_iarg_84_we1,
    input ap_bram_iarg_84_en1,
    //input AXI-Stream to BRAM interface 85
    input s_axis_bram_85_aclk,
    input s_axis_bram_85_aresetn,
    input s_axis_bram_85_tlast,
    input s_axis_bram_85_tvalid,
    input [S_AXIS_BRAM_85_DMWIDTH/8-1:0] s_axis_bram_85_tkeep,
    input [S_AXIS_BRAM_85_DMWIDTH/8-1:0] s_axis_bram_85_tstrb,
    input [S_AXIS_BRAM_85_DMWIDTH-1:0] s_axis_bram_85_tdata,
    output s_axis_bram_85_tready,
    input [S_AXIS_BRAM_85_ADDR_WIDTH-1:0] ap_bram_iarg_85_addr0,
    input [S_AXIS_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_din0,
    output [S_AXIS_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_dout0,
    input ap_bram_iarg_85_clk0,
    input ap_bram_iarg_85_rst0,
    input [S_AXIS_BRAM_85_WIDTH/8-1:0] ap_bram_iarg_85_we0,
    input ap_bram_iarg_85_en0,
    input [S_AXIS_BRAM_85_ADDR_WIDTH-1:0] ap_bram_iarg_85_addr1,
    input [S_AXIS_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_din1,
    output [S_AXIS_BRAM_85_WIDTH-1:0] ap_bram_iarg_85_dout1,
    input ap_bram_iarg_85_clk1,
    input ap_bram_iarg_85_rst1,
    input [S_AXIS_BRAM_85_WIDTH/8-1:0] ap_bram_iarg_85_we1,
    input ap_bram_iarg_85_en1,
    //input AXI-Stream to BRAM interface 86
    input s_axis_bram_86_aclk,
    input s_axis_bram_86_aresetn,
    input s_axis_bram_86_tlast,
    input s_axis_bram_86_tvalid,
    input [S_AXIS_BRAM_86_DMWIDTH/8-1:0] s_axis_bram_86_tkeep,
    input [S_AXIS_BRAM_86_DMWIDTH/8-1:0] s_axis_bram_86_tstrb,
    input [S_AXIS_BRAM_86_DMWIDTH-1:0] s_axis_bram_86_tdata,
    output s_axis_bram_86_tready,
    input [S_AXIS_BRAM_86_ADDR_WIDTH-1:0] ap_bram_iarg_86_addr0,
    input [S_AXIS_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_din0,
    output [S_AXIS_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_dout0,
    input ap_bram_iarg_86_clk0,
    input ap_bram_iarg_86_rst0,
    input [S_AXIS_BRAM_86_WIDTH/8-1:0] ap_bram_iarg_86_we0,
    input ap_bram_iarg_86_en0,
    input [S_AXIS_BRAM_86_ADDR_WIDTH-1:0] ap_bram_iarg_86_addr1,
    input [S_AXIS_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_din1,
    output [S_AXIS_BRAM_86_WIDTH-1:0] ap_bram_iarg_86_dout1,
    input ap_bram_iarg_86_clk1,
    input ap_bram_iarg_86_rst1,
    input [S_AXIS_BRAM_86_WIDTH/8-1:0] ap_bram_iarg_86_we1,
    input ap_bram_iarg_86_en1,
    //input AXI-Stream to BRAM interface 87
    input s_axis_bram_87_aclk,
    input s_axis_bram_87_aresetn,
    input s_axis_bram_87_tlast,
    input s_axis_bram_87_tvalid,
    input [S_AXIS_BRAM_87_DMWIDTH/8-1:0] s_axis_bram_87_tkeep,
    input [S_AXIS_BRAM_87_DMWIDTH/8-1:0] s_axis_bram_87_tstrb,
    input [S_AXIS_BRAM_87_DMWIDTH-1:0] s_axis_bram_87_tdata,
    output s_axis_bram_87_tready,
    input [S_AXIS_BRAM_87_ADDR_WIDTH-1:0] ap_bram_iarg_87_addr0,
    input [S_AXIS_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_din0,
    output [S_AXIS_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_dout0,
    input ap_bram_iarg_87_clk0,
    input ap_bram_iarg_87_rst0,
    input [S_AXIS_BRAM_87_WIDTH/8-1:0] ap_bram_iarg_87_we0,
    input ap_bram_iarg_87_en0,
    input [S_AXIS_BRAM_87_ADDR_WIDTH-1:0] ap_bram_iarg_87_addr1,
    input [S_AXIS_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_din1,
    output [S_AXIS_BRAM_87_WIDTH-1:0] ap_bram_iarg_87_dout1,
    input ap_bram_iarg_87_clk1,
    input ap_bram_iarg_87_rst1,
    input [S_AXIS_BRAM_87_WIDTH/8-1:0] ap_bram_iarg_87_we1,
    input ap_bram_iarg_87_en1,
    //input AXI-Stream to BRAM interface 88
    input s_axis_bram_88_aclk,
    input s_axis_bram_88_aresetn,
    input s_axis_bram_88_tlast,
    input s_axis_bram_88_tvalid,
    input [S_AXIS_BRAM_88_DMWIDTH/8-1:0] s_axis_bram_88_tkeep,
    input [S_AXIS_BRAM_88_DMWIDTH/8-1:0] s_axis_bram_88_tstrb,
    input [S_AXIS_BRAM_88_DMWIDTH-1:0] s_axis_bram_88_tdata,
    output s_axis_bram_88_tready,
    input [S_AXIS_BRAM_88_ADDR_WIDTH-1:0] ap_bram_iarg_88_addr0,
    input [S_AXIS_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_din0,
    output [S_AXIS_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_dout0,
    input ap_bram_iarg_88_clk0,
    input ap_bram_iarg_88_rst0,
    input [S_AXIS_BRAM_88_WIDTH/8-1:0] ap_bram_iarg_88_we0,
    input ap_bram_iarg_88_en0,
    input [S_AXIS_BRAM_88_ADDR_WIDTH-1:0] ap_bram_iarg_88_addr1,
    input [S_AXIS_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_din1,
    output [S_AXIS_BRAM_88_WIDTH-1:0] ap_bram_iarg_88_dout1,
    input ap_bram_iarg_88_clk1,
    input ap_bram_iarg_88_rst1,
    input [S_AXIS_BRAM_88_WIDTH/8-1:0] ap_bram_iarg_88_we1,
    input ap_bram_iarg_88_en1,
    //input AXI-Stream to BRAM interface 89
    input s_axis_bram_89_aclk,
    input s_axis_bram_89_aresetn,
    input s_axis_bram_89_tlast,
    input s_axis_bram_89_tvalid,
    input [S_AXIS_BRAM_89_DMWIDTH/8-1:0] s_axis_bram_89_tkeep,
    input [S_AXIS_BRAM_89_DMWIDTH/8-1:0] s_axis_bram_89_tstrb,
    input [S_AXIS_BRAM_89_DMWIDTH-1:0] s_axis_bram_89_tdata,
    output s_axis_bram_89_tready,
    input [S_AXIS_BRAM_89_ADDR_WIDTH-1:0] ap_bram_iarg_89_addr0,
    input [S_AXIS_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_din0,
    output [S_AXIS_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_dout0,
    input ap_bram_iarg_89_clk0,
    input ap_bram_iarg_89_rst0,
    input [S_AXIS_BRAM_89_WIDTH/8-1:0] ap_bram_iarg_89_we0,
    input ap_bram_iarg_89_en0,
    input [S_AXIS_BRAM_89_ADDR_WIDTH-1:0] ap_bram_iarg_89_addr1,
    input [S_AXIS_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_din1,
    output [S_AXIS_BRAM_89_WIDTH-1:0] ap_bram_iarg_89_dout1,
    input ap_bram_iarg_89_clk1,
    input ap_bram_iarg_89_rst1,
    input [S_AXIS_BRAM_89_WIDTH/8-1:0] ap_bram_iarg_89_we1,
    input ap_bram_iarg_89_en1,
    //input AXI-Stream to BRAM interface 90
    input s_axis_bram_90_aclk,
    input s_axis_bram_90_aresetn,
    input s_axis_bram_90_tlast,
    input s_axis_bram_90_tvalid,
    input [S_AXIS_BRAM_90_DMWIDTH/8-1:0] s_axis_bram_90_tkeep,
    input [S_AXIS_BRAM_90_DMWIDTH/8-1:0] s_axis_bram_90_tstrb,
    input [S_AXIS_BRAM_90_DMWIDTH-1:0] s_axis_bram_90_tdata,
    output s_axis_bram_90_tready,
    input [S_AXIS_BRAM_90_ADDR_WIDTH-1:0] ap_bram_iarg_90_addr0,
    input [S_AXIS_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_din0,
    output [S_AXIS_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_dout0,
    input ap_bram_iarg_90_clk0,
    input ap_bram_iarg_90_rst0,
    input [S_AXIS_BRAM_90_WIDTH/8-1:0] ap_bram_iarg_90_we0,
    input ap_bram_iarg_90_en0,
    input [S_AXIS_BRAM_90_ADDR_WIDTH-1:0] ap_bram_iarg_90_addr1,
    input [S_AXIS_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_din1,
    output [S_AXIS_BRAM_90_WIDTH-1:0] ap_bram_iarg_90_dout1,
    input ap_bram_iarg_90_clk1,
    input ap_bram_iarg_90_rst1,
    input [S_AXIS_BRAM_90_WIDTH/8-1:0] ap_bram_iarg_90_we1,
    input ap_bram_iarg_90_en1,
    //input AXI-Stream to BRAM interface 91
    input s_axis_bram_91_aclk,
    input s_axis_bram_91_aresetn,
    input s_axis_bram_91_tlast,
    input s_axis_bram_91_tvalid,
    input [S_AXIS_BRAM_91_DMWIDTH/8-1:0] s_axis_bram_91_tkeep,
    input [S_AXIS_BRAM_91_DMWIDTH/8-1:0] s_axis_bram_91_tstrb,
    input [S_AXIS_BRAM_91_DMWIDTH-1:0] s_axis_bram_91_tdata,
    output s_axis_bram_91_tready,
    input [S_AXIS_BRAM_91_ADDR_WIDTH-1:0] ap_bram_iarg_91_addr0,
    input [S_AXIS_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_din0,
    output [S_AXIS_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_dout0,
    input ap_bram_iarg_91_clk0,
    input ap_bram_iarg_91_rst0,
    input [S_AXIS_BRAM_91_WIDTH/8-1:0] ap_bram_iarg_91_we0,
    input ap_bram_iarg_91_en0,
    input [S_AXIS_BRAM_91_ADDR_WIDTH-1:0] ap_bram_iarg_91_addr1,
    input [S_AXIS_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_din1,
    output [S_AXIS_BRAM_91_WIDTH-1:0] ap_bram_iarg_91_dout1,
    input ap_bram_iarg_91_clk1,
    input ap_bram_iarg_91_rst1,
    input [S_AXIS_BRAM_91_WIDTH/8-1:0] ap_bram_iarg_91_we1,
    input ap_bram_iarg_91_en1,
    //input AXI-Stream to BRAM interface 92
    input s_axis_bram_92_aclk,
    input s_axis_bram_92_aresetn,
    input s_axis_bram_92_tlast,
    input s_axis_bram_92_tvalid,
    input [S_AXIS_BRAM_92_DMWIDTH/8-1:0] s_axis_bram_92_tkeep,
    input [S_AXIS_BRAM_92_DMWIDTH/8-1:0] s_axis_bram_92_tstrb,
    input [S_AXIS_BRAM_92_DMWIDTH-1:0] s_axis_bram_92_tdata,
    output s_axis_bram_92_tready,
    input [S_AXIS_BRAM_92_ADDR_WIDTH-1:0] ap_bram_iarg_92_addr0,
    input [S_AXIS_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_din0,
    output [S_AXIS_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_dout0,
    input ap_bram_iarg_92_clk0,
    input ap_bram_iarg_92_rst0,
    input [S_AXIS_BRAM_92_WIDTH/8-1:0] ap_bram_iarg_92_we0,
    input ap_bram_iarg_92_en0,
    input [S_AXIS_BRAM_92_ADDR_WIDTH-1:0] ap_bram_iarg_92_addr1,
    input [S_AXIS_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_din1,
    output [S_AXIS_BRAM_92_WIDTH-1:0] ap_bram_iarg_92_dout1,
    input ap_bram_iarg_92_clk1,
    input ap_bram_iarg_92_rst1,
    input [S_AXIS_BRAM_92_WIDTH/8-1:0] ap_bram_iarg_92_we1,
    input ap_bram_iarg_92_en1,
    //input AXI-Stream to BRAM interface 93
    input s_axis_bram_93_aclk,
    input s_axis_bram_93_aresetn,
    input s_axis_bram_93_tlast,
    input s_axis_bram_93_tvalid,
    input [S_AXIS_BRAM_93_DMWIDTH/8-1:0] s_axis_bram_93_tkeep,
    input [S_AXIS_BRAM_93_DMWIDTH/8-1:0] s_axis_bram_93_tstrb,
    input [S_AXIS_BRAM_93_DMWIDTH-1:0] s_axis_bram_93_tdata,
    output s_axis_bram_93_tready,
    input [S_AXIS_BRAM_93_ADDR_WIDTH-1:0] ap_bram_iarg_93_addr0,
    input [S_AXIS_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_din0,
    output [S_AXIS_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_dout0,
    input ap_bram_iarg_93_clk0,
    input ap_bram_iarg_93_rst0,
    input [S_AXIS_BRAM_93_WIDTH/8-1:0] ap_bram_iarg_93_we0,
    input ap_bram_iarg_93_en0,
    input [S_AXIS_BRAM_93_ADDR_WIDTH-1:0] ap_bram_iarg_93_addr1,
    input [S_AXIS_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_din1,
    output [S_AXIS_BRAM_93_WIDTH-1:0] ap_bram_iarg_93_dout1,
    input ap_bram_iarg_93_clk1,
    input ap_bram_iarg_93_rst1,
    input [S_AXIS_BRAM_93_WIDTH/8-1:0] ap_bram_iarg_93_we1,
    input ap_bram_iarg_93_en1,
    //input AXI-Stream to BRAM interface 94
    input s_axis_bram_94_aclk,
    input s_axis_bram_94_aresetn,
    input s_axis_bram_94_tlast,
    input s_axis_bram_94_tvalid,
    input [S_AXIS_BRAM_94_DMWIDTH/8-1:0] s_axis_bram_94_tkeep,
    input [S_AXIS_BRAM_94_DMWIDTH/8-1:0] s_axis_bram_94_tstrb,
    input [S_AXIS_BRAM_94_DMWIDTH-1:0] s_axis_bram_94_tdata,
    output s_axis_bram_94_tready,
    input [S_AXIS_BRAM_94_ADDR_WIDTH-1:0] ap_bram_iarg_94_addr0,
    input [S_AXIS_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_din0,
    output [S_AXIS_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_dout0,
    input ap_bram_iarg_94_clk0,
    input ap_bram_iarg_94_rst0,
    input [S_AXIS_BRAM_94_WIDTH/8-1:0] ap_bram_iarg_94_we0,
    input ap_bram_iarg_94_en0,
    input [S_AXIS_BRAM_94_ADDR_WIDTH-1:0] ap_bram_iarg_94_addr1,
    input [S_AXIS_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_din1,
    output [S_AXIS_BRAM_94_WIDTH-1:0] ap_bram_iarg_94_dout1,
    input ap_bram_iarg_94_clk1,
    input ap_bram_iarg_94_rst1,
    input [S_AXIS_BRAM_94_WIDTH/8-1:0] ap_bram_iarg_94_we1,
    input ap_bram_iarg_94_en1,
    //input AXI-Stream to BRAM interface 95
    input s_axis_bram_95_aclk,
    input s_axis_bram_95_aresetn,
    input s_axis_bram_95_tlast,
    input s_axis_bram_95_tvalid,
    input [S_AXIS_BRAM_95_DMWIDTH/8-1:0] s_axis_bram_95_tkeep,
    input [S_AXIS_BRAM_95_DMWIDTH/8-1:0] s_axis_bram_95_tstrb,
    input [S_AXIS_BRAM_95_DMWIDTH-1:0] s_axis_bram_95_tdata,
    output s_axis_bram_95_tready,
    input [S_AXIS_BRAM_95_ADDR_WIDTH-1:0] ap_bram_iarg_95_addr0,
    input [S_AXIS_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_din0,
    output [S_AXIS_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_dout0,
    input ap_bram_iarg_95_clk0,
    input ap_bram_iarg_95_rst0,
    input [S_AXIS_BRAM_95_WIDTH/8-1:0] ap_bram_iarg_95_we0,
    input ap_bram_iarg_95_en0,
    input [S_AXIS_BRAM_95_ADDR_WIDTH-1:0] ap_bram_iarg_95_addr1,
    input [S_AXIS_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_din1,
    output [S_AXIS_BRAM_95_WIDTH-1:0] ap_bram_iarg_95_dout1,
    input ap_bram_iarg_95_clk1,
    input ap_bram_iarg_95_rst1,
    input [S_AXIS_BRAM_95_WIDTH/8-1:0] ap_bram_iarg_95_we1,
    input ap_bram_iarg_95_en1,
    //input AXI-Stream to BRAM interface 96
    input s_axis_bram_96_aclk,
    input s_axis_bram_96_aresetn,
    input s_axis_bram_96_tlast,
    input s_axis_bram_96_tvalid,
    input [S_AXIS_BRAM_96_DMWIDTH/8-1:0] s_axis_bram_96_tkeep,
    input [S_AXIS_BRAM_96_DMWIDTH/8-1:0] s_axis_bram_96_tstrb,
    input [S_AXIS_BRAM_96_DMWIDTH-1:0] s_axis_bram_96_tdata,
    output s_axis_bram_96_tready,
    input [S_AXIS_BRAM_96_ADDR_WIDTH-1:0] ap_bram_iarg_96_addr0,
    input [S_AXIS_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_din0,
    output [S_AXIS_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_dout0,
    input ap_bram_iarg_96_clk0,
    input ap_bram_iarg_96_rst0,
    input [S_AXIS_BRAM_96_WIDTH/8-1:0] ap_bram_iarg_96_we0,
    input ap_bram_iarg_96_en0,
    input [S_AXIS_BRAM_96_ADDR_WIDTH-1:0] ap_bram_iarg_96_addr1,
    input [S_AXIS_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_din1,
    output [S_AXIS_BRAM_96_WIDTH-1:0] ap_bram_iarg_96_dout1,
    input ap_bram_iarg_96_clk1,
    input ap_bram_iarg_96_rst1,
    input [S_AXIS_BRAM_96_WIDTH/8-1:0] ap_bram_iarg_96_we1,
    input ap_bram_iarg_96_en1,
    //input AXI-Stream to BRAM interface 97
    input s_axis_bram_97_aclk,
    input s_axis_bram_97_aresetn,
    input s_axis_bram_97_tlast,
    input s_axis_bram_97_tvalid,
    input [S_AXIS_BRAM_97_DMWIDTH/8-1:0] s_axis_bram_97_tkeep,
    input [S_AXIS_BRAM_97_DMWIDTH/8-1:0] s_axis_bram_97_tstrb,
    input [S_AXIS_BRAM_97_DMWIDTH-1:0] s_axis_bram_97_tdata,
    output s_axis_bram_97_tready,
    input [S_AXIS_BRAM_97_ADDR_WIDTH-1:0] ap_bram_iarg_97_addr0,
    input [S_AXIS_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_din0,
    output [S_AXIS_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_dout0,
    input ap_bram_iarg_97_clk0,
    input ap_bram_iarg_97_rst0,
    input [S_AXIS_BRAM_97_WIDTH/8-1:0] ap_bram_iarg_97_we0,
    input ap_bram_iarg_97_en0,
    input [S_AXIS_BRAM_97_ADDR_WIDTH-1:0] ap_bram_iarg_97_addr1,
    input [S_AXIS_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_din1,
    output [S_AXIS_BRAM_97_WIDTH-1:0] ap_bram_iarg_97_dout1,
    input ap_bram_iarg_97_clk1,
    input ap_bram_iarg_97_rst1,
    input [S_AXIS_BRAM_97_WIDTH/8-1:0] ap_bram_iarg_97_we1,
    input ap_bram_iarg_97_en1,
    //input AXI-Stream to BRAM interface 98
    input s_axis_bram_98_aclk,
    input s_axis_bram_98_aresetn,
    input s_axis_bram_98_tlast,
    input s_axis_bram_98_tvalid,
    input [S_AXIS_BRAM_98_DMWIDTH/8-1:0] s_axis_bram_98_tkeep,
    input [S_AXIS_BRAM_98_DMWIDTH/8-1:0] s_axis_bram_98_tstrb,
    input [S_AXIS_BRAM_98_DMWIDTH-1:0] s_axis_bram_98_tdata,
    output s_axis_bram_98_tready,
    input [S_AXIS_BRAM_98_ADDR_WIDTH-1:0] ap_bram_iarg_98_addr0,
    input [S_AXIS_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_din0,
    output [S_AXIS_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_dout0,
    input ap_bram_iarg_98_clk0,
    input ap_bram_iarg_98_rst0,
    input [S_AXIS_BRAM_98_WIDTH/8-1:0] ap_bram_iarg_98_we0,
    input ap_bram_iarg_98_en0,
    input [S_AXIS_BRAM_98_ADDR_WIDTH-1:0] ap_bram_iarg_98_addr1,
    input [S_AXIS_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_din1,
    output [S_AXIS_BRAM_98_WIDTH-1:0] ap_bram_iarg_98_dout1,
    input ap_bram_iarg_98_clk1,
    input ap_bram_iarg_98_rst1,
    input [S_AXIS_BRAM_98_WIDTH/8-1:0] ap_bram_iarg_98_we1,
    input ap_bram_iarg_98_en1,
    //input AXI-Stream to BRAM interface 99
    input s_axis_bram_99_aclk,
    input s_axis_bram_99_aresetn,
    input s_axis_bram_99_tlast,
    input s_axis_bram_99_tvalid,
    input [S_AXIS_BRAM_99_DMWIDTH/8-1:0] s_axis_bram_99_tkeep,
    input [S_AXIS_BRAM_99_DMWIDTH/8-1:0] s_axis_bram_99_tstrb,
    input [S_AXIS_BRAM_99_DMWIDTH-1:0] s_axis_bram_99_tdata,
    output s_axis_bram_99_tready,
    input [S_AXIS_BRAM_99_ADDR_WIDTH-1:0] ap_bram_iarg_99_addr0,
    input [S_AXIS_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_din0,
    output [S_AXIS_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_dout0,
    input ap_bram_iarg_99_clk0,
    input ap_bram_iarg_99_rst0,
    input [S_AXIS_BRAM_99_WIDTH/8-1:0] ap_bram_iarg_99_we0,
    input ap_bram_iarg_99_en0,
    input [S_AXIS_BRAM_99_ADDR_WIDTH-1:0] ap_bram_iarg_99_addr1,
    input [S_AXIS_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_din1,
    output [S_AXIS_BRAM_99_WIDTH-1:0] ap_bram_iarg_99_dout1,
    input ap_bram_iarg_99_clk1,
    input ap_bram_iarg_99_rst1,
    input [S_AXIS_BRAM_99_WIDTH/8-1:0] ap_bram_iarg_99_we1,
    input ap_bram_iarg_99_en1,
    //input AXI-Stream to BRAM interface 100
    input s_axis_bram_100_aclk,
    input s_axis_bram_100_aresetn,
    input s_axis_bram_100_tlast,
    input s_axis_bram_100_tvalid,
    input [S_AXIS_BRAM_100_DMWIDTH/8-1:0] s_axis_bram_100_tkeep,
    input [S_AXIS_BRAM_100_DMWIDTH/8-1:0] s_axis_bram_100_tstrb,
    input [S_AXIS_BRAM_100_DMWIDTH-1:0] s_axis_bram_100_tdata,
    output s_axis_bram_100_tready,
    input [S_AXIS_BRAM_100_ADDR_WIDTH-1:0] ap_bram_iarg_100_addr0,
    input [S_AXIS_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_din0,
    output [S_AXIS_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_dout0,
    input ap_bram_iarg_100_clk0,
    input ap_bram_iarg_100_rst0,
    input [S_AXIS_BRAM_100_WIDTH/8-1:0] ap_bram_iarg_100_we0,
    input ap_bram_iarg_100_en0,
    input [S_AXIS_BRAM_100_ADDR_WIDTH-1:0] ap_bram_iarg_100_addr1,
    input [S_AXIS_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_din1,
    output [S_AXIS_BRAM_100_WIDTH-1:0] ap_bram_iarg_100_dout1,
    input ap_bram_iarg_100_clk1,
    input ap_bram_iarg_100_rst1,
    input [S_AXIS_BRAM_100_WIDTH/8-1:0] ap_bram_iarg_100_we1,
    input ap_bram_iarg_100_en1,
    //input AXI-Stream to BRAM interface 101
    input s_axis_bram_101_aclk,
    input s_axis_bram_101_aresetn,
    input s_axis_bram_101_tlast,
    input s_axis_bram_101_tvalid,
    input [S_AXIS_BRAM_101_DMWIDTH/8-1:0] s_axis_bram_101_tkeep,
    input [S_AXIS_BRAM_101_DMWIDTH/8-1:0] s_axis_bram_101_tstrb,
    input [S_AXIS_BRAM_101_DMWIDTH-1:0] s_axis_bram_101_tdata,
    output s_axis_bram_101_tready,
    input [S_AXIS_BRAM_101_ADDR_WIDTH-1:0] ap_bram_iarg_101_addr0,
    input [S_AXIS_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_din0,
    output [S_AXIS_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_dout0,
    input ap_bram_iarg_101_clk0,
    input ap_bram_iarg_101_rst0,
    input [S_AXIS_BRAM_101_WIDTH/8-1:0] ap_bram_iarg_101_we0,
    input ap_bram_iarg_101_en0,
    input [S_AXIS_BRAM_101_ADDR_WIDTH-1:0] ap_bram_iarg_101_addr1,
    input [S_AXIS_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_din1,
    output [S_AXIS_BRAM_101_WIDTH-1:0] ap_bram_iarg_101_dout1,
    input ap_bram_iarg_101_clk1,
    input ap_bram_iarg_101_rst1,
    input [S_AXIS_BRAM_101_WIDTH/8-1:0] ap_bram_iarg_101_we1,
    input ap_bram_iarg_101_en1,
    //input AXI-Stream to BRAM interface 102
    input s_axis_bram_102_aclk,
    input s_axis_bram_102_aresetn,
    input s_axis_bram_102_tlast,
    input s_axis_bram_102_tvalid,
    input [S_AXIS_BRAM_102_DMWIDTH/8-1:0] s_axis_bram_102_tkeep,
    input [S_AXIS_BRAM_102_DMWIDTH/8-1:0] s_axis_bram_102_tstrb,
    input [S_AXIS_BRAM_102_DMWIDTH-1:0] s_axis_bram_102_tdata,
    output s_axis_bram_102_tready,
    input [S_AXIS_BRAM_102_ADDR_WIDTH-1:0] ap_bram_iarg_102_addr0,
    input [S_AXIS_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_din0,
    output [S_AXIS_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_dout0,
    input ap_bram_iarg_102_clk0,
    input ap_bram_iarg_102_rst0,
    input [S_AXIS_BRAM_102_WIDTH/8-1:0] ap_bram_iarg_102_we0,
    input ap_bram_iarg_102_en0,
    input [S_AXIS_BRAM_102_ADDR_WIDTH-1:0] ap_bram_iarg_102_addr1,
    input [S_AXIS_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_din1,
    output [S_AXIS_BRAM_102_WIDTH-1:0] ap_bram_iarg_102_dout1,
    input ap_bram_iarg_102_clk1,
    input ap_bram_iarg_102_rst1,
    input [S_AXIS_BRAM_102_WIDTH/8-1:0] ap_bram_iarg_102_we1,
    input ap_bram_iarg_102_en1,
    //input AXI-Stream to BRAM interface 103
    input s_axis_bram_103_aclk,
    input s_axis_bram_103_aresetn,
    input s_axis_bram_103_tlast,
    input s_axis_bram_103_tvalid,
    input [S_AXIS_BRAM_103_DMWIDTH/8-1:0] s_axis_bram_103_tkeep,
    input [S_AXIS_BRAM_103_DMWIDTH/8-1:0] s_axis_bram_103_tstrb,
    input [S_AXIS_BRAM_103_DMWIDTH-1:0] s_axis_bram_103_tdata,
    output s_axis_bram_103_tready,
    input [S_AXIS_BRAM_103_ADDR_WIDTH-1:0] ap_bram_iarg_103_addr0,
    input [S_AXIS_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_din0,
    output [S_AXIS_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_dout0,
    input ap_bram_iarg_103_clk0,
    input ap_bram_iarg_103_rst0,
    input [S_AXIS_BRAM_103_WIDTH/8-1:0] ap_bram_iarg_103_we0,
    input ap_bram_iarg_103_en0,
    input [S_AXIS_BRAM_103_ADDR_WIDTH-1:0] ap_bram_iarg_103_addr1,
    input [S_AXIS_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_din1,
    output [S_AXIS_BRAM_103_WIDTH-1:0] ap_bram_iarg_103_dout1,
    input ap_bram_iarg_103_clk1,
    input ap_bram_iarg_103_rst1,
    input [S_AXIS_BRAM_103_WIDTH/8-1:0] ap_bram_iarg_103_we1,
    input ap_bram_iarg_103_en1,
    //input AXI-Stream to BRAM interface 104
    input s_axis_bram_104_aclk,
    input s_axis_bram_104_aresetn,
    input s_axis_bram_104_tlast,
    input s_axis_bram_104_tvalid,
    input [S_AXIS_BRAM_104_DMWIDTH/8-1:0] s_axis_bram_104_tkeep,
    input [S_AXIS_BRAM_104_DMWIDTH/8-1:0] s_axis_bram_104_tstrb,
    input [S_AXIS_BRAM_104_DMWIDTH-1:0] s_axis_bram_104_tdata,
    output s_axis_bram_104_tready,
    input [S_AXIS_BRAM_104_ADDR_WIDTH-1:0] ap_bram_iarg_104_addr0,
    input [S_AXIS_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_din0,
    output [S_AXIS_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_dout0,
    input ap_bram_iarg_104_clk0,
    input ap_bram_iarg_104_rst0,
    input [S_AXIS_BRAM_104_WIDTH/8-1:0] ap_bram_iarg_104_we0,
    input ap_bram_iarg_104_en0,
    input [S_AXIS_BRAM_104_ADDR_WIDTH-1:0] ap_bram_iarg_104_addr1,
    input [S_AXIS_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_din1,
    output [S_AXIS_BRAM_104_WIDTH-1:0] ap_bram_iarg_104_dout1,
    input ap_bram_iarg_104_clk1,
    input ap_bram_iarg_104_rst1,
    input [S_AXIS_BRAM_104_WIDTH/8-1:0] ap_bram_iarg_104_we1,
    input ap_bram_iarg_104_en1,
    //input AXI-Stream to BRAM interface 105
    input s_axis_bram_105_aclk,
    input s_axis_bram_105_aresetn,
    input s_axis_bram_105_tlast,
    input s_axis_bram_105_tvalid,
    input [S_AXIS_BRAM_105_DMWIDTH/8-1:0] s_axis_bram_105_tkeep,
    input [S_AXIS_BRAM_105_DMWIDTH/8-1:0] s_axis_bram_105_tstrb,
    input [S_AXIS_BRAM_105_DMWIDTH-1:0] s_axis_bram_105_tdata,
    output s_axis_bram_105_tready,
    input [S_AXIS_BRAM_105_ADDR_WIDTH-1:0] ap_bram_iarg_105_addr0,
    input [S_AXIS_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_din0,
    output [S_AXIS_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_dout0,
    input ap_bram_iarg_105_clk0,
    input ap_bram_iarg_105_rst0,
    input [S_AXIS_BRAM_105_WIDTH/8-1:0] ap_bram_iarg_105_we0,
    input ap_bram_iarg_105_en0,
    input [S_AXIS_BRAM_105_ADDR_WIDTH-1:0] ap_bram_iarg_105_addr1,
    input [S_AXIS_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_din1,
    output [S_AXIS_BRAM_105_WIDTH-1:0] ap_bram_iarg_105_dout1,
    input ap_bram_iarg_105_clk1,
    input ap_bram_iarg_105_rst1,
    input [S_AXIS_BRAM_105_WIDTH/8-1:0] ap_bram_iarg_105_we1,
    input ap_bram_iarg_105_en1,
    //input AXI-Stream to BRAM interface 106
    input s_axis_bram_106_aclk,
    input s_axis_bram_106_aresetn,
    input s_axis_bram_106_tlast,
    input s_axis_bram_106_tvalid,
    input [S_AXIS_BRAM_106_DMWIDTH/8-1:0] s_axis_bram_106_tkeep,
    input [S_AXIS_BRAM_106_DMWIDTH/8-1:0] s_axis_bram_106_tstrb,
    input [S_AXIS_BRAM_106_DMWIDTH-1:0] s_axis_bram_106_tdata,
    output s_axis_bram_106_tready,
    input [S_AXIS_BRAM_106_ADDR_WIDTH-1:0] ap_bram_iarg_106_addr0,
    input [S_AXIS_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_din0,
    output [S_AXIS_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_dout0,
    input ap_bram_iarg_106_clk0,
    input ap_bram_iarg_106_rst0,
    input [S_AXIS_BRAM_106_WIDTH/8-1:0] ap_bram_iarg_106_we0,
    input ap_bram_iarg_106_en0,
    input [S_AXIS_BRAM_106_ADDR_WIDTH-1:0] ap_bram_iarg_106_addr1,
    input [S_AXIS_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_din1,
    output [S_AXIS_BRAM_106_WIDTH-1:0] ap_bram_iarg_106_dout1,
    input ap_bram_iarg_106_clk1,
    input ap_bram_iarg_106_rst1,
    input [S_AXIS_BRAM_106_WIDTH/8-1:0] ap_bram_iarg_106_we1,
    input ap_bram_iarg_106_en1,
    //input AXI-Stream to BRAM interface 107
    input s_axis_bram_107_aclk,
    input s_axis_bram_107_aresetn,
    input s_axis_bram_107_tlast,
    input s_axis_bram_107_tvalid,
    input [S_AXIS_BRAM_107_DMWIDTH/8-1:0] s_axis_bram_107_tkeep,
    input [S_AXIS_BRAM_107_DMWIDTH/8-1:0] s_axis_bram_107_tstrb,
    input [S_AXIS_BRAM_107_DMWIDTH-1:0] s_axis_bram_107_tdata,
    output s_axis_bram_107_tready,
    input [S_AXIS_BRAM_107_ADDR_WIDTH-1:0] ap_bram_iarg_107_addr0,
    input [S_AXIS_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_din0,
    output [S_AXIS_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_dout0,
    input ap_bram_iarg_107_clk0,
    input ap_bram_iarg_107_rst0,
    input [S_AXIS_BRAM_107_WIDTH/8-1:0] ap_bram_iarg_107_we0,
    input ap_bram_iarg_107_en0,
    input [S_AXIS_BRAM_107_ADDR_WIDTH-1:0] ap_bram_iarg_107_addr1,
    input [S_AXIS_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_din1,
    output [S_AXIS_BRAM_107_WIDTH-1:0] ap_bram_iarg_107_dout1,
    input ap_bram_iarg_107_clk1,
    input ap_bram_iarg_107_rst1,
    input [S_AXIS_BRAM_107_WIDTH/8-1:0] ap_bram_iarg_107_we1,
    input ap_bram_iarg_107_en1,
    //input AXI-Stream to BRAM interface 108
    input s_axis_bram_108_aclk,
    input s_axis_bram_108_aresetn,
    input s_axis_bram_108_tlast,
    input s_axis_bram_108_tvalid,
    input [S_AXIS_BRAM_108_DMWIDTH/8-1:0] s_axis_bram_108_tkeep,
    input [S_AXIS_BRAM_108_DMWIDTH/8-1:0] s_axis_bram_108_tstrb,
    input [S_AXIS_BRAM_108_DMWIDTH-1:0] s_axis_bram_108_tdata,
    output s_axis_bram_108_tready,
    input [S_AXIS_BRAM_108_ADDR_WIDTH-1:0] ap_bram_iarg_108_addr0,
    input [S_AXIS_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_din0,
    output [S_AXIS_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_dout0,
    input ap_bram_iarg_108_clk0,
    input ap_bram_iarg_108_rst0,
    input [S_AXIS_BRAM_108_WIDTH/8-1:0] ap_bram_iarg_108_we0,
    input ap_bram_iarg_108_en0,
    input [S_AXIS_BRAM_108_ADDR_WIDTH-1:0] ap_bram_iarg_108_addr1,
    input [S_AXIS_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_din1,
    output [S_AXIS_BRAM_108_WIDTH-1:0] ap_bram_iarg_108_dout1,
    input ap_bram_iarg_108_clk1,
    input ap_bram_iarg_108_rst1,
    input [S_AXIS_BRAM_108_WIDTH/8-1:0] ap_bram_iarg_108_we1,
    input ap_bram_iarg_108_en1,
    //input AXI-Stream to BRAM interface 109
    input s_axis_bram_109_aclk,
    input s_axis_bram_109_aresetn,
    input s_axis_bram_109_tlast,
    input s_axis_bram_109_tvalid,
    input [S_AXIS_BRAM_109_DMWIDTH/8-1:0] s_axis_bram_109_tkeep,
    input [S_AXIS_BRAM_109_DMWIDTH/8-1:0] s_axis_bram_109_tstrb,
    input [S_AXIS_BRAM_109_DMWIDTH-1:0] s_axis_bram_109_tdata,
    output s_axis_bram_109_tready,
    input [S_AXIS_BRAM_109_ADDR_WIDTH-1:0] ap_bram_iarg_109_addr0,
    input [S_AXIS_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_din0,
    output [S_AXIS_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_dout0,
    input ap_bram_iarg_109_clk0,
    input ap_bram_iarg_109_rst0,
    input [S_AXIS_BRAM_109_WIDTH/8-1:0] ap_bram_iarg_109_we0,
    input ap_bram_iarg_109_en0,
    input [S_AXIS_BRAM_109_ADDR_WIDTH-1:0] ap_bram_iarg_109_addr1,
    input [S_AXIS_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_din1,
    output [S_AXIS_BRAM_109_WIDTH-1:0] ap_bram_iarg_109_dout1,
    input ap_bram_iarg_109_clk1,
    input ap_bram_iarg_109_rst1,
    input [S_AXIS_BRAM_109_WIDTH/8-1:0] ap_bram_iarg_109_we1,
    input ap_bram_iarg_109_en1,
    //input AXI-Stream to BRAM interface 110
    input s_axis_bram_110_aclk,
    input s_axis_bram_110_aresetn,
    input s_axis_bram_110_tlast,
    input s_axis_bram_110_tvalid,
    input [S_AXIS_BRAM_110_DMWIDTH/8-1:0] s_axis_bram_110_tkeep,
    input [S_AXIS_BRAM_110_DMWIDTH/8-1:0] s_axis_bram_110_tstrb,
    input [S_AXIS_BRAM_110_DMWIDTH-1:0] s_axis_bram_110_tdata,
    output s_axis_bram_110_tready,
    input [S_AXIS_BRAM_110_ADDR_WIDTH-1:0] ap_bram_iarg_110_addr0,
    input [S_AXIS_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_din0,
    output [S_AXIS_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_dout0,
    input ap_bram_iarg_110_clk0,
    input ap_bram_iarg_110_rst0,
    input [S_AXIS_BRAM_110_WIDTH/8-1:0] ap_bram_iarg_110_we0,
    input ap_bram_iarg_110_en0,
    input [S_AXIS_BRAM_110_ADDR_WIDTH-1:0] ap_bram_iarg_110_addr1,
    input [S_AXIS_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_din1,
    output [S_AXIS_BRAM_110_WIDTH-1:0] ap_bram_iarg_110_dout1,
    input ap_bram_iarg_110_clk1,
    input ap_bram_iarg_110_rst1,
    input [S_AXIS_BRAM_110_WIDTH/8-1:0] ap_bram_iarg_110_we1,
    input ap_bram_iarg_110_en1,
    //input AXI-Stream to BRAM interface 111
    input s_axis_bram_111_aclk,
    input s_axis_bram_111_aresetn,
    input s_axis_bram_111_tlast,
    input s_axis_bram_111_tvalid,
    input [S_AXIS_BRAM_111_DMWIDTH/8-1:0] s_axis_bram_111_tkeep,
    input [S_AXIS_BRAM_111_DMWIDTH/8-1:0] s_axis_bram_111_tstrb,
    input [S_AXIS_BRAM_111_DMWIDTH-1:0] s_axis_bram_111_tdata,
    output s_axis_bram_111_tready,
    input [S_AXIS_BRAM_111_ADDR_WIDTH-1:0] ap_bram_iarg_111_addr0,
    input [S_AXIS_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_din0,
    output [S_AXIS_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_dout0,
    input ap_bram_iarg_111_clk0,
    input ap_bram_iarg_111_rst0,
    input [S_AXIS_BRAM_111_WIDTH/8-1:0] ap_bram_iarg_111_we0,
    input ap_bram_iarg_111_en0,
    input [S_AXIS_BRAM_111_ADDR_WIDTH-1:0] ap_bram_iarg_111_addr1,
    input [S_AXIS_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_din1,
    output [S_AXIS_BRAM_111_WIDTH-1:0] ap_bram_iarg_111_dout1,
    input ap_bram_iarg_111_clk1,
    input ap_bram_iarg_111_rst1,
    input [S_AXIS_BRAM_111_WIDTH/8-1:0] ap_bram_iarg_111_we1,
    input ap_bram_iarg_111_en1,
    //input AXI-Stream to BRAM interface 112
    input s_axis_bram_112_aclk,
    input s_axis_bram_112_aresetn,
    input s_axis_bram_112_tlast,
    input s_axis_bram_112_tvalid,
    input [S_AXIS_BRAM_112_DMWIDTH/8-1:0] s_axis_bram_112_tkeep,
    input [S_AXIS_BRAM_112_DMWIDTH/8-1:0] s_axis_bram_112_tstrb,
    input [S_AXIS_BRAM_112_DMWIDTH-1:0] s_axis_bram_112_tdata,
    output s_axis_bram_112_tready,
    input [S_AXIS_BRAM_112_ADDR_WIDTH-1:0] ap_bram_iarg_112_addr0,
    input [S_AXIS_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_din0,
    output [S_AXIS_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_dout0,
    input ap_bram_iarg_112_clk0,
    input ap_bram_iarg_112_rst0,
    input [S_AXIS_BRAM_112_WIDTH/8-1:0] ap_bram_iarg_112_we0,
    input ap_bram_iarg_112_en0,
    input [S_AXIS_BRAM_112_ADDR_WIDTH-1:0] ap_bram_iarg_112_addr1,
    input [S_AXIS_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_din1,
    output [S_AXIS_BRAM_112_WIDTH-1:0] ap_bram_iarg_112_dout1,
    input ap_bram_iarg_112_clk1,
    input ap_bram_iarg_112_rst1,
    input [S_AXIS_BRAM_112_WIDTH/8-1:0] ap_bram_iarg_112_we1,
    input ap_bram_iarg_112_en1,
    //input AXI-Stream to BRAM interface 113
    input s_axis_bram_113_aclk,
    input s_axis_bram_113_aresetn,
    input s_axis_bram_113_tlast,
    input s_axis_bram_113_tvalid,
    input [S_AXIS_BRAM_113_DMWIDTH/8-1:0] s_axis_bram_113_tkeep,
    input [S_AXIS_BRAM_113_DMWIDTH/8-1:0] s_axis_bram_113_tstrb,
    input [S_AXIS_BRAM_113_DMWIDTH-1:0] s_axis_bram_113_tdata,
    output s_axis_bram_113_tready,
    input [S_AXIS_BRAM_113_ADDR_WIDTH-1:0] ap_bram_iarg_113_addr0,
    input [S_AXIS_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_din0,
    output [S_AXIS_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_dout0,
    input ap_bram_iarg_113_clk0,
    input ap_bram_iarg_113_rst0,
    input [S_AXIS_BRAM_113_WIDTH/8-1:0] ap_bram_iarg_113_we0,
    input ap_bram_iarg_113_en0,
    input [S_AXIS_BRAM_113_ADDR_WIDTH-1:0] ap_bram_iarg_113_addr1,
    input [S_AXIS_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_din1,
    output [S_AXIS_BRAM_113_WIDTH-1:0] ap_bram_iarg_113_dout1,
    input ap_bram_iarg_113_clk1,
    input ap_bram_iarg_113_rst1,
    input [S_AXIS_BRAM_113_WIDTH/8-1:0] ap_bram_iarg_113_we1,
    input ap_bram_iarg_113_en1,
    //input AXI-Stream to BRAM interface 114
    input s_axis_bram_114_aclk,
    input s_axis_bram_114_aresetn,
    input s_axis_bram_114_tlast,
    input s_axis_bram_114_tvalid,
    input [S_AXIS_BRAM_114_DMWIDTH/8-1:0] s_axis_bram_114_tkeep,
    input [S_AXIS_BRAM_114_DMWIDTH/8-1:0] s_axis_bram_114_tstrb,
    input [S_AXIS_BRAM_114_DMWIDTH-1:0] s_axis_bram_114_tdata,
    output s_axis_bram_114_tready,
    input [S_AXIS_BRAM_114_ADDR_WIDTH-1:0] ap_bram_iarg_114_addr0,
    input [S_AXIS_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_din0,
    output [S_AXIS_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_dout0,
    input ap_bram_iarg_114_clk0,
    input ap_bram_iarg_114_rst0,
    input [S_AXIS_BRAM_114_WIDTH/8-1:0] ap_bram_iarg_114_we0,
    input ap_bram_iarg_114_en0,
    input [S_AXIS_BRAM_114_ADDR_WIDTH-1:0] ap_bram_iarg_114_addr1,
    input [S_AXIS_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_din1,
    output [S_AXIS_BRAM_114_WIDTH-1:0] ap_bram_iarg_114_dout1,
    input ap_bram_iarg_114_clk1,
    input ap_bram_iarg_114_rst1,
    input [S_AXIS_BRAM_114_WIDTH/8-1:0] ap_bram_iarg_114_we1,
    input ap_bram_iarg_114_en1,
    //input AXI-Stream to BRAM interface 115
    input s_axis_bram_115_aclk,
    input s_axis_bram_115_aresetn,
    input s_axis_bram_115_tlast,
    input s_axis_bram_115_tvalid,
    input [S_AXIS_BRAM_115_DMWIDTH/8-1:0] s_axis_bram_115_tkeep,
    input [S_AXIS_BRAM_115_DMWIDTH/8-1:0] s_axis_bram_115_tstrb,
    input [S_AXIS_BRAM_115_DMWIDTH-1:0] s_axis_bram_115_tdata,
    output s_axis_bram_115_tready,
    input [S_AXIS_BRAM_115_ADDR_WIDTH-1:0] ap_bram_iarg_115_addr0,
    input [S_AXIS_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_din0,
    output [S_AXIS_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_dout0,
    input ap_bram_iarg_115_clk0,
    input ap_bram_iarg_115_rst0,
    input [S_AXIS_BRAM_115_WIDTH/8-1:0] ap_bram_iarg_115_we0,
    input ap_bram_iarg_115_en0,
    input [S_AXIS_BRAM_115_ADDR_WIDTH-1:0] ap_bram_iarg_115_addr1,
    input [S_AXIS_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_din1,
    output [S_AXIS_BRAM_115_WIDTH-1:0] ap_bram_iarg_115_dout1,
    input ap_bram_iarg_115_clk1,
    input ap_bram_iarg_115_rst1,
    input [S_AXIS_BRAM_115_WIDTH/8-1:0] ap_bram_iarg_115_we1,
    input ap_bram_iarg_115_en1,
    //input AXI-Stream to BRAM interface 116
    input s_axis_bram_116_aclk,
    input s_axis_bram_116_aresetn,
    input s_axis_bram_116_tlast,
    input s_axis_bram_116_tvalid,
    input [S_AXIS_BRAM_116_DMWIDTH/8-1:0] s_axis_bram_116_tkeep,
    input [S_AXIS_BRAM_116_DMWIDTH/8-1:0] s_axis_bram_116_tstrb,
    input [S_AXIS_BRAM_116_DMWIDTH-1:0] s_axis_bram_116_tdata,
    output s_axis_bram_116_tready,
    input [S_AXIS_BRAM_116_ADDR_WIDTH-1:0] ap_bram_iarg_116_addr0,
    input [S_AXIS_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_din0,
    output [S_AXIS_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_dout0,
    input ap_bram_iarg_116_clk0,
    input ap_bram_iarg_116_rst0,
    input [S_AXIS_BRAM_116_WIDTH/8-1:0] ap_bram_iarg_116_we0,
    input ap_bram_iarg_116_en0,
    input [S_AXIS_BRAM_116_ADDR_WIDTH-1:0] ap_bram_iarg_116_addr1,
    input [S_AXIS_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_din1,
    output [S_AXIS_BRAM_116_WIDTH-1:0] ap_bram_iarg_116_dout1,
    input ap_bram_iarg_116_clk1,
    input ap_bram_iarg_116_rst1,
    input [S_AXIS_BRAM_116_WIDTH/8-1:0] ap_bram_iarg_116_we1,
    input ap_bram_iarg_116_en1,
    //input AXI-Stream to BRAM interface 117
    input s_axis_bram_117_aclk,
    input s_axis_bram_117_aresetn,
    input s_axis_bram_117_tlast,
    input s_axis_bram_117_tvalid,
    input [S_AXIS_BRAM_117_DMWIDTH/8-1:0] s_axis_bram_117_tkeep,
    input [S_AXIS_BRAM_117_DMWIDTH/8-1:0] s_axis_bram_117_tstrb,
    input [S_AXIS_BRAM_117_DMWIDTH-1:0] s_axis_bram_117_tdata,
    output s_axis_bram_117_tready,
    input [S_AXIS_BRAM_117_ADDR_WIDTH-1:0] ap_bram_iarg_117_addr0,
    input [S_AXIS_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_din0,
    output [S_AXIS_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_dout0,
    input ap_bram_iarg_117_clk0,
    input ap_bram_iarg_117_rst0,
    input [S_AXIS_BRAM_117_WIDTH/8-1:0] ap_bram_iarg_117_we0,
    input ap_bram_iarg_117_en0,
    input [S_AXIS_BRAM_117_ADDR_WIDTH-1:0] ap_bram_iarg_117_addr1,
    input [S_AXIS_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_din1,
    output [S_AXIS_BRAM_117_WIDTH-1:0] ap_bram_iarg_117_dout1,
    input ap_bram_iarg_117_clk1,
    input ap_bram_iarg_117_rst1,
    input [S_AXIS_BRAM_117_WIDTH/8-1:0] ap_bram_iarg_117_we1,
    input ap_bram_iarg_117_en1,
    //input AXI-Stream to BRAM interface 118
    input s_axis_bram_118_aclk,
    input s_axis_bram_118_aresetn,
    input s_axis_bram_118_tlast,
    input s_axis_bram_118_tvalid,
    input [S_AXIS_BRAM_118_DMWIDTH/8-1:0] s_axis_bram_118_tkeep,
    input [S_AXIS_BRAM_118_DMWIDTH/8-1:0] s_axis_bram_118_tstrb,
    input [S_AXIS_BRAM_118_DMWIDTH-1:0] s_axis_bram_118_tdata,
    output s_axis_bram_118_tready,
    input [S_AXIS_BRAM_118_ADDR_WIDTH-1:0] ap_bram_iarg_118_addr0,
    input [S_AXIS_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_din0,
    output [S_AXIS_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_dout0,
    input ap_bram_iarg_118_clk0,
    input ap_bram_iarg_118_rst0,
    input [S_AXIS_BRAM_118_WIDTH/8-1:0] ap_bram_iarg_118_we0,
    input ap_bram_iarg_118_en0,
    input [S_AXIS_BRAM_118_ADDR_WIDTH-1:0] ap_bram_iarg_118_addr1,
    input [S_AXIS_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_din1,
    output [S_AXIS_BRAM_118_WIDTH-1:0] ap_bram_iarg_118_dout1,
    input ap_bram_iarg_118_clk1,
    input ap_bram_iarg_118_rst1,
    input [S_AXIS_BRAM_118_WIDTH/8-1:0] ap_bram_iarg_118_we1,
    input ap_bram_iarg_118_en1,
    //input AXI-Stream to BRAM interface 119
    input s_axis_bram_119_aclk,
    input s_axis_bram_119_aresetn,
    input s_axis_bram_119_tlast,
    input s_axis_bram_119_tvalid,
    input [S_AXIS_BRAM_119_DMWIDTH/8-1:0] s_axis_bram_119_tkeep,
    input [S_AXIS_BRAM_119_DMWIDTH/8-1:0] s_axis_bram_119_tstrb,
    input [S_AXIS_BRAM_119_DMWIDTH-1:0] s_axis_bram_119_tdata,
    output s_axis_bram_119_tready,
    input [S_AXIS_BRAM_119_ADDR_WIDTH-1:0] ap_bram_iarg_119_addr0,
    input [S_AXIS_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_din0,
    output [S_AXIS_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_dout0,
    input ap_bram_iarg_119_clk0,
    input ap_bram_iarg_119_rst0,
    input [S_AXIS_BRAM_119_WIDTH/8-1:0] ap_bram_iarg_119_we0,
    input ap_bram_iarg_119_en0,
    input [S_AXIS_BRAM_119_ADDR_WIDTH-1:0] ap_bram_iarg_119_addr1,
    input [S_AXIS_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_din1,
    output [S_AXIS_BRAM_119_WIDTH-1:0] ap_bram_iarg_119_dout1,
    input ap_bram_iarg_119_clk1,
    input ap_bram_iarg_119_rst1,
    input [S_AXIS_BRAM_119_WIDTH/8-1:0] ap_bram_iarg_119_we1,
    input ap_bram_iarg_119_en1,
    //input AXI-Stream to BRAM interface 120
    input s_axis_bram_120_aclk,
    input s_axis_bram_120_aresetn,
    input s_axis_bram_120_tlast,
    input s_axis_bram_120_tvalid,
    input [S_AXIS_BRAM_120_DMWIDTH/8-1:0] s_axis_bram_120_tkeep,
    input [S_AXIS_BRAM_120_DMWIDTH/8-1:0] s_axis_bram_120_tstrb,
    input [S_AXIS_BRAM_120_DMWIDTH-1:0] s_axis_bram_120_tdata,
    output s_axis_bram_120_tready,
    input [S_AXIS_BRAM_120_ADDR_WIDTH-1:0] ap_bram_iarg_120_addr0,
    input [S_AXIS_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_din0,
    output [S_AXIS_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_dout0,
    input ap_bram_iarg_120_clk0,
    input ap_bram_iarg_120_rst0,
    input [S_AXIS_BRAM_120_WIDTH/8-1:0] ap_bram_iarg_120_we0,
    input ap_bram_iarg_120_en0,
    input [S_AXIS_BRAM_120_ADDR_WIDTH-1:0] ap_bram_iarg_120_addr1,
    input [S_AXIS_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_din1,
    output [S_AXIS_BRAM_120_WIDTH-1:0] ap_bram_iarg_120_dout1,
    input ap_bram_iarg_120_clk1,
    input ap_bram_iarg_120_rst1,
    input [S_AXIS_BRAM_120_WIDTH/8-1:0] ap_bram_iarg_120_we1,
    input ap_bram_iarg_120_en1,
    //input AXI-Stream to BRAM interface 121
    input s_axis_bram_121_aclk,
    input s_axis_bram_121_aresetn,
    input s_axis_bram_121_tlast,
    input s_axis_bram_121_tvalid,
    input [S_AXIS_BRAM_121_DMWIDTH/8-1:0] s_axis_bram_121_tkeep,
    input [S_AXIS_BRAM_121_DMWIDTH/8-1:0] s_axis_bram_121_tstrb,
    input [S_AXIS_BRAM_121_DMWIDTH-1:0] s_axis_bram_121_tdata,
    output s_axis_bram_121_tready,
    input [S_AXIS_BRAM_121_ADDR_WIDTH-1:0] ap_bram_iarg_121_addr0,
    input [S_AXIS_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_din0,
    output [S_AXIS_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_dout0,
    input ap_bram_iarg_121_clk0,
    input ap_bram_iarg_121_rst0,
    input [S_AXIS_BRAM_121_WIDTH/8-1:0] ap_bram_iarg_121_we0,
    input ap_bram_iarg_121_en0,
    input [S_AXIS_BRAM_121_ADDR_WIDTH-1:0] ap_bram_iarg_121_addr1,
    input [S_AXIS_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_din1,
    output [S_AXIS_BRAM_121_WIDTH-1:0] ap_bram_iarg_121_dout1,
    input ap_bram_iarg_121_clk1,
    input ap_bram_iarg_121_rst1,
    input [S_AXIS_BRAM_121_WIDTH/8-1:0] ap_bram_iarg_121_we1,
    input ap_bram_iarg_121_en1,
    //input AXI-Stream to BRAM interface 122
    input s_axis_bram_122_aclk,
    input s_axis_bram_122_aresetn,
    input s_axis_bram_122_tlast,
    input s_axis_bram_122_tvalid,
    input [S_AXIS_BRAM_122_DMWIDTH/8-1:0] s_axis_bram_122_tkeep,
    input [S_AXIS_BRAM_122_DMWIDTH/8-1:0] s_axis_bram_122_tstrb,
    input [S_AXIS_BRAM_122_DMWIDTH-1:0] s_axis_bram_122_tdata,
    output s_axis_bram_122_tready,
    input [S_AXIS_BRAM_122_ADDR_WIDTH-1:0] ap_bram_iarg_122_addr0,
    input [S_AXIS_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_din0,
    output [S_AXIS_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_dout0,
    input ap_bram_iarg_122_clk0,
    input ap_bram_iarg_122_rst0,
    input [S_AXIS_BRAM_122_WIDTH/8-1:0] ap_bram_iarg_122_we0,
    input ap_bram_iarg_122_en0,
    input [S_AXIS_BRAM_122_ADDR_WIDTH-1:0] ap_bram_iarg_122_addr1,
    input [S_AXIS_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_din1,
    output [S_AXIS_BRAM_122_WIDTH-1:0] ap_bram_iarg_122_dout1,
    input ap_bram_iarg_122_clk1,
    input ap_bram_iarg_122_rst1,
    input [S_AXIS_BRAM_122_WIDTH/8-1:0] ap_bram_iarg_122_we1,
    input ap_bram_iarg_122_en1,
    //input AXI-Stream to BRAM interface 123
    input s_axis_bram_123_aclk,
    input s_axis_bram_123_aresetn,
    input s_axis_bram_123_tlast,
    input s_axis_bram_123_tvalid,
    input [S_AXIS_BRAM_123_DMWIDTH/8-1:0] s_axis_bram_123_tkeep,
    input [S_AXIS_BRAM_123_DMWIDTH/8-1:0] s_axis_bram_123_tstrb,
    input [S_AXIS_BRAM_123_DMWIDTH-1:0] s_axis_bram_123_tdata,
    output s_axis_bram_123_tready,
    input [S_AXIS_BRAM_123_ADDR_WIDTH-1:0] ap_bram_iarg_123_addr0,
    input [S_AXIS_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_din0,
    output [S_AXIS_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_dout0,
    input ap_bram_iarg_123_clk0,
    input ap_bram_iarg_123_rst0,
    input [S_AXIS_BRAM_123_WIDTH/8-1:0] ap_bram_iarg_123_we0,
    input ap_bram_iarg_123_en0,
    input [S_AXIS_BRAM_123_ADDR_WIDTH-1:0] ap_bram_iarg_123_addr1,
    input [S_AXIS_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_din1,
    output [S_AXIS_BRAM_123_WIDTH-1:0] ap_bram_iarg_123_dout1,
    input ap_bram_iarg_123_clk1,
    input ap_bram_iarg_123_rst1,
    input [S_AXIS_BRAM_123_WIDTH/8-1:0] ap_bram_iarg_123_we1,
    input ap_bram_iarg_123_en1,
    //input AXI-Stream to BRAM interface 124
    input s_axis_bram_124_aclk,
    input s_axis_bram_124_aresetn,
    input s_axis_bram_124_tlast,
    input s_axis_bram_124_tvalid,
    input [S_AXIS_BRAM_124_DMWIDTH/8-1:0] s_axis_bram_124_tkeep,
    input [S_AXIS_BRAM_124_DMWIDTH/8-1:0] s_axis_bram_124_tstrb,
    input [S_AXIS_BRAM_124_DMWIDTH-1:0] s_axis_bram_124_tdata,
    output s_axis_bram_124_tready,
    input [S_AXIS_BRAM_124_ADDR_WIDTH-1:0] ap_bram_iarg_124_addr0,
    input [S_AXIS_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_din0,
    output [S_AXIS_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_dout0,
    input ap_bram_iarg_124_clk0,
    input ap_bram_iarg_124_rst0,
    input [S_AXIS_BRAM_124_WIDTH/8-1:0] ap_bram_iarg_124_we0,
    input ap_bram_iarg_124_en0,
    input [S_AXIS_BRAM_124_ADDR_WIDTH-1:0] ap_bram_iarg_124_addr1,
    input [S_AXIS_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_din1,
    output [S_AXIS_BRAM_124_WIDTH-1:0] ap_bram_iarg_124_dout1,
    input ap_bram_iarg_124_clk1,
    input ap_bram_iarg_124_rst1,
    input [S_AXIS_BRAM_124_WIDTH/8-1:0] ap_bram_iarg_124_we1,
    input ap_bram_iarg_124_en1,
    //input AXI-Stream to BRAM interface 125
    input s_axis_bram_125_aclk,
    input s_axis_bram_125_aresetn,
    input s_axis_bram_125_tlast,
    input s_axis_bram_125_tvalid,
    input [S_AXIS_BRAM_125_DMWIDTH/8-1:0] s_axis_bram_125_tkeep,
    input [S_AXIS_BRAM_125_DMWIDTH/8-1:0] s_axis_bram_125_tstrb,
    input [S_AXIS_BRAM_125_DMWIDTH-1:0] s_axis_bram_125_tdata,
    output s_axis_bram_125_tready,
    input [S_AXIS_BRAM_125_ADDR_WIDTH-1:0] ap_bram_iarg_125_addr0,
    input [S_AXIS_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_din0,
    output [S_AXIS_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_dout0,
    input ap_bram_iarg_125_clk0,
    input ap_bram_iarg_125_rst0,
    input [S_AXIS_BRAM_125_WIDTH/8-1:0] ap_bram_iarg_125_we0,
    input ap_bram_iarg_125_en0,
    input [S_AXIS_BRAM_125_ADDR_WIDTH-1:0] ap_bram_iarg_125_addr1,
    input [S_AXIS_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_din1,
    output [S_AXIS_BRAM_125_WIDTH-1:0] ap_bram_iarg_125_dout1,
    input ap_bram_iarg_125_clk1,
    input ap_bram_iarg_125_rst1,
    input [S_AXIS_BRAM_125_WIDTH/8-1:0] ap_bram_iarg_125_we1,
    input ap_bram_iarg_125_en1,
    //input AXI-Stream to BRAM interface 126
    input s_axis_bram_126_aclk,
    input s_axis_bram_126_aresetn,
    input s_axis_bram_126_tlast,
    input s_axis_bram_126_tvalid,
    input [S_AXIS_BRAM_126_DMWIDTH/8-1:0] s_axis_bram_126_tkeep,
    input [S_AXIS_BRAM_126_DMWIDTH/8-1:0] s_axis_bram_126_tstrb,
    input [S_AXIS_BRAM_126_DMWIDTH-1:0] s_axis_bram_126_tdata,
    output s_axis_bram_126_tready,
    input [S_AXIS_BRAM_126_ADDR_WIDTH-1:0] ap_bram_iarg_126_addr0,
    input [S_AXIS_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_din0,
    output [S_AXIS_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_dout0,
    input ap_bram_iarg_126_clk0,
    input ap_bram_iarg_126_rst0,
    input [S_AXIS_BRAM_126_WIDTH/8-1:0] ap_bram_iarg_126_we0,
    input ap_bram_iarg_126_en0,
    input [S_AXIS_BRAM_126_ADDR_WIDTH-1:0] ap_bram_iarg_126_addr1,
    input [S_AXIS_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_din1,
    output [S_AXIS_BRAM_126_WIDTH-1:0] ap_bram_iarg_126_dout1,
    input ap_bram_iarg_126_clk1,
    input ap_bram_iarg_126_rst1,
    input [S_AXIS_BRAM_126_WIDTH/8-1:0] ap_bram_iarg_126_we1,
    input ap_bram_iarg_126_en1,
    //input AXI-Stream to BRAM interface 127
    input s_axis_bram_127_aclk,
    input s_axis_bram_127_aresetn,
    input s_axis_bram_127_tlast,
    input s_axis_bram_127_tvalid,
    input [S_AXIS_BRAM_127_DMWIDTH/8-1:0] s_axis_bram_127_tkeep,
    input [S_AXIS_BRAM_127_DMWIDTH/8-1:0] s_axis_bram_127_tstrb,
    input [S_AXIS_BRAM_127_DMWIDTH-1:0] s_axis_bram_127_tdata,
    output s_axis_bram_127_tready,
    input [S_AXIS_BRAM_127_ADDR_WIDTH-1:0] ap_bram_iarg_127_addr0,
    input [S_AXIS_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_din0,
    output [S_AXIS_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_dout0,
    input ap_bram_iarg_127_clk0,
    input ap_bram_iarg_127_rst0,
    input [S_AXIS_BRAM_127_WIDTH/8-1:0] ap_bram_iarg_127_we0,
    input ap_bram_iarg_127_en0,
    input [S_AXIS_BRAM_127_ADDR_WIDTH-1:0] ap_bram_iarg_127_addr1,
    input [S_AXIS_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_din1,
    output [S_AXIS_BRAM_127_WIDTH-1:0] ap_bram_iarg_127_dout1,
    input ap_bram_iarg_127_clk1,
    input ap_bram_iarg_127_rst1,
    input [S_AXIS_BRAM_127_WIDTH/8-1:0] ap_bram_iarg_127_we1,
    input ap_bram_iarg_127_en1,
    //-----------------------------------------------------------
    //in-out BRAM AXI-Stream output interface 0
    input m_axis_bramio_0_aclk,
    input m_axis_bramio_0_aresetn,
    output m_axis_bramio_0_tlast,
    output m_axis_bramio_0_tvalid,
    output [M_AXIS_BRAMIO_0_DMWIDTH/8-1:0] m_axis_bramio_0_tkeep,
    output [M_AXIS_BRAMIO_0_DMWIDTH/8-1:0] m_axis_bramio_0_tstrb,
    output [M_AXIS_BRAMIO_0_DMWIDTH-1:0] m_axis_bramio_0_tdata,
    input m_axis_bramio_0_tready,
    //in-out BRAM AXI-Stream output interface 1
    input m_axis_bramio_1_aclk,
    input m_axis_bramio_1_aresetn,
    output m_axis_bramio_1_tlast,
    output m_axis_bramio_1_tvalid,
    output [M_AXIS_BRAMIO_1_DMWIDTH/8-1:0] m_axis_bramio_1_tkeep,
    output [M_AXIS_BRAMIO_1_DMWIDTH/8-1:0] m_axis_bramio_1_tstrb,
    output [M_AXIS_BRAMIO_1_DMWIDTH-1:0] m_axis_bramio_1_tdata,
    input m_axis_bramio_1_tready,
    //in-out BRAM AXI-Stream output interface 2
    input m_axis_bramio_2_aclk,
    input m_axis_bramio_2_aresetn,
    output m_axis_bramio_2_tlast,
    output m_axis_bramio_2_tvalid,
    output [M_AXIS_BRAMIO_2_DMWIDTH/8-1:0] m_axis_bramio_2_tkeep,
    output [M_AXIS_BRAMIO_2_DMWIDTH/8-1:0] m_axis_bramio_2_tstrb,
    output [M_AXIS_BRAMIO_2_DMWIDTH-1:0] m_axis_bramio_2_tdata,
    input m_axis_bramio_2_tready,
    //in-out BRAM AXI-Stream output interface 3
    input m_axis_bramio_3_aclk,
    input m_axis_bramio_3_aresetn,
    output m_axis_bramio_3_tlast,
    output m_axis_bramio_3_tvalid,
    output [M_AXIS_BRAMIO_3_DMWIDTH/8-1:0] m_axis_bramio_3_tkeep,
    output [M_AXIS_BRAMIO_3_DMWIDTH/8-1:0] m_axis_bramio_3_tstrb,
    output [M_AXIS_BRAMIO_3_DMWIDTH-1:0] m_axis_bramio_3_tdata,
    input m_axis_bramio_3_tready,
    //in-out BRAM AXI-Stream output interface 4
    input m_axis_bramio_4_aclk,
    input m_axis_bramio_4_aresetn,
    output m_axis_bramio_4_tlast,
    output m_axis_bramio_4_tvalid,
    output [M_AXIS_BRAMIO_4_DMWIDTH/8-1:0] m_axis_bramio_4_tkeep,
    output [M_AXIS_BRAMIO_4_DMWIDTH/8-1:0] m_axis_bramio_4_tstrb,
    output [M_AXIS_BRAMIO_4_DMWIDTH-1:0] m_axis_bramio_4_tdata,
    input m_axis_bramio_4_tready,
    //in-out BRAM AXI-Stream output interface 5
    input m_axis_bramio_5_aclk,
    input m_axis_bramio_5_aresetn,
    output m_axis_bramio_5_tlast,
    output m_axis_bramio_5_tvalid,
    output [M_AXIS_BRAMIO_5_DMWIDTH/8-1:0] m_axis_bramio_5_tkeep,
    output [M_AXIS_BRAMIO_5_DMWIDTH/8-1:0] m_axis_bramio_5_tstrb,
    output [M_AXIS_BRAMIO_5_DMWIDTH-1:0] m_axis_bramio_5_tdata,
    input m_axis_bramio_5_tready,
    //in-out BRAM AXI-Stream output interface 6
    input m_axis_bramio_6_aclk,
    input m_axis_bramio_6_aresetn,
    output m_axis_bramio_6_tlast,
    output m_axis_bramio_6_tvalid,
    output [M_AXIS_BRAMIO_6_DMWIDTH/8-1:0] m_axis_bramio_6_tkeep,
    output [M_AXIS_BRAMIO_6_DMWIDTH/8-1:0] m_axis_bramio_6_tstrb,
    output [M_AXIS_BRAMIO_6_DMWIDTH-1:0] m_axis_bramio_6_tdata,
    input m_axis_bramio_6_tready,
    //in-out BRAM AXI-Stream output interface 7
    input m_axis_bramio_7_aclk,
    input m_axis_bramio_7_aresetn,
    output m_axis_bramio_7_tlast,
    output m_axis_bramio_7_tvalid,
    output [M_AXIS_BRAMIO_7_DMWIDTH/8-1:0] m_axis_bramio_7_tkeep,
    output [M_AXIS_BRAMIO_7_DMWIDTH/8-1:0] m_axis_bramio_7_tstrb,
    output [M_AXIS_BRAMIO_7_DMWIDTH-1:0] m_axis_bramio_7_tdata,
    input m_axis_bramio_7_tready,
    //in-out BRAM AXI-Stream output interface 8
    input m_axis_bramio_8_aclk,
    input m_axis_bramio_8_aresetn,
    output m_axis_bramio_8_tlast,
    output m_axis_bramio_8_tvalid,
    output [M_AXIS_BRAMIO_8_DMWIDTH/8-1:0] m_axis_bramio_8_tkeep,
    output [M_AXIS_BRAMIO_8_DMWIDTH/8-1:0] m_axis_bramio_8_tstrb,
    output [M_AXIS_BRAMIO_8_DMWIDTH-1:0] m_axis_bramio_8_tdata,
    input m_axis_bramio_8_tready,
    //in-out BRAM AXI-Stream output interface 9
    input m_axis_bramio_9_aclk,
    input m_axis_bramio_9_aresetn,
    output m_axis_bramio_9_tlast,
    output m_axis_bramio_9_tvalid,
    output [M_AXIS_BRAMIO_9_DMWIDTH/8-1:0] m_axis_bramio_9_tkeep,
    output [M_AXIS_BRAMIO_9_DMWIDTH/8-1:0] m_axis_bramio_9_tstrb,
    output [M_AXIS_BRAMIO_9_DMWIDTH-1:0] m_axis_bramio_9_tdata,
    input m_axis_bramio_9_tready,
    //in-out BRAM AXI-Stream output interface 10
    input m_axis_bramio_10_aclk,
    input m_axis_bramio_10_aresetn,
    output m_axis_bramio_10_tlast,
    output m_axis_bramio_10_tvalid,
    output [M_AXIS_BRAMIO_10_DMWIDTH/8-1:0] m_axis_bramio_10_tkeep,
    output [M_AXIS_BRAMIO_10_DMWIDTH/8-1:0] m_axis_bramio_10_tstrb,
    output [M_AXIS_BRAMIO_10_DMWIDTH-1:0] m_axis_bramio_10_tdata,
    input m_axis_bramio_10_tready,
    //in-out BRAM AXI-Stream output interface 11
    input m_axis_bramio_11_aclk,
    input m_axis_bramio_11_aresetn,
    output m_axis_bramio_11_tlast,
    output m_axis_bramio_11_tvalid,
    output [M_AXIS_BRAMIO_11_DMWIDTH/8-1:0] m_axis_bramio_11_tkeep,
    output [M_AXIS_BRAMIO_11_DMWIDTH/8-1:0] m_axis_bramio_11_tstrb,
    output [M_AXIS_BRAMIO_11_DMWIDTH-1:0] m_axis_bramio_11_tdata,
    input m_axis_bramio_11_tready,
    //in-out BRAM AXI-Stream output interface 12
    input m_axis_bramio_12_aclk,
    input m_axis_bramio_12_aresetn,
    output m_axis_bramio_12_tlast,
    output m_axis_bramio_12_tvalid,
    output [M_AXIS_BRAMIO_12_DMWIDTH/8-1:0] m_axis_bramio_12_tkeep,
    output [M_AXIS_BRAMIO_12_DMWIDTH/8-1:0] m_axis_bramio_12_tstrb,
    output [M_AXIS_BRAMIO_12_DMWIDTH-1:0] m_axis_bramio_12_tdata,
    input m_axis_bramio_12_tready,
    //in-out BRAM AXI-Stream output interface 13
    input m_axis_bramio_13_aclk,
    input m_axis_bramio_13_aresetn,
    output m_axis_bramio_13_tlast,
    output m_axis_bramio_13_tvalid,
    output [M_AXIS_BRAMIO_13_DMWIDTH/8-1:0] m_axis_bramio_13_tkeep,
    output [M_AXIS_BRAMIO_13_DMWIDTH/8-1:0] m_axis_bramio_13_tstrb,
    output [M_AXIS_BRAMIO_13_DMWIDTH-1:0] m_axis_bramio_13_tdata,
    input m_axis_bramio_13_tready,
    //in-out BRAM AXI-Stream output interface 14
    input m_axis_bramio_14_aclk,
    input m_axis_bramio_14_aresetn,
    output m_axis_bramio_14_tlast,
    output m_axis_bramio_14_tvalid,
    output [M_AXIS_BRAMIO_14_DMWIDTH/8-1:0] m_axis_bramio_14_tkeep,
    output [M_AXIS_BRAMIO_14_DMWIDTH/8-1:0] m_axis_bramio_14_tstrb,
    output [M_AXIS_BRAMIO_14_DMWIDTH-1:0] m_axis_bramio_14_tdata,
    input m_axis_bramio_14_tready,
    //in-out BRAM AXI-Stream output interface 15
    input m_axis_bramio_15_aclk,
    input m_axis_bramio_15_aresetn,
    output m_axis_bramio_15_tlast,
    output m_axis_bramio_15_tvalid,
    output [M_AXIS_BRAMIO_15_DMWIDTH/8-1:0] m_axis_bramio_15_tkeep,
    output [M_AXIS_BRAMIO_15_DMWIDTH/8-1:0] m_axis_bramio_15_tstrb,
    output [M_AXIS_BRAMIO_15_DMWIDTH-1:0] m_axis_bramio_15_tdata,
    input m_axis_bramio_15_tready,
    //in-out BRAM AXI-Stream output interface 16
    input m_axis_bramio_16_aclk,
    input m_axis_bramio_16_aresetn,
    output m_axis_bramio_16_tlast,
    output m_axis_bramio_16_tvalid,
    output [M_AXIS_BRAMIO_16_DMWIDTH/8-1:0] m_axis_bramio_16_tkeep,
    output [M_AXIS_BRAMIO_16_DMWIDTH/8-1:0] m_axis_bramio_16_tstrb,
    output [M_AXIS_BRAMIO_16_DMWIDTH-1:0] m_axis_bramio_16_tdata,
    input m_axis_bramio_16_tready,
    //in-out BRAM AXI-Stream output interface 17
    input m_axis_bramio_17_aclk,
    input m_axis_bramio_17_aresetn,
    output m_axis_bramio_17_tlast,
    output m_axis_bramio_17_tvalid,
    output [M_AXIS_BRAMIO_17_DMWIDTH/8-1:0] m_axis_bramio_17_tkeep,
    output [M_AXIS_BRAMIO_17_DMWIDTH/8-1:0] m_axis_bramio_17_tstrb,
    output [M_AXIS_BRAMIO_17_DMWIDTH-1:0] m_axis_bramio_17_tdata,
    input m_axis_bramio_17_tready,
    //in-out BRAM AXI-Stream output interface 18
    input m_axis_bramio_18_aclk,
    input m_axis_bramio_18_aresetn,
    output m_axis_bramio_18_tlast,
    output m_axis_bramio_18_tvalid,
    output [M_AXIS_BRAMIO_18_DMWIDTH/8-1:0] m_axis_bramio_18_tkeep,
    output [M_AXIS_BRAMIO_18_DMWIDTH/8-1:0] m_axis_bramio_18_tstrb,
    output [M_AXIS_BRAMIO_18_DMWIDTH-1:0] m_axis_bramio_18_tdata,
    input m_axis_bramio_18_tready,
    //in-out BRAM AXI-Stream output interface 19
    input m_axis_bramio_19_aclk,
    input m_axis_bramio_19_aresetn,
    output m_axis_bramio_19_tlast,
    output m_axis_bramio_19_tvalid,
    output [M_AXIS_BRAMIO_19_DMWIDTH/8-1:0] m_axis_bramio_19_tkeep,
    output [M_AXIS_BRAMIO_19_DMWIDTH/8-1:0] m_axis_bramio_19_tstrb,
    output [M_AXIS_BRAMIO_19_DMWIDTH-1:0] m_axis_bramio_19_tdata,
    input m_axis_bramio_19_tready,
    //in-out BRAM AXI-Stream output interface 20
    input m_axis_bramio_20_aclk,
    input m_axis_bramio_20_aresetn,
    output m_axis_bramio_20_tlast,
    output m_axis_bramio_20_tvalid,
    output [M_AXIS_BRAMIO_20_DMWIDTH/8-1:0] m_axis_bramio_20_tkeep,
    output [M_AXIS_BRAMIO_20_DMWIDTH/8-1:0] m_axis_bramio_20_tstrb,
    output [M_AXIS_BRAMIO_20_DMWIDTH-1:0] m_axis_bramio_20_tdata,
    input m_axis_bramio_20_tready,
    //in-out BRAM AXI-Stream output interface 21
    input m_axis_bramio_21_aclk,
    input m_axis_bramio_21_aresetn,
    output m_axis_bramio_21_tlast,
    output m_axis_bramio_21_tvalid,
    output [M_AXIS_BRAMIO_21_DMWIDTH/8-1:0] m_axis_bramio_21_tkeep,
    output [M_AXIS_BRAMIO_21_DMWIDTH/8-1:0] m_axis_bramio_21_tstrb,
    output [M_AXIS_BRAMIO_21_DMWIDTH-1:0] m_axis_bramio_21_tdata,
    input m_axis_bramio_21_tready,
    //in-out BRAM AXI-Stream output interface 22
    input m_axis_bramio_22_aclk,
    input m_axis_bramio_22_aresetn,
    output m_axis_bramio_22_tlast,
    output m_axis_bramio_22_tvalid,
    output [M_AXIS_BRAMIO_22_DMWIDTH/8-1:0] m_axis_bramio_22_tkeep,
    output [M_AXIS_BRAMIO_22_DMWIDTH/8-1:0] m_axis_bramio_22_tstrb,
    output [M_AXIS_BRAMIO_22_DMWIDTH-1:0] m_axis_bramio_22_tdata,
    input m_axis_bramio_22_tready,
    //in-out BRAM AXI-Stream output interface 23
    input m_axis_bramio_23_aclk,
    input m_axis_bramio_23_aresetn,
    output m_axis_bramio_23_tlast,
    output m_axis_bramio_23_tvalid,
    output [M_AXIS_BRAMIO_23_DMWIDTH/8-1:0] m_axis_bramio_23_tkeep,
    output [M_AXIS_BRAMIO_23_DMWIDTH/8-1:0] m_axis_bramio_23_tstrb,
    output [M_AXIS_BRAMIO_23_DMWIDTH-1:0] m_axis_bramio_23_tdata,
    input m_axis_bramio_23_tready,
    //in-out BRAM AXI-Stream output interface 24
    input m_axis_bramio_24_aclk,
    input m_axis_bramio_24_aresetn,
    output m_axis_bramio_24_tlast,
    output m_axis_bramio_24_tvalid,
    output [M_AXIS_BRAMIO_24_DMWIDTH/8-1:0] m_axis_bramio_24_tkeep,
    output [M_AXIS_BRAMIO_24_DMWIDTH/8-1:0] m_axis_bramio_24_tstrb,
    output [M_AXIS_BRAMIO_24_DMWIDTH-1:0] m_axis_bramio_24_tdata,
    input m_axis_bramio_24_tready,
    //in-out BRAM AXI-Stream output interface 25
    input m_axis_bramio_25_aclk,
    input m_axis_bramio_25_aresetn,
    output m_axis_bramio_25_tlast,
    output m_axis_bramio_25_tvalid,
    output [M_AXIS_BRAMIO_25_DMWIDTH/8-1:0] m_axis_bramio_25_tkeep,
    output [M_AXIS_BRAMIO_25_DMWIDTH/8-1:0] m_axis_bramio_25_tstrb,
    output [M_AXIS_BRAMIO_25_DMWIDTH-1:0] m_axis_bramio_25_tdata,
    input m_axis_bramio_25_tready,
    //in-out BRAM AXI-Stream output interface 26
    input m_axis_bramio_26_aclk,
    input m_axis_bramio_26_aresetn,
    output m_axis_bramio_26_tlast,
    output m_axis_bramio_26_tvalid,
    output [M_AXIS_BRAMIO_26_DMWIDTH/8-1:0] m_axis_bramio_26_tkeep,
    output [M_AXIS_BRAMIO_26_DMWIDTH/8-1:0] m_axis_bramio_26_tstrb,
    output [M_AXIS_BRAMIO_26_DMWIDTH-1:0] m_axis_bramio_26_tdata,
    input m_axis_bramio_26_tready,
    //in-out BRAM AXI-Stream output interface 27
    input m_axis_bramio_27_aclk,
    input m_axis_bramio_27_aresetn,
    output m_axis_bramio_27_tlast,
    output m_axis_bramio_27_tvalid,
    output [M_AXIS_BRAMIO_27_DMWIDTH/8-1:0] m_axis_bramio_27_tkeep,
    output [M_AXIS_BRAMIO_27_DMWIDTH/8-1:0] m_axis_bramio_27_tstrb,
    output [M_AXIS_BRAMIO_27_DMWIDTH-1:0] m_axis_bramio_27_tdata,
    input m_axis_bramio_27_tready,
    //in-out BRAM AXI-Stream output interface 28
    input m_axis_bramio_28_aclk,
    input m_axis_bramio_28_aresetn,
    output m_axis_bramio_28_tlast,
    output m_axis_bramio_28_tvalid,
    output [M_AXIS_BRAMIO_28_DMWIDTH/8-1:0] m_axis_bramio_28_tkeep,
    output [M_AXIS_BRAMIO_28_DMWIDTH/8-1:0] m_axis_bramio_28_tstrb,
    output [M_AXIS_BRAMIO_28_DMWIDTH-1:0] m_axis_bramio_28_tdata,
    input m_axis_bramio_28_tready,
    //in-out BRAM AXI-Stream output interface 29
    input m_axis_bramio_29_aclk,
    input m_axis_bramio_29_aresetn,
    output m_axis_bramio_29_tlast,
    output m_axis_bramio_29_tvalid,
    output [M_AXIS_BRAMIO_29_DMWIDTH/8-1:0] m_axis_bramio_29_tkeep,
    output [M_AXIS_BRAMIO_29_DMWIDTH/8-1:0] m_axis_bramio_29_tstrb,
    output [M_AXIS_BRAMIO_29_DMWIDTH-1:0] m_axis_bramio_29_tdata,
    input m_axis_bramio_29_tready,
    //in-out BRAM AXI-Stream output interface 30
    input m_axis_bramio_30_aclk,
    input m_axis_bramio_30_aresetn,
    output m_axis_bramio_30_tlast,
    output m_axis_bramio_30_tvalid,
    output [M_AXIS_BRAMIO_30_DMWIDTH/8-1:0] m_axis_bramio_30_tkeep,
    output [M_AXIS_BRAMIO_30_DMWIDTH/8-1:0] m_axis_bramio_30_tstrb,
    output [M_AXIS_BRAMIO_30_DMWIDTH-1:0] m_axis_bramio_30_tdata,
    input m_axis_bramio_30_tready,
    //in-out BRAM AXI-Stream output interface 31
    input m_axis_bramio_31_aclk,
    input m_axis_bramio_31_aresetn,
    output m_axis_bramio_31_tlast,
    output m_axis_bramio_31_tvalid,
    output [M_AXIS_BRAMIO_31_DMWIDTH/8-1:0] m_axis_bramio_31_tkeep,
    output [M_AXIS_BRAMIO_31_DMWIDTH/8-1:0] m_axis_bramio_31_tstrb,
    output [M_AXIS_BRAMIO_31_DMWIDTH-1:0] m_axis_bramio_31_tdata,
    input m_axis_bramio_31_tready,
    //in-out BRAM AXI-Stream output interface 32
    input m_axis_bramio_32_aclk,
    input m_axis_bramio_32_aresetn,
    output m_axis_bramio_32_tlast,
    output m_axis_bramio_32_tvalid,
    output [M_AXIS_BRAMIO_32_DMWIDTH/8-1:0] m_axis_bramio_32_tkeep,
    output [M_AXIS_BRAMIO_32_DMWIDTH/8-1:0] m_axis_bramio_32_tstrb,
    output [M_AXIS_BRAMIO_32_DMWIDTH-1:0] m_axis_bramio_32_tdata,
    input m_axis_bramio_32_tready,
    //in-out BRAM AXI-Stream output interface 33
    input m_axis_bramio_33_aclk,
    input m_axis_bramio_33_aresetn,
    output m_axis_bramio_33_tlast,
    output m_axis_bramio_33_tvalid,
    output [M_AXIS_BRAMIO_33_DMWIDTH/8-1:0] m_axis_bramio_33_tkeep,
    output [M_AXIS_BRAMIO_33_DMWIDTH/8-1:0] m_axis_bramio_33_tstrb,
    output [M_AXIS_BRAMIO_33_DMWIDTH-1:0] m_axis_bramio_33_tdata,
    input m_axis_bramio_33_tready,
    //in-out BRAM AXI-Stream output interface 34
    input m_axis_bramio_34_aclk,
    input m_axis_bramio_34_aresetn,
    output m_axis_bramio_34_tlast,
    output m_axis_bramio_34_tvalid,
    output [M_AXIS_BRAMIO_34_DMWIDTH/8-1:0] m_axis_bramio_34_tkeep,
    output [M_AXIS_BRAMIO_34_DMWIDTH/8-1:0] m_axis_bramio_34_tstrb,
    output [M_AXIS_BRAMIO_34_DMWIDTH-1:0] m_axis_bramio_34_tdata,
    input m_axis_bramio_34_tready,
    //in-out BRAM AXI-Stream output interface 35
    input m_axis_bramio_35_aclk,
    input m_axis_bramio_35_aresetn,
    output m_axis_bramio_35_tlast,
    output m_axis_bramio_35_tvalid,
    output [M_AXIS_BRAMIO_35_DMWIDTH/8-1:0] m_axis_bramio_35_tkeep,
    output [M_AXIS_BRAMIO_35_DMWIDTH/8-1:0] m_axis_bramio_35_tstrb,
    output [M_AXIS_BRAMIO_35_DMWIDTH-1:0] m_axis_bramio_35_tdata,
    input m_axis_bramio_35_tready,
    //in-out BRAM AXI-Stream output interface 36
    input m_axis_bramio_36_aclk,
    input m_axis_bramio_36_aresetn,
    output m_axis_bramio_36_tlast,
    output m_axis_bramio_36_tvalid,
    output [M_AXIS_BRAMIO_36_DMWIDTH/8-1:0] m_axis_bramio_36_tkeep,
    output [M_AXIS_BRAMIO_36_DMWIDTH/8-1:0] m_axis_bramio_36_tstrb,
    output [M_AXIS_BRAMIO_36_DMWIDTH-1:0] m_axis_bramio_36_tdata,
    input m_axis_bramio_36_tready,
    //in-out BRAM AXI-Stream output interface 37
    input m_axis_bramio_37_aclk,
    input m_axis_bramio_37_aresetn,
    output m_axis_bramio_37_tlast,
    output m_axis_bramio_37_tvalid,
    output [M_AXIS_BRAMIO_37_DMWIDTH/8-1:0] m_axis_bramio_37_tkeep,
    output [M_AXIS_BRAMIO_37_DMWIDTH/8-1:0] m_axis_bramio_37_tstrb,
    output [M_AXIS_BRAMIO_37_DMWIDTH-1:0] m_axis_bramio_37_tdata,
    input m_axis_bramio_37_tready,
    //in-out BRAM AXI-Stream output interface 38
    input m_axis_bramio_38_aclk,
    input m_axis_bramio_38_aresetn,
    output m_axis_bramio_38_tlast,
    output m_axis_bramio_38_tvalid,
    output [M_AXIS_BRAMIO_38_DMWIDTH/8-1:0] m_axis_bramio_38_tkeep,
    output [M_AXIS_BRAMIO_38_DMWIDTH/8-1:0] m_axis_bramio_38_tstrb,
    output [M_AXIS_BRAMIO_38_DMWIDTH-1:0] m_axis_bramio_38_tdata,
    input m_axis_bramio_38_tready,
    //in-out BRAM AXI-Stream output interface 39
    input m_axis_bramio_39_aclk,
    input m_axis_bramio_39_aresetn,
    output m_axis_bramio_39_tlast,
    output m_axis_bramio_39_tvalid,
    output [M_AXIS_BRAMIO_39_DMWIDTH/8-1:0] m_axis_bramio_39_tkeep,
    output [M_AXIS_BRAMIO_39_DMWIDTH/8-1:0] m_axis_bramio_39_tstrb,
    output [M_AXIS_BRAMIO_39_DMWIDTH-1:0] m_axis_bramio_39_tdata,
    input m_axis_bramio_39_tready,
    //in-out BRAM AXI-Stream output interface 40
    input m_axis_bramio_40_aclk,
    input m_axis_bramio_40_aresetn,
    output m_axis_bramio_40_tlast,
    output m_axis_bramio_40_tvalid,
    output [M_AXIS_BRAMIO_40_DMWIDTH/8-1:0] m_axis_bramio_40_tkeep,
    output [M_AXIS_BRAMIO_40_DMWIDTH/8-1:0] m_axis_bramio_40_tstrb,
    output [M_AXIS_BRAMIO_40_DMWIDTH-1:0] m_axis_bramio_40_tdata,
    input m_axis_bramio_40_tready,
    //in-out BRAM AXI-Stream output interface 41
    input m_axis_bramio_41_aclk,
    input m_axis_bramio_41_aresetn,
    output m_axis_bramio_41_tlast,
    output m_axis_bramio_41_tvalid,
    output [M_AXIS_BRAMIO_41_DMWIDTH/8-1:0] m_axis_bramio_41_tkeep,
    output [M_AXIS_BRAMIO_41_DMWIDTH/8-1:0] m_axis_bramio_41_tstrb,
    output [M_AXIS_BRAMIO_41_DMWIDTH-1:0] m_axis_bramio_41_tdata,
    input m_axis_bramio_41_tready,
    //in-out BRAM AXI-Stream output interface 42
    input m_axis_bramio_42_aclk,
    input m_axis_bramio_42_aresetn,
    output m_axis_bramio_42_tlast,
    output m_axis_bramio_42_tvalid,
    output [M_AXIS_BRAMIO_42_DMWIDTH/8-1:0] m_axis_bramio_42_tkeep,
    output [M_AXIS_BRAMIO_42_DMWIDTH/8-1:0] m_axis_bramio_42_tstrb,
    output [M_AXIS_BRAMIO_42_DMWIDTH-1:0] m_axis_bramio_42_tdata,
    input m_axis_bramio_42_tready,
    //in-out BRAM AXI-Stream output interface 43
    input m_axis_bramio_43_aclk,
    input m_axis_bramio_43_aresetn,
    output m_axis_bramio_43_tlast,
    output m_axis_bramio_43_tvalid,
    output [M_AXIS_BRAMIO_43_DMWIDTH/8-1:0] m_axis_bramio_43_tkeep,
    output [M_AXIS_BRAMIO_43_DMWIDTH/8-1:0] m_axis_bramio_43_tstrb,
    output [M_AXIS_BRAMIO_43_DMWIDTH-1:0] m_axis_bramio_43_tdata,
    input m_axis_bramio_43_tready,
    //in-out BRAM AXI-Stream output interface 44
    input m_axis_bramio_44_aclk,
    input m_axis_bramio_44_aresetn,
    output m_axis_bramio_44_tlast,
    output m_axis_bramio_44_tvalid,
    output [M_AXIS_BRAMIO_44_DMWIDTH/8-1:0] m_axis_bramio_44_tkeep,
    output [M_AXIS_BRAMIO_44_DMWIDTH/8-1:0] m_axis_bramio_44_tstrb,
    output [M_AXIS_BRAMIO_44_DMWIDTH-1:0] m_axis_bramio_44_tdata,
    input m_axis_bramio_44_tready,
    //in-out BRAM AXI-Stream output interface 45
    input m_axis_bramio_45_aclk,
    input m_axis_bramio_45_aresetn,
    output m_axis_bramio_45_tlast,
    output m_axis_bramio_45_tvalid,
    output [M_AXIS_BRAMIO_45_DMWIDTH/8-1:0] m_axis_bramio_45_tkeep,
    output [M_AXIS_BRAMIO_45_DMWIDTH/8-1:0] m_axis_bramio_45_tstrb,
    output [M_AXIS_BRAMIO_45_DMWIDTH-1:0] m_axis_bramio_45_tdata,
    input m_axis_bramio_45_tready,
    //in-out BRAM AXI-Stream output interface 46
    input m_axis_bramio_46_aclk,
    input m_axis_bramio_46_aresetn,
    output m_axis_bramio_46_tlast,
    output m_axis_bramio_46_tvalid,
    output [M_AXIS_BRAMIO_46_DMWIDTH/8-1:0] m_axis_bramio_46_tkeep,
    output [M_AXIS_BRAMIO_46_DMWIDTH/8-1:0] m_axis_bramio_46_tstrb,
    output [M_AXIS_BRAMIO_46_DMWIDTH-1:0] m_axis_bramio_46_tdata,
    input m_axis_bramio_46_tready,
    //in-out BRAM AXI-Stream output interface 47
    input m_axis_bramio_47_aclk,
    input m_axis_bramio_47_aresetn,
    output m_axis_bramio_47_tlast,
    output m_axis_bramio_47_tvalid,
    output [M_AXIS_BRAMIO_47_DMWIDTH/8-1:0] m_axis_bramio_47_tkeep,
    output [M_AXIS_BRAMIO_47_DMWIDTH/8-1:0] m_axis_bramio_47_tstrb,
    output [M_AXIS_BRAMIO_47_DMWIDTH-1:0] m_axis_bramio_47_tdata,
    input m_axis_bramio_47_tready,
    //in-out BRAM AXI-Stream output interface 48
    input m_axis_bramio_48_aclk,
    input m_axis_bramio_48_aresetn,
    output m_axis_bramio_48_tlast,
    output m_axis_bramio_48_tvalid,
    output [M_AXIS_BRAMIO_48_DMWIDTH/8-1:0] m_axis_bramio_48_tkeep,
    output [M_AXIS_BRAMIO_48_DMWIDTH/8-1:0] m_axis_bramio_48_tstrb,
    output [M_AXIS_BRAMIO_48_DMWIDTH-1:0] m_axis_bramio_48_tdata,
    input m_axis_bramio_48_tready,
    //in-out BRAM AXI-Stream output interface 49
    input m_axis_bramio_49_aclk,
    input m_axis_bramio_49_aresetn,
    output m_axis_bramio_49_tlast,
    output m_axis_bramio_49_tvalid,
    output [M_AXIS_BRAMIO_49_DMWIDTH/8-1:0] m_axis_bramio_49_tkeep,
    output [M_AXIS_BRAMIO_49_DMWIDTH/8-1:0] m_axis_bramio_49_tstrb,
    output [M_AXIS_BRAMIO_49_DMWIDTH-1:0] m_axis_bramio_49_tdata,
    input m_axis_bramio_49_tready,
    //in-out BRAM AXI-Stream output interface 50
    input m_axis_bramio_50_aclk,
    input m_axis_bramio_50_aresetn,
    output m_axis_bramio_50_tlast,
    output m_axis_bramio_50_tvalid,
    output [M_AXIS_BRAMIO_50_DMWIDTH/8-1:0] m_axis_bramio_50_tkeep,
    output [M_AXIS_BRAMIO_50_DMWIDTH/8-1:0] m_axis_bramio_50_tstrb,
    output [M_AXIS_BRAMIO_50_DMWIDTH-1:0] m_axis_bramio_50_tdata,
    input m_axis_bramio_50_tready,
    //in-out BRAM AXI-Stream output interface 51
    input m_axis_bramio_51_aclk,
    input m_axis_bramio_51_aresetn,
    output m_axis_bramio_51_tlast,
    output m_axis_bramio_51_tvalid,
    output [M_AXIS_BRAMIO_51_DMWIDTH/8-1:0] m_axis_bramio_51_tkeep,
    output [M_AXIS_BRAMIO_51_DMWIDTH/8-1:0] m_axis_bramio_51_tstrb,
    output [M_AXIS_BRAMIO_51_DMWIDTH-1:0] m_axis_bramio_51_tdata,
    input m_axis_bramio_51_tready,
    //in-out BRAM AXI-Stream output interface 52
    input m_axis_bramio_52_aclk,
    input m_axis_bramio_52_aresetn,
    output m_axis_bramio_52_tlast,
    output m_axis_bramio_52_tvalid,
    output [M_AXIS_BRAMIO_52_DMWIDTH/8-1:0] m_axis_bramio_52_tkeep,
    output [M_AXIS_BRAMIO_52_DMWIDTH/8-1:0] m_axis_bramio_52_tstrb,
    output [M_AXIS_BRAMIO_52_DMWIDTH-1:0] m_axis_bramio_52_tdata,
    input m_axis_bramio_52_tready,
    //in-out BRAM AXI-Stream output interface 53
    input m_axis_bramio_53_aclk,
    input m_axis_bramio_53_aresetn,
    output m_axis_bramio_53_tlast,
    output m_axis_bramio_53_tvalid,
    output [M_AXIS_BRAMIO_53_DMWIDTH/8-1:0] m_axis_bramio_53_tkeep,
    output [M_AXIS_BRAMIO_53_DMWIDTH/8-1:0] m_axis_bramio_53_tstrb,
    output [M_AXIS_BRAMIO_53_DMWIDTH-1:0] m_axis_bramio_53_tdata,
    input m_axis_bramio_53_tready,
    //in-out BRAM AXI-Stream output interface 54
    input m_axis_bramio_54_aclk,
    input m_axis_bramio_54_aresetn,
    output m_axis_bramio_54_tlast,
    output m_axis_bramio_54_tvalid,
    output [M_AXIS_BRAMIO_54_DMWIDTH/8-1:0] m_axis_bramio_54_tkeep,
    output [M_AXIS_BRAMIO_54_DMWIDTH/8-1:0] m_axis_bramio_54_tstrb,
    output [M_AXIS_BRAMIO_54_DMWIDTH-1:0] m_axis_bramio_54_tdata,
    input m_axis_bramio_54_tready,
    //in-out BRAM AXI-Stream output interface 55
    input m_axis_bramio_55_aclk,
    input m_axis_bramio_55_aresetn,
    output m_axis_bramio_55_tlast,
    output m_axis_bramio_55_tvalid,
    output [M_AXIS_BRAMIO_55_DMWIDTH/8-1:0] m_axis_bramio_55_tkeep,
    output [M_AXIS_BRAMIO_55_DMWIDTH/8-1:0] m_axis_bramio_55_tstrb,
    output [M_AXIS_BRAMIO_55_DMWIDTH-1:0] m_axis_bramio_55_tdata,
    input m_axis_bramio_55_tready,
    //in-out BRAM AXI-Stream output interface 56
    input m_axis_bramio_56_aclk,
    input m_axis_bramio_56_aresetn,
    output m_axis_bramio_56_tlast,
    output m_axis_bramio_56_tvalid,
    output [M_AXIS_BRAMIO_56_DMWIDTH/8-1:0] m_axis_bramio_56_tkeep,
    output [M_AXIS_BRAMIO_56_DMWIDTH/8-1:0] m_axis_bramio_56_tstrb,
    output [M_AXIS_BRAMIO_56_DMWIDTH-1:0] m_axis_bramio_56_tdata,
    input m_axis_bramio_56_tready,
    //in-out BRAM AXI-Stream output interface 57
    input m_axis_bramio_57_aclk,
    input m_axis_bramio_57_aresetn,
    output m_axis_bramio_57_tlast,
    output m_axis_bramio_57_tvalid,
    output [M_AXIS_BRAMIO_57_DMWIDTH/8-1:0] m_axis_bramio_57_tkeep,
    output [M_AXIS_BRAMIO_57_DMWIDTH/8-1:0] m_axis_bramio_57_tstrb,
    output [M_AXIS_BRAMIO_57_DMWIDTH-1:0] m_axis_bramio_57_tdata,
    input m_axis_bramio_57_tready,
    //in-out BRAM AXI-Stream output interface 58
    input m_axis_bramio_58_aclk,
    input m_axis_bramio_58_aresetn,
    output m_axis_bramio_58_tlast,
    output m_axis_bramio_58_tvalid,
    output [M_AXIS_BRAMIO_58_DMWIDTH/8-1:0] m_axis_bramio_58_tkeep,
    output [M_AXIS_BRAMIO_58_DMWIDTH/8-1:0] m_axis_bramio_58_tstrb,
    output [M_AXIS_BRAMIO_58_DMWIDTH-1:0] m_axis_bramio_58_tdata,
    input m_axis_bramio_58_tready,
    //in-out BRAM AXI-Stream output interface 59
    input m_axis_bramio_59_aclk,
    input m_axis_bramio_59_aresetn,
    output m_axis_bramio_59_tlast,
    output m_axis_bramio_59_tvalid,
    output [M_AXIS_BRAMIO_59_DMWIDTH/8-1:0] m_axis_bramio_59_tkeep,
    output [M_AXIS_BRAMIO_59_DMWIDTH/8-1:0] m_axis_bramio_59_tstrb,
    output [M_AXIS_BRAMIO_59_DMWIDTH-1:0] m_axis_bramio_59_tdata,
    input m_axis_bramio_59_tready,
    //in-out BRAM AXI-Stream output interface 60
    input m_axis_bramio_60_aclk,
    input m_axis_bramio_60_aresetn,
    output m_axis_bramio_60_tlast,
    output m_axis_bramio_60_tvalid,
    output [M_AXIS_BRAMIO_60_DMWIDTH/8-1:0] m_axis_bramio_60_tkeep,
    output [M_AXIS_BRAMIO_60_DMWIDTH/8-1:0] m_axis_bramio_60_tstrb,
    output [M_AXIS_BRAMIO_60_DMWIDTH-1:0] m_axis_bramio_60_tdata,
    input m_axis_bramio_60_tready,
    //in-out BRAM AXI-Stream output interface 61
    input m_axis_bramio_61_aclk,
    input m_axis_bramio_61_aresetn,
    output m_axis_bramio_61_tlast,
    output m_axis_bramio_61_tvalid,
    output [M_AXIS_BRAMIO_61_DMWIDTH/8-1:0] m_axis_bramio_61_tkeep,
    output [M_AXIS_BRAMIO_61_DMWIDTH/8-1:0] m_axis_bramio_61_tstrb,
    output [M_AXIS_BRAMIO_61_DMWIDTH-1:0] m_axis_bramio_61_tdata,
    input m_axis_bramio_61_tready,
    //in-out BRAM AXI-Stream output interface 62
    input m_axis_bramio_62_aclk,
    input m_axis_bramio_62_aresetn,
    output m_axis_bramio_62_tlast,
    output m_axis_bramio_62_tvalid,
    output [M_AXIS_BRAMIO_62_DMWIDTH/8-1:0] m_axis_bramio_62_tkeep,
    output [M_AXIS_BRAMIO_62_DMWIDTH/8-1:0] m_axis_bramio_62_tstrb,
    output [M_AXIS_BRAMIO_62_DMWIDTH-1:0] m_axis_bramio_62_tdata,
    input m_axis_bramio_62_tready,
    //in-out BRAM AXI-Stream output interface 63
    input m_axis_bramio_63_aclk,
    input m_axis_bramio_63_aresetn,
    output m_axis_bramio_63_tlast,
    output m_axis_bramio_63_tvalid,
    output [M_AXIS_BRAMIO_63_DMWIDTH/8-1:0] m_axis_bramio_63_tkeep,
    output [M_AXIS_BRAMIO_63_DMWIDTH/8-1:0] m_axis_bramio_63_tstrb,
    output [M_AXIS_BRAMIO_63_DMWIDTH-1:0] m_axis_bramio_63_tdata,
    input m_axis_bramio_63_tready,
    //in-out BRAM AXI-Stream output interface 64
    input m_axis_bramio_64_aclk,
    input m_axis_bramio_64_aresetn,
    output m_axis_bramio_64_tlast,
    output m_axis_bramio_64_tvalid,
    output [M_AXIS_BRAMIO_64_DMWIDTH/8-1:0] m_axis_bramio_64_tkeep,
    output [M_AXIS_BRAMIO_64_DMWIDTH/8-1:0] m_axis_bramio_64_tstrb,
    output [M_AXIS_BRAMIO_64_DMWIDTH-1:0] m_axis_bramio_64_tdata,
    input m_axis_bramio_64_tready,
    //in-out BRAM AXI-Stream output interface 65
    input m_axis_bramio_65_aclk,
    input m_axis_bramio_65_aresetn,
    output m_axis_bramio_65_tlast,
    output m_axis_bramio_65_tvalid,
    output [M_AXIS_BRAMIO_65_DMWIDTH/8-1:0] m_axis_bramio_65_tkeep,
    output [M_AXIS_BRAMIO_65_DMWIDTH/8-1:0] m_axis_bramio_65_tstrb,
    output [M_AXIS_BRAMIO_65_DMWIDTH-1:0] m_axis_bramio_65_tdata,
    input m_axis_bramio_65_tready,
    //in-out BRAM AXI-Stream output interface 66
    input m_axis_bramio_66_aclk,
    input m_axis_bramio_66_aresetn,
    output m_axis_bramio_66_tlast,
    output m_axis_bramio_66_tvalid,
    output [M_AXIS_BRAMIO_66_DMWIDTH/8-1:0] m_axis_bramio_66_tkeep,
    output [M_AXIS_BRAMIO_66_DMWIDTH/8-1:0] m_axis_bramio_66_tstrb,
    output [M_AXIS_BRAMIO_66_DMWIDTH-1:0] m_axis_bramio_66_tdata,
    input m_axis_bramio_66_tready,
    //in-out BRAM AXI-Stream output interface 67
    input m_axis_bramio_67_aclk,
    input m_axis_bramio_67_aresetn,
    output m_axis_bramio_67_tlast,
    output m_axis_bramio_67_tvalid,
    output [M_AXIS_BRAMIO_67_DMWIDTH/8-1:0] m_axis_bramio_67_tkeep,
    output [M_AXIS_BRAMIO_67_DMWIDTH/8-1:0] m_axis_bramio_67_tstrb,
    output [M_AXIS_BRAMIO_67_DMWIDTH-1:0] m_axis_bramio_67_tdata,
    input m_axis_bramio_67_tready,
    //in-out BRAM AXI-Stream output interface 68
    input m_axis_bramio_68_aclk,
    input m_axis_bramio_68_aresetn,
    output m_axis_bramio_68_tlast,
    output m_axis_bramio_68_tvalid,
    output [M_AXIS_BRAMIO_68_DMWIDTH/8-1:0] m_axis_bramio_68_tkeep,
    output [M_AXIS_BRAMIO_68_DMWIDTH/8-1:0] m_axis_bramio_68_tstrb,
    output [M_AXIS_BRAMIO_68_DMWIDTH-1:0] m_axis_bramio_68_tdata,
    input m_axis_bramio_68_tready,
    //in-out BRAM AXI-Stream output interface 69
    input m_axis_bramio_69_aclk,
    input m_axis_bramio_69_aresetn,
    output m_axis_bramio_69_tlast,
    output m_axis_bramio_69_tvalid,
    output [M_AXIS_BRAMIO_69_DMWIDTH/8-1:0] m_axis_bramio_69_tkeep,
    output [M_AXIS_BRAMIO_69_DMWIDTH/8-1:0] m_axis_bramio_69_tstrb,
    output [M_AXIS_BRAMIO_69_DMWIDTH-1:0] m_axis_bramio_69_tdata,
    input m_axis_bramio_69_tready,
    //in-out BRAM AXI-Stream output interface 70
    input m_axis_bramio_70_aclk,
    input m_axis_bramio_70_aresetn,
    output m_axis_bramio_70_tlast,
    output m_axis_bramio_70_tvalid,
    output [M_AXIS_BRAMIO_70_DMWIDTH/8-1:0] m_axis_bramio_70_tkeep,
    output [M_AXIS_BRAMIO_70_DMWIDTH/8-1:0] m_axis_bramio_70_tstrb,
    output [M_AXIS_BRAMIO_70_DMWIDTH-1:0] m_axis_bramio_70_tdata,
    input m_axis_bramio_70_tready,
    //in-out BRAM AXI-Stream output interface 71
    input m_axis_bramio_71_aclk,
    input m_axis_bramio_71_aresetn,
    output m_axis_bramio_71_tlast,
    output m_axis_bramio_71_tvalid,
    output [M_AXIS_BRAMIO_71_DMWIDTH/8-1:0] m_axis_bramio_71_tkeep,
    output [M_AXIS_BRAMIO_71_DMWIDTH/8-1:0] m_axis_bramio_71_tstrb,
    output [M_AXIS_BRAMIO_71_DMWIDTH-1:0] m_axis_bramio_71_tdata,
    input m_axis_bramio_71_tready,
    //in-out BRAM AXI-Stream output interface 72
    input m_axis_bramio_72_aclk,
    input m_axis_bramio_72_aresetn,
    output m_axis_bramio_72_tlast,
    output m_axis_bramio_72_tvalid,
    output [M_AXIS_BRAMIO_72_DMWIDTH/8-1:0] m_axis_bramio_72_tkeep,
    output [M_AXIS_BRAMIO_72_DMWIDTH/8-1:0] m_axis_bramio_72_tstrb,
    output [M_AXIS_BRAMIO_72_DMWIDTH-1:0] m_axis_bramio_72_tdata,
    input m_axis_bramio_72_tready,
    //in-out BRAM AXI-Stream output interface 73
    input m_axis_bramio_73_aclk,
    input m_axis_bramio_73_aresetn,
    output m_axis_bramio_73_tlast,
    output m_axis_bramio_73_tvalid,
    output [M_AXIS_BRAMIO_73_DMWIDTH/8-1:0] m_axis_bramio_73_tkeep,
    output [M_AXIS_BRAMIO_73_DMWIDTH/8-1:0] m_axis_bramio_73_tstrb,
    output [M_AXIS_BRAMIO_73_DMWIDTH-1:0] m_axis_bramio_73_tdata,
    input m_axis_bramio_73_tready,
    //in-out BRAM AXI-Stream output interface 74
    input m_axis_bramio_74_aclk,
    input m_axis_bramio_74_aresetn,
    output m_axis_bramio_74_tlast,
    output m_axis_bramio_74_tvalid,
    output [M_AXIS_BRAMIO_74_DMWIDTH/8-1:0] m_axis_bramio_74_tkeep,
    output [M_AXIS_BRAMIO_74_DMWIDTH/8-1:0] m_axis_bramio_74_tstrb,
    output [M_AXIS_BRAMIO_74_DMWIDTH-1:0] m_axis_bramio_74_tdata,
    input m_axis_bramio_74_tready,
    //in-out BRAM AXI-Stream output interface 75
    input m_axis_bramio_75_aclk,
    input m_axis_bramio_75_aresetn,
    output m_axis_bramio_75_tlast,
    output m_axis_bramio_75_tvalid,
    output [M_AXIS_BRAMIO_75_DMWIDTH/8-1:0] m_axis_bramio_75_tkeep,
    output [M_AXIS_BRAMIO_75_DMWIDTH/8-1:0] m_axis_bramio_75_tstrb,
    output [M_AXIS_BRAMIO_75_DMWIDTH-1:0] m_axis_bramio_75_tdata,
    input m_axis_bramio_75_tready,
    //in-out BRAM AXI-Stream output interface 76
    input m_axis_bramio_76_aclk,
    input m_axis_bramio_76_aresetn,
    output m_axis_bramio_76_tlast,
    output m_axis_bramio_76_tvalid,
    output [M_AXIS_BRAMIO_76_DMWIDTH/8-1:0] m_axis_bramio_76_tkeep,
    output [M_AXIS_BRAMIO_76_DMWIDTH/8-1:0] m_axis_bramio_76_tstrb,
    output [M_AXIS_BRAMIO_76_DMWIDTH-1:0] m_axis_bramio_76_tdata,
    input m_axis_bramio_76_tready,
    //in-out BRAM AXI-Stream output interface 77
    input m_axis_bramio_77_aclk,
    input m_axis_bramio_77_aresetn,
    output m_axis_bramio_77_tlast,
    output m_axis_bramio_77_tvalid,
    output [M_AXIS_BRAMIO_77_DMWIDTH/8-1:0] m_axis_bramio_77_tkeep,
    output [M_AXIS_BRAMIO_77_DMWIDTH/8-1:0] m_axis_bramio_77_tstrb,
    output [M_AXIS_BRAMIO_77_DMWIDTH-1:0] m_axis_bramio_77_tdata,
    input m_axis_bramio_77_tready,
    //in-out BRAM AXI-Stream output interface 78
    input m_axis_bramio_78_aclk,
    input m_axis_bramio_78_aresetn,
    output m_axis_bramio_78_tlast,
    output m_axis_bramio_78_tvalid,
    output [M_AXIS_BRAMIO_78_DMWIDTH/8-1:0] m_axis_bramio_78_tkeep,
    output [M_AXIS_BRAMIO_78_DMWIDTH/8-1:0] m_axis_bramio_78_tstrb,
    output [M_AXIS_BRAMIO_78_DMWIDTH-1:0] m_axis_bramio_78_tdata,
    input m_axis_bramio_78_tready,
    //in-out BRAM AXI-Stream output interface 79
    input m_axis_bramio_79_aclk,
    input m_axis_bramio_79_aresetn,
    output m_axis_bramio_79_tlast,
    output m_axis_bramio_79_tvalid,
    output [M_AXIS_BRAMIO_79_DMWIDTH/8-1:0] m_axis_bramio_79_tkeep,
    output [M_AXIS_BRAMIO_79_DMWIDTH/8-1:0] m_axis_bramio_79_tstrb,
    output [M_AXIS_BRAMIO_79_DMWIDTH-1:0] m_axis_bramio_79_tdata,
    input m_axis_bramio_79_tready,
    //in-out BRAM AXI-Stream output interface 80
    input m_axis_bramio_80_aclk,
    input m_axis_bramio_80_aresetn,
    output m_axis_bramio_80_tlast,
    output m_axis_bramio_80_tvalid,
    output [M_AXIS_BRAMIO_80_DMWIDTH/8-1:0] m_axis_bramio_80_tkeep,
    output [M_AXIS_BRAMIO_80_DMWIDTH/8-1:0] m_axis_bramio_80_tstrb,
    output [M_AXIS_BRAMIO_80_DMWIDTH-1:0] m_axis_bramio_80_tdata,
    input m_axis_bramio_80_tready,
    //in-out BRAM AXI-Stream output interface 81
    input m_axis_bramio_81_aclk,
    input m_axis_bramio_81_aresetn,
    output m_axis_bramio_81_tlast,
    output m_axis_bramio_81_tvalid,
    output [M_AXIS_BRAMIO_81_DMWIDTH/8-1:0] m_axis_bramio_81_tkeep,
    output [M_AXIS_BRAMIO_81_DMWIDTH/8-1:0] m_axis_bramio_81_tstrb,
    output [M_AXIS_BRAMIO_81_DMWIDTH-1:0] m_axis_bramio_81_tdata,
    input m_axis_bramio_81_tready,
    //in-out BRAM AXI-Stream output interface 82
    input m_axis_bramio_82_aclk,
    input m_axis_bramio_82_aresetn,
    output m_axis_bramio_82_tlast,
    output m_axis_bramio_82_tvalid,
    output [M_AXIS_BRAMIO_82_DMWIDTH/8-1:0] m_axis_bramio_82_tkeep,
    output [M_AXIS_BRAMIO_82_DMWIDTH/8-1:0] m_axis_bramio_82_tstrb,
    output [M_AXIS_BRAMIO_82_DMWIDTH-1:0] m_axis_bramio_82_tdata,
    input m_axis_bramio_82_tready,
    //in-out BRAM AXI-Stream output interface 83
    input m_axis_bramio_83_aclk,
    input m_axis_bramio_83_aresetn,
    output m_axis_bramio_83_tlast,
    output m_axis_bramio_83_tvalid,
    output [M_AXIS_BRAMIO_83_DMWIDTH/8-1:0] m_axis_bramio_83_tkeep,
    output [M_AXIS_BRAMIO_83_DMWIDTH/8-1:0] m_axis_bramio_83_tstrb,
    output [M_AXIS_BRAMIO_83_DMWIDTH-1:0] m_axis_bramio_83_tdata,
    input m_axis_bramio_83_tready,
    //in-out BRAM AXI-Stream output interface 84
    input m_axis_bramio_84_aclk,
    input m_axis_bramio_84_aresetn,
    output m_axis_bramio_84_tlast,
    output m_axis_bramio_84_tvalid,
    output [M_AXIS_BRAMIO_84_DMWIDTH/8-1:0] m_axis_bramio_84_tkeep,
    output [M_AXIS_BRAMIO_84_DMWIDTH/8-1:0] m_axis_bramio_84_tstrb,
    output [M_AXIS_BRAMIO_84_DMWIDTH-1:0] m_axis_bramio_84_tdata,
    input m_axis_bramio_84_tready,
    //in-out BRAM AXI-Stream output interface 85
    input m_axis_bramio_85_aclk,
    input m_axis_bramio_85_aresetn,
    output m_axis_bramio_85_tlast,
    output m_axis_bramio_85_tvalid,
    output [M_AXIS_BRAMIO_85_DMWIDTH/8-1:0] m_axis_bramio_85_tkeep,
    output [M_AXIS_BRAMIO_85_DMWIDTH/8-1:0] m_axis_bramio_85_tstrb,
    output [M_AXIS_BRAMIO_85_DMWIDTH-1:0] m_axis_bramio_85_tdata,
    input m_axis_bramio_85_tready,
    //in-out BRAM AXI-Stream output interface 86
    input m_axis_bramio_86_aclk,
    input m_axis_bramio_86_aresetn,
    output m_axis_bramio_86_tlast,
    output m_axis_bramio_86_tvalid,
    output [M_AXIS_BRAMIO_86_DMWIDTH/8-1:0] m_axis_bramio_86_tkeep,
    output [M_AXIS_BRAMIO_86_DMWIDTH/8-1:0] m_axis_bramio_86_tstrb,
    output [M_AXIS_BRAMIO_86_DMWIDTH-1:0] m_axis_bramio_86_tdata,
    input m_axis_bramio_86_tready,
    //in-out BRAM AXI-Stream output interface 87
    input m_axis_bramio_87_aclk,
    input m_axis_bramio_87_aresetn,
    output m_axis_bramio_87_tlast,
    output m_axis_bramio_87_tvalid,
    output [M_AXIS_BRAMIO_87_DMWIDTH/8-1:0] m_axis_bramio_87_tkeep,
    output [M_AXIS_BRAMIO_87_DMWIDTH/8-1:0] m_axis_bramio_87_tstrb,
    output [M_AXIS_BRAMIO_87_DMWIDTH-1:0] m_axis_bramio_87_tdata,
    input m_axis_bramio_87_tready,
    //in-out BRAM AXI-Stream output interface 88
    input m_axis_bramio_88_aclk,
    input m_axis_bramio_88_aresetn,
    output m_axis_bramio_88_tlast,
    output m_axis_bramio_88_tvalid,
    output [M_AXIS_BRAMIO_88_DMWIDTH/8-1:0] m_axis_bramio_88_tkeep,
    output [M_AXIS_BRAMIO_88_DMWIDTH/8-1:0] m_axis_bramio_88_tstrb,
    output [M_AXIS_BRAMIO_88_DMWIDTH-1:0] m_axis_bramio_88_tdata,
    input m_axis_bramio_88_tready,
    //in-out BRAM AXI-Stream output interface 89
    input m_axis_bramio_89_aclk,
    input m_axis_bramio_89_aresetn,
    output m_axis_bramio_89_tlast,
    output m_axis_bramio_89_tvalid,
    output [M_AXIS_BRAMIO_89_DMWIDTH/8-1:0] m_axis_bramio_89_tkeep,
    output [M_AXIS_BRAMIO_89_DMWIDTH/8-1:0] m_axis_bramio_89_tstrb,
    output [M_AXIS_BRAMIO_89_DMWIDTH-1:0] m_axis_bramio_89_tdata,
    input m_axis_bramio_89_tready,
    //in-out BRAM AXI-Stream output interface 90
    input m_axis_bramio_90_aclk,
    input m_axis_bramio_90_aresetn,
    output m_axis_bramio_90_tlast,
    output m_axis_bramio_90_tvalid,
    output [M_AXIS_BRAMIO_90_DMWIDTH/8-1:0] m_axis_bramio_90_tkeep,
    output [M_AXIS_BRAMIO_90_DMWIDTH/8-1:0] m_axis_bramio_90_tstrb,
    output [M_AXIS_BRAMIO_90_DMWIDTH-1:0] m_axis_bramio_90_tdata,
    input m_axis_bramio_90_tready,
    //in-out BRAM AXI-Stream output interface 91
    input m_axis_bramio_91_aclk,
    input m_axis_bramio_91_aresetn,
    output m_axis_bramio_91_tlast,
    output m_axis_bramio_91_tvalid,
    output [M_AXIS_BRAMIO_91_DMWIDTH/8-1:0] m_axis_bramio_91_tkeep,
    output [M_AXIS_BRAMIO_91_DMWIDTH/8-1:0] m_axis_bramio_91_tstrb,
    output [M_AXIS_BRAMIO_91_DMWIDTH-1:0] m_axis_bramio_91_tdata,
    input m_axis_bramio_91_tready,
    //in-out BRAM AXI-Stream output interface 92
    input m_axis_bramio_92_aclk,
    input m_axis_bramio_92_aresetn,
    output m_axis_bramio_92_tlast,
    output m_axis_bramio_92_tvalid,
    output [M_AXIS_BRAMIO_92_DMWIDTH/8-1:0] m_axis_bramio_92_tkeep,
    output [M_AXIS_BRAMIO_92_DMWIDTH/8-1:0] m_axis_bramio_92_tstrb,
    output [M_AXIS_BRAMIO_92_DMWIDTH-1:0] m_axis_bramio_92_tdata,
    input m_axis_bramio_92_tready,
    //in-out BRAM AXI-Stream output interface 93
    input m_axis_bramio_93_aclk,
    input m_axis_bramio_93_aresetn,
    output m_axis_bramio_93_tlast,
    output m_axis_bramio_93_tvalid,
    output [M_AXIS_BRAMIO_93_DMWIDTH/8-1:0] m_axis_bramio_93_tkeep,
    output [M_AXIS_BRAMIO_93_DMWIDTH/8-1:0] m_axis_bramio_93_tstrb,
    output [M_AXIS_BRAMIO_93_DMWIDTH-1:0] m_axis_bramio_93_tdata,
    input m_axis_bramio_93_tready,
    //in-out BRAM AXI-Stream output interface 94
    input m_axis_bramio_94_aclk,
    input m_axis_bramio_94_aresetn,
    output m_axis_bramio_94_tlast,
    output m_axis_bramio_94_tvalid,
    output [M_AXIS_BRAMIO_94_DMWIDTH/8-1:0] m_axis_bramio_94_tkeep,
    output [M_AXIS_BRAMIO_94_DMWIDTH/8-1:0] m_axis_bramio_94_tstrb,
    output [M_AXIS_BRAMIO_94_DMWIDTH-1:0] m_axis_bramio_94_tdata,
    input m_axis_bramio_94_tready,
    //in-out BRAM AXI-Stream output interface 95
    input m_axis_bramio_95_aclk,
    input m_axis_bramio_95_aresetn,
    output m_axis_bramio_95_tlast,
    output m_axis_bramio_95_tvalid,
    output [M_AXIS_BRAMIO_95_DMWIDTH/8-1:0] m_axis_bramio_95_tkeep,
    output [M_AXIS_BRAMIO_95_DMWIDTH/8-1:0] m_axis_bramio_95_tstrb,
    output [M_AXIS_BRAMIO_95_DMWIDTH-1:0] m_axis_bramio_95_tdata,
    input m_axis_bramio_95_tready,
    //in-out BRAM AXI-Stream output interface 96
    input m_axis_bramio_96_aclk,
    input m_axis_bramio_96_aresetn,
    output m_axis_bramio_96_tlast,
    output m_axis_bramio_96_tvalid,
    output [M_AXIS_BRAMIO_96_DMWIDTH/8-1:0] m_axis_bramio_96_tkeep,
    output [M_AXIS_BRAMIO_96_DMWIDTH/8-1:0] m_axis_bramio_96_tstrb,
    output [M_AXIS_BRAMIO_96_DMWIDTH-1:0] m_axis_bramio_96_tdata,
    input m_axis_bramio_96_tready,
    //in-out BRAM AXI-Stream output interface 97
    input m_axis_bramio_97_aclk,
    input m_axis_bramio_97_aresetn,
    output m_axis_bramio_97_tlast,
    output m_axis_bramio_97_tvalid,
    output [M_AXIS_BRAMIO_97_DMWIDTH/8-1:0] m_axis_bramio_97_tkeep,
    output [M_AXIS_BRAMIO_97_DMWIDTH/8-1:0] m_axis_bramio_97_tstrb,
    output [M_AXIS_BRAMIO_97_DMWIDTH-1:0] m_axis_bramio_97_tdata,
    input m_axis_bramio_97_tready,
    //in-out BRAM AXI-Stream output interface 98
    input m_axis_bramio_98_aclk,
    input m_axis_bramio_98_aresetn,
    output m_axis_bramio_98_tlast,
    output m_axis_bramio_98_tvalid,
    output [M_AXIS_BRAMIO_98_DMWIDTH/8-1:0] m_axis_bramio_98_tkeep,
    output [M_AXIS_BRAMIO_98_DMWIDTH/8-1:0] m_axis_bramio_98_tstrb,
    output [M_AXIS_BRAMIO_98_DMWIDTH-1:0] m_axis_bramio_98_tdata,
    input m_axis_bramio_98_tready,
    //in-out BRAM AXI-Stream output interface 99
    input m_axis_bramio_99_aclk,
    input m_axis_bramio_99_aresetn,
    output m_axis_bramio_99_tlast,
    output m_axis_bramio_99_tvalid,
    output [M_AXIS_BRAMIO_99_DMWIDTH/8-1:0] m_axis_bramio_99_tkeep,
    output [M_AXIS_BRAMIO_99_DMWIDTH/8-1:0] m_axis_bramio_99_tstrb,
    output [M_AXIS_BRAMIO_99_DMWIDTH-1:0] m_axis_bramio_99_tdata,
    input m_axis_bramio_99_tready,
    //in-out BRAM AXI-Stream output interface 100
    input m_axis_bramio_100_aclk,
    input m_axis_bramio_100_aresetn,
    output m_axis_bramio_100_tlast,
    output m_axis_bramio_100_tvalid,
    output [M_AXIS_BRAMIO_100_DMWIDTH/8-1:0] m_axis_bramio_100_tkeep,
    output [M_AXIS_BRAMIO_100_DMWIDTH/8-1:0] m_axis_bramio_100_tstrb,
    output [M_AXIS_BRAMIO_100_DMWIDTH-1:0] m_axis_bramio_100_tdata,
    input m_axis_bramio_100_tready,
    //in-out BRAM AXI-Stream output interface 101
    input m_axis_bramio_101_aclk,
    input m_axis_bramio_101_aresetn,
    output m_axis_bramio_101_tlast,
    output m_axis_bramio_101_tvalid,
    output [M_AXIS_BRAMIO_101_DMWIDTH/8-1:0] m_axis_bramio_101_tkeep,
    output [M_AXIS_BRAMIO_101_DMWIDTH/8-1:0] m_axis_bramio_101_tstrb,
    output [M_AXIS_BRAMIO_101_DMWIDTH-1:0] m_axis_bramio_101_tdata,
    input m_axis_bramio_101_tready,
    //in-out BRAM AXI-Stream output interface 102
    input m_axis_bramio_102_aclk,
    input m_axis_bramio_102_aresetn,
    output m_axis_bramio_102_tlast,
    output m_axis_bramio_102_tvalid,
    output [M_AXIS_BRAMIO_102_DMWIDTH/8-1:0] m_axis_bramio_102_tkeep,
    output [M_AXIS_BRAMIO_102_DMWIDTH/8-1:0] m_axis_bramio_102_tstrb,
    output [M_AXIS_BRAMIO_102_DMWIDTH-1:0] m_axis_bramio_102_tdata,
    input m_axis_bramio_102_tready,
    //in-out BRAM AXI-Stream output interface 103
    input m_axis_bramio_103_aclk,
    input m_axis_bramio_103_aresetn,
    output m_axis_bramio_103_tlast,
    output m_axis_bramio_103_tvalid,
    output [M_AXIS_BRAMIO_103_DMWIDTH/8-1:0] m_axis_bramio_103_tkeep,
    output [M_AXIS_BRAMIO_103_DMWIDTH/8-1:0] m_axis_bramio_103_tstrb,
    output [M_AXIS_BRAMIO_103_DMWIDTH-1:0] m_axis_bramio_103_tdata,
    input m_axis_bramio_103_tready,
    //in-out BRAM AXI-Stream output interface 104
    input m_axis_bramio_104_aclk,
    input m_axis_bramio_104_aresetn,
    output m_axis_bramio_104_tlast,
    output m_axis_bramio_104_tvalid,
    output [M_AXIS_BRAMIO_104_DMWIDTH/8-1:0] m_axis_bramio_104_tkeep,
    output [M_AXIS_BRAMIO_104_DMWIDTH/8-1:0] m_axis_bramio_104_tstrb,
    output [M_AXIS_BRAMIO_104_DMWIDTH-1:0] m_axis_bramio_104_tdata,
    input m_axis_bramio_104_tready,
    //in-out BRAM AXI-Stream output interface 105
    input m_axis_bramio_105_aclk,
    input m_axis_bramio_105_aresetn,
    output m_axis_bramio_105_tlast,
    output m_axis_bramio_105_tvalid,
    output [M_AXIS_BRAMIO_105_DMWIDTH/8-1:0] m_axis_bramio_105_tkeep,
    output [M_AXIS_BRAMIO_105_DMWIDTH/8-1:0] m_axis_bramio_105_tstrb,
    output [M_AXIS_BRAMIO_105_DMWIDTH-1:0] m_axis_bramio_105_tdata,
    input m_axis_bramio_105_tready,
    //in-out BRAM AXI-Stream output interface 106
    input m_axis_bramio_106_aclk,
    input m_axis_bramio_106_aresetn,
    output m_axis_bramio_106_tlast,
    output m_axis_bramio_106_tvalid,
    output [M_AXIS_BRAMIO_106_DMWIDTH/8-1:0] m_axis_bramio_106_tkeep,
    output [M_AXIS_BRAMIO_106_DMWIDTH/8-1:0] m_axis_bramio_106_tstrb,
    output [M_AXIS_BRAMIO_106_DMWIDTH-1:0] m_axis_bramio_106_tdata,
    input m_axis_bramio_106_tready,
    //in-out BRAM AXI-Stream output interface 107
    input m_axis_bramio_107_aclk,
    input m_axis_bramio_107_aresetn,
    output m_axis_bramio_107_tlast,
    output m_axis_bramio_107_tvalid,
    output [M_AXIS_BRAMIO_107_DMWIDTH/8-1:0] m_axis_bramio_107_tkeep,
    output [M_AXIS_BRAMIO_107_DMWIDTH/8-1:0] m_axis_bramio_107_tstrb,
    output [M_AXIS_BRAMIO_107_DMWIDTH-1:0] m_axis_bramio_107_tdata,
    input m_axis_bramio_107_tready,
    //in-out BRAM AXI-Stream output interface 108
    input m_axis_bramio_108_aclk,
    input m_axis_bramio_108_aresetn,
    output m_axis_bramio_108_tlast,
    output m_axis_bramio_108_tvalid,
    output [M_AXIS_BRAMIO_108_DMWIDTH/8-1:0] m_axis_bramio_108_tkeep,
    output [M_AXIS_BRAMIO_108_DMWIDTH/8-1:0] m_axis_bramio_108_tstrb,
    output [M_AXIS_BRAMIO_108_DMWIDTH-1:0] m_axis_bramio_108_tdata,
    input m_axis_bramio_108_tready,
    //in-out BRAM AXI-Stream output interface 109
    input m_axis_bramio_109_aclk,
    input m_axis_bramio_109_aresetn,
    output m_axis_bramio_109_tlast,
    output m_axis_bramio_109_tvalid,
    output [M_AXIS_BRAMIO_109_DMWIDTH/8-1:0] m_axis_bramio_109_tkeep,
    output [M_AXIS_BRAMIO_109_DMWIDTH/8-1:0] m_axis_bramio_109_tstrb,
    output [M_AXIS_BRAMIO_109_DMWIDTH-1:0] m_axis_bramio_109_tdata,
    input m_axis_bramio_109_tready,
    //in-out BRAM AXI-Stream output interface 110
    input m_axis_bramio_110_aclk,
    input m_axis_bramio_110_aresetn,
    output m_axis_bramio_110_tlast,
    output m_axis_bramio_110_tvalid,
    output [M_AXIS_BRAMIO_110_DMWIDTH/8-1:0] m_axis_bramio_110_tkeep,
    output [M_AXIS_BRAMIO_110_DMWIDTH/8-1:0] m_axis_bramio_110_tstrb,
    output [M_AXIS_BRAMIO_110_DMWIDTH-1:0] m_axis_bramio_110_tdata,
    input m_axis_bramio_110_tready,
    //in-out BRAM AXI-Stream output interface 111
    input m_axis_bramio_111_aclk,
    input m_axis_bramio_111_aresetn,
    output m_axis_bramio_111_tlast,
    output m_axis_bramio_111_tvalid,
    output [M_AXIS_BRAMIO_111_DMWIDTH/8-1:0] m_axis_bramio_111_tkeep,
    output [M_AXIS_BRAMIO_111_DMWIDTH/8-1:0] m_axis_bramio_111_tstrb,
    output [M_AXIS_BRAMIO_111_DMWIDTH-1:0] m_axis_bramio_111_tdata,
    input m_axis_bramio_111_tready,
    //in-out BRAM AXI-Stream output interface 112
    input m_axis_bramio_112_aclk,
    input m_axis_bramio_112_aresetn,
    output m_axis_bramio_112_tlast,
    output m_axis_bramio_112_tvalid,
    output [M_AXIS_BRAMIO_112_DMWIDTH/8-1:0] m_axis_bramio_112_tkeep,
    output [M_AXIS_BRAMIO_112_DMWIDTH/8-1:0] m_axis_bramio_112_tstrb,
    output [M_AXIS_BRAMIO_112_DMWIDTH-1:0] m_axis_bramio_112_tdata,
    input m_axis_bramio_112_tready,
    //in-out BRAM AXI-Stream output interface 113
    input m_axis_bramio_113_aclk,
    input m_axis_bramio_113_aresetn,
    output m_axis_bramio_113_tlast,
    output m_axis_bramio_113_tvalid,
    output [M_AXIS_BRAMIO_113_DMWIDTH/8-1:0] m_axis_bramio_113_tkeep,
    output [M_AXIS_BRAMIO_113_DMWIDTH/8-1:0] m_axis_bramio_113_tstrb,
    output [M_AXIS_BRAMIO_113_DMWIDTH-1:0] m_axis_bramio_113_tdata,
    input m_axis_bramio_113_tready,
    //in-out BRAM AXI-Stream output interface 114
    input m_axis_bramio_114_aclk,
    input m_axis_bramio_114_aresetn,
    output m_axis_bramio_114_tlast,
    output m_axis_bramio_114_tvalid,
    output [M_AXIS_BRAMIO_114_DMWIDTH/8-1:0] m_axis_bramio_114_tkeep,
    output [M_AXIS_BRAMIO_114_DMWIDTH/8-1:0] m_axis_bramio_114_tstrb,
    output [M_AXIS_BRAMIO_114_DMWIDTH-1:0] m_axis_bramio_114_tdata,
    input m_axis_bramio_114_tready,
    //in-out BRAM AXI-Stream output interface 115
    input m_axis_bramio_115_aclk,
    input m_axis_bramio_115_aresetn,
    output m_axis_bramio_115_tlast,
    output m_axis_bramio_115_tvalid,
    output [M_AXIS_BRAMIO_115_DMWIDTH/8-1:0] m_axis_bramio_115_tkeep,
    output [M_AXIS_BRAMIO_115_DMWIDTH/8-1:0] m_axis_bramio_115_tstrb,
    output [M_AXIS_BRAMIO_115_DMWIDTH-1:0] m_axis_bramio_115_tdata,
    input m_axis_bramio_115_tready,
    //in-out BRAM AXI-Stream output interface 116
    input m_axis_bramio_116_aclk,
    input m_axis_bramio_116_aresetn,
    output m_axis_bramio_116_tlast,
    output m_axis_bramio_116_tvalid,
    output [M_AXIS_BRAMIO_116_DMWIDTH/8-1:0] m_axis_bramio_116_tkeep,
    output [M_AXIS_BRAMIO_116_DMWIDTH/8-1:0] m_axis_bramio_116_tstrb,
    output [M_AXIS_BRAMIO_116_DMWIDTH-1:0] m_axis_bramio_116_tdata,
    input m_axis_bramio_116_tready,
    //in-out BRAM AXI-Stream output interface 117
    input m_axis_bramio_117_aclk,
    input m_axis_bramio_117_aresetn,
    output m_axis_bramio_117_tlast,
    output m_axis_bramio_117_tvalid,
    output [M_AXIS_BRAMIO_117_DMWIDTH/8-1:0] m_axis_bramio_117_tkeep,
    output [M_AXIS_BRAMIO_117_DMWIDTH/8-1:0] m_axis_bramio_117_tstrb,
    output [M_AXIS_BRAMIO_117_DMWIDTH-1:0] m_axis_bramio_117_tdata,
    input m_axis_bramio_117_tready,
    //in-out BRAM AXI-Stream output interface 118
    input m_axis_bramio_118_aclk,
    input m_axis_bramio_118_aresetn,
    output m_axis_bramio_118_tlast,
    output m_axis_bramio_118_tvalid,
    output [M_AXIS_BRAMIO_118_DMWIDTH/8-1:0] m_axis_bramio_118_tkeep,
    output [M_AXIS_BRAMIO_118_DMWIDTH/8-1:0] m_axis_bramio_118_tstrb,
    output [M_AXIS_BRAMIO_118_DMWIDTH-1:0] m_axis_bramio_118_tdata,
    input m_axis_bramio_118_tready,
    //in-out BRAM AXI-Stream output interface 119
    input m_axis_bramio_119_aclk,
    input m_axis_bramio_119_aresetn,
    output m_axis_bramio_119_tlast,
    output m_axis_bramio_119_tvalid,
    output [M_AXIS_BRAMIO_119_DMWIDTH/8-1:0] m_axis_bramio_119_tkeep,
    output [M_AXIS_BRAMIO_119_DMWIDTH/8-1:0] m_axis_bramio_119_tstrb,
    output [M_AXIS_BRAMIO_119_DMWIDTH-1:0] m_axis_bramio_119_tdata,
    input m_axis_bramio_119_tready,
    //in-out BRAM AXI-Stream output interface 120
    input m_axis_bramio_120_aclk,
    input m_axis_bramio_120_aresetn,
    output m_axis_bramio_120_tlast,
    output m_axis_bramio_120_tvalid,
    output [M_AXIS_BRAMIO_120_DMWIDTH/8-1:0] m_axis_bramio_120_tkeep,
    output [M_AXIS_BRAMIO_120_DMWIDTH/8-1:0] m_axis_bramio_120_tstrb,
    output [M_AXIS_BRAMIO_120_DMWIDTH-1:0] m_axis_bramio_120_tdata,
    input m_axis_bramio_120_tready,
    //in-out BRAM AXI-Stream output interface 121
    input m_axis_bramio_121_aclk,
    input m_axis_bramio_121_aresetn,
    output m_axis_bramio_121_tlast,
    output m_axis_bramio_121_tvalid,
    output [M_AXIS_BRAMIO_121_DMWIDTH/8-1:0] m_axis_bramio_121_tkeep,
    output [M_AXIS_BRAMIO_121_DMWIDTH/8-1:0] m_axis_bramio_121_tstrb,
    output [M_AXIS_BRAMIO_121_DMWIDTH-1:0] m_axis_bramio_121_tdata,
    input m_axis_bramio_121_tready,
    //in-out BRAM AXI-Stream output interface 122
    input m_axis_bramio_122_aclk,
    input m_axis_bramio_122_aresetn,
    output m_axis_bramio_122_tlast,
    output m_axis_bramio_122_tvalid,
    output [M_AXIS_BRAMIO_122_DMWIDTH/8-1:0] m_axis_bramio_122_tkeep,
    output [M_AXIS_BRAMIO_122_DMWIDTH/8-1:0] m_axis_bramio_122_tstrb,
    output [M_AXIS_BRAMIO_122_DMWIDTH-1:0] m_axis_bramio_122_tdata,
    input m_axis_bramio_122_tready,
    //in-out BRAM AXI-Stream output interface 123
    input m_axis_bramio_123_aclk,
    input m_axis_bramio_123_aresetn,
    output m_axis_bramio_123_tlast,
    output m_axis_bramio_123_tvalid,
    output [M_AXIS_BRAMIO_123_DMWIDTH/8-1:0] m_axis_bramio_123_tkeep,
    output [M_AXIS_BRAMIO_123_DMWIDTH/8-1:0] m_axis_bramio_123_tstrb,
    output [M_AXIS_BRAMIO_123_DMWIDTH-1:0] m_axis_bramio_123_tdata,
    input m_axis_bramio_123_tready,
    //in-out BRAM AXI-Stream output interface 124
    input m_axis_bramio_124_aclk,
    input m_axis_bramio_124_aresetn,
    output m_axis_bramio_124_tlast,
    output m_axis_bramio_124_tvalid,
    output [M_AXIS_BRAMIO_124_DMWIDTH/8-1:0] m_axis_bramio_124_tkeep,
    output [M_AXIS_BRAMIO_124_DMWIDTH/8-1:0] m_axis_bramio_124_tstrb,
    output [M_AXIS_BRAMIO_124_DMWIDTH-1:0] m_axis_bramio_124_tdata,
    input m_axis_bramio_124_tready,
    //in-out BRAM AXI-Stream output interface 125
    input m_axis_bramio_125_aclk,
    input m_axis_bramio_125_aresetn,
    output m_axis_bramio_125_tlast,
    output m_axis_bramio_125_tvalid,
    output [M_AXIS_BRAMIO_125_DMWIDTH/8-1:0] m_axis_bramio_125_tkeep,
    output [M_AXIS_BRAMIO_125_DMWIDTH/8-1:0] m_axis_bramio_125_tstrb,
    output [M_AXIS_BRAMIO_125_DMWIDTH-1:0] m_axis_bramio_125_tdata,
    input m_axis_bramio_125_tready,
    //in-out BRAM AXI-Stream output interface 126
    input m_axis_bramio_126_aclk,
    input m_axis_bramio_126_aresetn,
    output m_axis_bramio_126_tlast,
    output m_axis_bramio_126_tvalid,
    output [M_AXIS_BRAMIO_126_DMWIDTH/8-1:0] m_axis_bramio_126_tkeep,
    output [M_AXIS_BRAMIO_126_DMWIDTH/8-1:0] m_axis_bramio_126_tstrb,
    output [M_AXIS_BRAMIO_126_DMWIDTH-1:0] m_axis_bramio_126_tdata,
    input m_axis_bramio_126_tready,
    //in-out BRAM AXI-Stream output interface 127
    input m_axis_bramio_127_aclk,
    input m_axis_bramio_127_aresetn,
    output m_axis_bramio_127_tlast,
    output m_axis_bramio_127_tvalid,
    output [M_AXIS_BRAMIO_127_DMWIDTH/8-1:0] m_axis_bramio_127_tkeep,
    output [M_AXIS_BRAMIO_127_DMWIDTH/8-1:0] m_axis_bramio_127_tstrb,
    output [M_AXIS_BRAMIO_127_DMWIDTH-1:0] m_axis_bramio_127_tdata,
    input m_axis_bramio_127_tready,
    //-----------------------------------------------------------
    //out BRAM to AXI-Stream interface 0
    input m_axis_bram_0_aclk,
    input m_axis_bram_0_aresetn,
    output m_axis_bram_0_tlast,
    output m_axis_bram_0_tvalid,
    output [M_AXIS_BRAM_0_DMWIDTH/8-1:0] m_axis_bram_0_tkeep,
    output [M_AXIS_BRAM_0_DMWIDTH/8-1:0] m_axis_bram_0_tstrb,
    output [M_AXIS_BRAM_0_DMWIDTH-1:0] m_axis_bram_0_tdata,
    input m_axis_bram_0_tready,
    input [M_AXIS_BRAM_0_ADDR_WIDTH-1:0] ap_bram_oarg_0_addr0,
    input [M_AXIS_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_din0,
    output [M_AXIS_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_dout0,
    input ap_bram_oarg_0_clk0,
    input ap_bram_oarg_0_rst0,
    input [M_AXIS_BRAM_0_WIDTH/8-1:0] ap_bram_oarg_0_we0,
    input ap_bram_oarg_0_en0,
    input [M_AXIS_BRAM_0_ADDR_WIDTH-1:0] ap_bram_oarg_0_addr1,
    input [M_AXIS_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_din1,
    output [M_AXIS_BRAM_0_WIDTH-1:0] ap_bram_oarg_0_dout1,
    input ap_bram_oarg_0_clk1,
    input ap_bram_oarg_0_rst1,
    input [M_AXIS_BRAM_0_WIDTH/8-1:0] ap_bram_oarg_0_we1,
    input ap_bram_oarg_0_en1,
    //out BRAM to AXI-Stream interface 1
    input m_axis_bram_1_aclk,
    input m_axis_bram_1_aresetn,
    output m_axis_bram_1_tlast,
    output m_axis_bram_1_tvalid,
    output [M_AXIS_BRAM_1_DMWIDTH/8-1:0] m_axis_bram_1_tkeep,
    output [M_AXIS_BRAM_1_DMWIDTH/8-1:0] m_axis_bram_1_tstrb,
    output [M_AXIS_BRAM_1_DMWIDTH-1:0] m_axis_bram_1_tdata,
    input m_axis_bram_1_tready,
    input [M_AXIS_BRAM_1_ADDR_WIDTH-1:0] ap_bram_oarg_1_addr0,
    input [M_AXIS_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_din0,
    output [M_AXIS_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_dout0,
    input ap_bram_oarg_1_clk0,
    input ap_bram_oarg_1_rst0,
    input [M_AXIS_BRAM_1_WIDTH/8-1:0] ap_bram_oarg_1_we0,
    input ap_bram_oarg_1_en0,
    input [M_AXIS_BRAM_1_ADDR_WIDTH-1:0] ap_bram_oarg_1_addr1,
    input [M_AXIS_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_din1,
    output [M_AXIS_BRAM_1_WIDTH-1:0] ap_bram_oarg_1_dout1,
    input ap_bram_oarg_1_clk1,
    input ap_bram_oarg_1_rst1,
    input [M_AXIS_BRAM_1_WIDTH/8-1:0] ap_bram_oarg_1_we1,
    input ap_bram_oarg_1_en1,
    //out BRAM to AXI-Stream interface 2
    input m_axis_bram_2_aclk,
    input m_axis_bram_2_aresetn,
    output m_axis_bram_2_tlast,
    output m_axis_bram_2_tvalid,
    output [M_AXIS_BRAM_2_DMWIDTH/8-1:0] m_axis_bram_2_tkeep,
    output [M_AXIS_BRAM_2_DMWIDTH/8-1:0] m_axis_bram_2_tstrb,
    output [M_AXIS_BRAM_2_DMWIDTH-1:0] m_axis_bram_2_tdata,
    input m_axis_bram_2_tready,
    input [M_AXIS_BRAM_2_ADDR_WIDTH-1:0] ap_bram_oarg_2_addr0,
    input [M_AXIS_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_din0,
    output [M_AXIS_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_dout0,
    input ap_bram_oarg_2_clk0,
    input ap_bram_oarg_2_rst0,
    input [M_AXIS_BRAM_2_WIDTH/8-1:0] ap_bram_oarg_2_we0,
    input ap_bram_oarg_2_en0,
    input [M_AXIS_BRAM_2_ADDR_WIDTH-1:0] ap_bram_oarg_2_addr1,
    input [M_AXIS_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_din1,
    output [M_AXIS_BRAM_2_WIDTH-1:0] ap_bram_oarg_2_dout1,
    input ap_bram_oarg_2_clk1,
    input ap_bram_oarg_2_rst1,
    input [M_AXIS_BRAM_2_WIDTH/8-1:0] ap_bram_oarg_2_we1,
    input ap_bram_oarg_2_en1,
    //out BRAM to AXI-Stream interface 3
    input m_axis_bram_3_aclk,
    input m_axis_bram_3_aresetn,
    output m_axis_bram_3_tlast,
    output m_axis_bram_3_tvalid,
    output [M_AXIS_BRAM_3_DMWIDTH/8-1:0] m_axis_bram_3_tkeep,
    output [M_AXIS_BRAM_3_DMWIDTH/8-1:0] m_axis_bram_3_tstrb,
    output [M_AXIS_BRAM_3_DMWIDTH-1:0] m_axis_bram_3_tdata,
    input m_axis_bram_3_tready,
    input [M_AXIS_BRAM_3_ADDR_WIDTH-1:0] ap_bram_oarg_3_addr0,
    input [M_AXIS_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_din0,
    output [M_AXIS_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_dout0,
    input ap_bram_oarg_3_clk0,
    input ap_bram_oarg_3_rst0,
    input [M_AXIS_BRAM_3_WIDTH/8-1:0] ap_bram_oarg_3_we0,
    input ap_bram_oarg_3_en0,
    input [M_AXIS_BRAM_3_ADDR_WIDTH-1:0] ap_bram_oarg_3_addr1,
    input [M_AXIS_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_din1,
    output [M_AXIS_BRAM_3_WIDTH-1:0] ap_bram_oarg_3_dout1,
    input ap_bram_oarg_3_clk1,
    input ap_bram_oarg_3_rst1,
    input [M_AXIS_BRAM_3_WIDTH/8-1:0] ap_bram_oarg_3_we1,
    input ap_bram_oarg_3_en1,
    //out BRAM to AXI-Stream interface 4
    input m_axis_bram_4_aclk,
    input m_axis_bram_4_aresetn,
    output m_axis_bram_4_tlast,
    output m_axis_bram_4_tvalid,
    output [M_AXIS_BRAM_4_DMWIDTH/8-1:0] m_axis_bram_4_tkeep,
    output [M_AXIS_BRAM_4_DMWIDTH/8-1:0] m_axis_bram_4_tstrb,
    output [M_AXIS_BRAM_4_DMWIDTH-1:0] m_axis_bram_4_tdata,
    input m_axis_bram_4_tready,
    input [M_AXIS_BRAM_4_ADDR_WIDTH-1:0] ap_bram_oarg_4_addr0,
    input [M_AXIS_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_din0,
    output [M_AXIS_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_dout0,
    input ap_bram_oarg_4_clk0,
    input ap_bram_oarg_4_rst0,
    input [M_AXIS_BRAM_4_WIDTH/8-1:0] ap_bram_oarg_4_we0,
    input ap_bram_oarg_4_en0,
    input [M_AXIS_BRAM_4_ADDR_WIDTH-1:0] ap_bram_oarg_4_addr1,
    input [M_AXIS_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_din1,
    output [M_AXIS_BRAM_4_WIDTH-1:0] ap_bram_oarg_4_dout1,
    input ap_bram_oarg_4_clk1,
    input ap_bram_oarg_4_rst1,
    input [M_AXIS_BRAM_4_WIDTH/8-1:0] ap_bram_oarg_4_we1,
    input ap_bram_oarg_4_en1,
    //out BRAM to AXI-Stream interface 5
    input m_axis_bram_5_aclk,
    input m_axis_bram_5_aresetn,
    output m_axis_bram_5_tlast,
    output m_axis_bram_5_tvalid,
    output [M_AXIS_BRAM_5_DMWIDTH/8-1:0] m_axis_bram_5_tkeep,
    output [M_AXIS_BRAM_5_DMWIDTH/8-1:0] m_axis_bram_5_tstrb,
    output [M_AXIS_BRAM_5_DMWIDTH-1:0] m_axis_bram_5_tdata,
    input m_axis_bram_5_tready,
    input [M_AXIS_BRAM_5_ADDR_WIDTH-1:0] ap_bram_oarg_5_addr0,
    input [M_AXIS_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_din0,
    output [M_AXIS_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_dout0,
    input ap_bram_oarg_5_clk0,
    input ap_bram_oarg_5_rst0,
    input [M_AXIS_BRAM_5_WIDTH/8-1:0] ap_bram_oarg_5_we0,
    input ap_bram_oarg_5_en0,
    input [M_AXIS_BRAM_5_ADDR_WIDTH-1:0] ap_bram_oarg_5_addr1,
    input [M_AXIS_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_din1,
    output [M_AXIS_BRAM_5_WIDTH-1:0] ap_bram_oarg_5_dout1,
    input ap_bram_oarg_5_clk1,
    input ap_bram_oarg_5_rst1,
    input [M_AXIS_BRAM_5_WIDTH/8-1:0] ap_bram_oarg_5_we1,
    input ap_bram_oarg_5_en1,
    //out BRAM to AXI-Stream interface 6
    input m_axis_bram_6_aclk,
    input m_axis_bram_6_aresetn,
    output m_axis_bram_6_tlast,
    output m_axis_bram_6_tvalid,
    output [M_AXIS_BRAM_6_DMWIDTH/8-1:0] m_axis_bram_6_tkeep,
    output [M_AXIS_BRAM_6_DMWIDTH/8-1:0] m_axis_bram_6_tstrb,
    output [M_AXIS_BRAM_6_DMWIDTH-1:0] m_axis_bram_6_tdata,
    input m_axis_bram_6_tready,
    input [M_AXIS_BRAM_6_ADDR_WIDTH-1:0] ap_bram_oarg_6_addr0,
    input [M_AXIS_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_din0,
    output [M_AXIS_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_dout0,
    input ap_bram_oarg_6_clk0,
    input ap_bram_oarg_6_rst0,
    input [M_AXIS_BRAM_6_WIDTH/8-1:0] ap_bram_oarg_6_we0,
    input ap_bram_oarg_6_en0,
    input [M_AXIS_BRAM_6_ADDR_WIDTH-1:0] ap_bram_oarg_6_addr1,
    input [M_AXIS_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_din1,
    output [M_AXIS_BRAM_6_WIDTH-1:0] ap_bram_oarg_6_dout1,
    input ap_bram_oarg_6_clk1,
    input ap_bram_oarg_6_rst1,
    input [M_AXIS_BRAM_6_WIDTH/8-1:0] ap_bram_oarg_6_we1,
    input ap_bram_oarg_6_en1,
    //out BRAM to AXI-Stream interface 7
    input m_axis_bram_7_aclk,
    input m_axis_bram_7_aresetn,
    output m_axis_bram_7_tlast,
    output m_axis_bram_7_tvalid,
    output [M_AXIS_BRAM_7_DMWIDTH/8-1:0] m_axis_bram_7_tkeep,
    output [M_AXIS_BRAM_7_DMWIDTH/8-1:0] m_axis_bram_7_tstrb,
    output [M_AXIS_BRAM_7_DMWIDTH-1:0] m_axis_bram_7_tdata,
    input m_axis_bram_7_tready,
    input [M_AXIS_BRAM_7_ADDR_WIDTH-1:0] ap_bram_oarg_7_addr0,
    input [M_AXIS_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_din0,
    output [M_AXIS_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_dout0,
    input ap_bram_oarg_7_clk0,
    input ap_bram_oarg_7_rst0,
    input [M_AXIS_BRAM_7_WIDTH/8-1:0] ap_bram_oarg_7_we0,
    input ap_bram_oarg_7_en0,
    input [M_AXIS_BRAM_7_ADDR_WIDTH-1:0] ap_bram_oarg_7_addr1,
    input [M_AXIS_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_din1,
    output [M_AXIS_BRAM_7_WIDTH-1:0] ap_bram_oarg_7_dout1,
    input ap_bram_oarg_7_clk1,
    input ap_bram_oarg_7_rst1,
    input [M_AXIS_BRAM_7_WIDTH/8-1:0] ap_bram_oarg_7_we1,
    input ap_bram_oarg_7_en1,
    //out BRAM to AXI-Stream interface 8
    input m_axis_bram_8_aclk,
    input m_axis_bram_8_aresetn,
    output m_axis_bram_8_tlast,
    output m_axis_bram_8_tvalid,
    output [M_AXIS_BRAM_8_DMWIDTH/8-1:0] m_axis_bram_8_tkeep,
    output [M_AXIS_BRAM_8_DMWIDTH/8-1:0] m_axis_bram_8_tstrb,
    output [M_AXIS_BRAM_8_DMWIDTH-1:0] m_axis_bram_8_tdata,
    input m_axis_bram_8_tready,
    input [M_AXIS_BRAM_8_ADDR_WIDTH-1:0] ap_bram_oarg_8_addr0,
    input [M_AXIS_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_din0,
    output [M_AXIS_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_dout0,
    input ap_bram_oarg_8_clk0,
    input ap_bram_oarg_8_rst0,
    input [M_AXIS_BRAM_8_WIDTH/8-1:0] ap_bram_oarg_8_we0,
    input ap_bram_oarg_8_en0,
    input [M_AXIS_BRAM_8_ADDR_WIDTH-1:0] ap_bram_oarg_8_addr1,
    input [M_AXIS_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_din1,
    output [M_AXIS_BRAM_8_WIDTH-1:0] ap_bram_oarg_8_dout1,
    input ap_bram_oarg_8_clk1,
    input ap_bram_oarg_8_rst1,
    input [M_AXIS_BRAM_8_WIDTH/8-1:0] ap_bram_oarg_8_we1,
    input ap_bram_oarg_8_en1,
    //out BRAM to AXI-Stream interface 9
    input m_axis_bram_9_aclk,
    input m_axis_bram_9_aresetn,
    output m_axis_bram_9_tlast,
    output m_axis_bram_9_tvalid,
    output [M_AXIS_BRAM_9_DMWIDTH/8-1:0] m_axis_bram_9_tkeep,
    output [M_AXIS_BRAM_9_DMWIDTH/8-1:0] m_axis_bram_9_tstrb,
    output [M_AXIS_BRAM_9_DMWIDTH-1:0] m_axis_bram_9_tdata,
    input m_axis_bram_9_tready,
    input [M_AXIS_BRAM_9_ADDR_WIDTH-1:0] ap_bram_oarg_9_addr0,
    input [M_AXIS_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_din0,
    output [M_AXIS_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_dout0,
    input ap_bram_oarg_9_clk0,
    input ap_bram_oarg_9_rst0,
    input [M_AXIS_BRAM_9_WIDTH/8-1:0] ap_bram_oarg_9_we0,
    input ap_bram_oarg_9_en0,
    input [M_AXIS_BRAM_9_ADDR_WIDTH-1:0] ap_bram_oarg_9_addr1,
    input [M_AXIS_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_din1,
    output [M_AXIS_BRAM_9_WIDTH-1:0] ap_bram_oarg_9_dout1,
    input ap_bram_oarg_9_clk1,
    input ap_bram_oarg_9_rst1,
    input [M_AXIS_BRAM_9_WIDTH/8-1:0] ap_bram_oarg_9_we1,
    input ap_bram_oarg_9_en1,
    //out BRAM to AXI-Stream interface 10
    input m_axis_bram_10_aclk,
    input m_axis_bram_10_aresetn,
    output m_axis_bram_10_tlast,
    output m_axis_bram_10_tvalid,
    output [M_AXIS_BRAM_10_DMWIDTH/8-1:0] m_axis_bram_10_tkeep,
    output [M_AXIS_BRAM_10_DMWIDTH/8-1:0] m_axis_bram_10_tstrb,
    output [M_AXIS_BRAM_10_DMWIDTH-1:0] m_axis_bram_10_tdata,
    input m_axis_bram_10_tready,
    input [M_AXIS_BRAM_10_ADDR_WIDTH-1:0] ap_bram_oarg_10_addr0,
    input [M_AXIS_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_din0,
    output [M_AXIS_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_dout0,
    input ap_bram_oarg_10_clk0,
    input ap_bram_oarg_10_rst0,
    input [M_AXIS_BRAM_10_WIDTH/8-1:0] ap_bram_oarg_10_we0,
    input ap_bram_oarg_10_en0,
    input [M_AXIS_BRAM_10_ADDR_WIDTH-1:0] ap_bram_oarg_10_addr1,
    input [M_AXIS_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_din1,
    output [M_AXIS_BRAM_10_WIDTH-1:0] ap_bram_oarg_10_dout1,
    input ap_bram_oarg_10_clk1,
    input ap_bram_oarg_10_rst1,
    input [M_AXIS_BRAM_10_WIDTH/8-1:0] ap_bram_oarg_10_we1,
    input ap_bram_oarg_10_en1,
    //out BRAM to AXI-Stream interface 11
    input m_axis_bram_11_aclk,
    input m_axis_bram_11_aresetn,
    output m_axis_bram_11_tlast,
    output m_axis_bram_11_tvalid,
    output [M_AXIS_BRAM_11_DMWIDTH/8-1:0] m_axis_bram_11_tkeep,
    output [M_AXIS_BRAM_11_DMWIDTH/8-1:0] m_axis_bram_11_tstrb,
    output [M_AXIS_BRAM_11_DMWIDTH-1:0] m_axis_bram_11_tdata,
    input m_axis_bram_11_tready,
    input [M_AXIS_BRAM_11_ADDR_WIDTH-1:0] ap_bram_oarg_11_addr0,
    input [M_AXIS_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_din0,
    output [M_AXIS_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_dout0,
    input ap_bram_oarg_11_clk0,
    input ap_bram_oarg_11_rst0,
    input [M_AXIS_BRAM_11_WIDTH/8-1:0] ap_bram_oarg_11_we0,
    input ap_bram_oarg_11_en0,
    input [M_AXIS_BRAM_11_ADDR_WIDTH-1:0] ap_bram_oarg_11_addr1,
    input [M_AXIS_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_din1,
    output [M_AXIS_BRAM_11_WIDTH-1:0] ap_bram_oarg_11_dout1,
    input ap_bram_oarg_11_clk1,
    input ap_bram_oarg_11_rst1,
    input [M_AXIS_BRAM_11_WIDTH/8-1:0] ap_bram_oarg_11_we1,
    input ap_bram_oarg_11_en1,
    //out BRAM to AXI-Stream interface 12
    input m_axis_bram_12_aclk,
    input m_axis_bram_12_aresetn,
    output m_axis_bram_12_tlast,
    output m_axis_bram_12_tvalid,
    output [M_AXIS_BRAM_12_DMWIDTH/8-1:0] m_axis_bram_12_tkeep,
    output [M_AXIS_BRAM_12_DMWIDTH/8-1:0] m_axis_bram_12_tstrb,
    output [M_AXIS_BRAM_12_DMWIDTH-1:0] m_axis_bram_12_tdata,
    input m_axis_bram_12_tready,
    input [M_AXIS_BRAM_12_ADDR_WIDTH-1:0] ap_bram_oarg_12_addr0,
    input [M_AXIS_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_din0,
    output [M_AXIS_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_dout0,
    input ap_bram_oarg_12_clk0,
    input ap_bram_oarg_12_rst0,
    input [M_AXIS_BRAM_12_WIDTH/8-1:0] ap_bram_oarg_12_we0,
    input ap_bram_oarg_12_en0,
    input [M_AXIS_BRAM_12_ADDR_WIDTH-1:0] ap_bram_oarg_12_addr1,
    input [M_AXIS_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_din1,
    output [M_AXIS_BRAM_12_WIDTH-1:0] ap_bram_oarg_12_dout1,
    input ap_bram_oarg_12_clk1,
    input ap_bram_oarg_12_rst1,
    input [M_AXIS_BRAM_12_WIDTH/8-1:0] ap_bram_oarg_12_we1,
    input ap_bram_oarg_12_en1,
    //out BRAM to AXI-Stream interface 13
    input m_axis_bram_13_aclk,
    input m_axis_bram_13_aresetn,
    output m_axis_bram_13_tlast,
    output m_axis_bram_13_tvalid,
    output [M_AXIS_BRAM_13_DMWIDTH/8-1:0] m_axis_bram_13_tkeep,
    output [M_AXIS_BRAM_13_DMWIDTH/8-1:0] m_axis_bram_13_tstrb,
    output [M_AXIS_BRAM_13_DMWIDTH-1:0] m_axis_bram_13_tdata,
    input m_axis_bram_13_tready,
    input [M_AXIS_BRAM_13_ADDR_WIDTH-1:0] ap_bram_oarg_13_addr0,
    input [M_AXIS_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_din0,
    output [M_AXIS_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_dout0,
    input ap_bram_oarg_13_clk0,
    input ap_bram_oarg_13_rst0,
    input [M_AXIS_BRAM_13_WIDTH/8-1:0] ap_bram_oarg_13_we0,
    input ap_bram_oarg_13_en0,
    input [M_AXIS_BRAM_13_ADDR_WIDTH-1:0] ap_bram_oarg_13_addr1,
    input [M_AXIS_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_din1,
    output [M_AXIS_BRAM_13_WIDTH-1:0] ap_bram_oarg_13_dout1,
    input ap_bram_oarg_13_clk1,
    input ap_bram_oarg_13_rst1,
    input [M_AXIS_BRAM_13_WIDTH/8-1:0] ap_bram_oarg_13_we1,
    input ap_bram_oarg_13_en1,
    //out BRAM to AXI-Stream interface 14
    input m_axis_bram_14_aclk,
    input m_axis_bram_14_aresetn,
    output m_axis_bram_14_tlast,
    output m_axis_bram_14_tvalid,
    output [M_AXIS_BRAM_14_DMWIDTH/8-1:0] m_axis_bram_14_tkeep,
    output [M_AXIS_BRAM_14_DMWIDTH/8-1:0] m_axis_bram_14_tstrb,
    output [M_AXIS_BRAM_14_DMWIDTH-1:0] m_axis_bram_14_tdata,
    input m_axis_bram_14_tready,
    input [M_AXIS_BRAM_14_ADDR_WIDTH-1:0] ap_bram_oarg_14_addr0,
    input [M_AXIS_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_din0,
    output [M_AXIS_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_dout0,
    input ap_bram_oarg_14_clk0,
    input ap_bram_oarg_14_rst0,
    input [M_AXIS_BRAM_14_WIDTH/8-1:0] ap_bram_oarg_14_we0,
    input ap_bram_oarg_14_en0,
    input [M_AXIS_BRAM_14_ADDR_WIDTH-1:0] ap_bram_oarg_14_addr1,
    input [M_AXIS_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_din1,
    output [M_AXIS_BRAM_14_WIDTH-1:0] ap_bram_oarg_14_dout1,
    input ap_bram_oarg_14_clk1,
    input ap_bram_oarg_14_rst1,
    input [M_AXIS_BRAM_14_WIDTH/8-1:0] ap_bram_oarg_14_we1,
    input ap_bram_oarg_14_en1,
    //out BRAM to AXI-Stream interface 15
    input m_axis_bram_15_aclk,
    input m_axis_bram_15_aresetn,
    output m_axis_bram_15_tlast,
    output m_axis_bram_15_tvalid,
    output [M_AXIS_BRAM_15_DMWIDTH/8-1:0] m_axis_bram_15_tkeep,
    output [M_AXIS_BRAM_15_DMWIDTH/8-1:0] m_axis_bram_15_tstrb,
    output [M_AXIS_BRAM_15_DMWIDTH-1:0] m_axis_bram_15_tdata,
    input m_axis_bram_15_tready,
    input [M_AXIS_BRAM_15_ADDR_WIDTH-1:0] ap_bram_oarg_15_addr0,
    input [M_AXIS_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_din0,
    output [M_AXIS_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_dout0,
    input ap_bram_oarg_15_clk0,
    input ap_bram_oarg_15_rst0,
    input [M_AXIS_BRAM_15_WIDTH/8-1:0] ap_bram_oarg_15_we0,
    input ap_bram_oarg_15_en0,
    input [M_AXIS_BRAM_15_ADDR_WIDTH-1:0] ap_bram_oarg_15_addr1,
    input [M_AXIS_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_din1,
    output [M_AXIS_BRAM_15_WIDTH-1:0] ap_bram_oarg_15_dout1,
    input ap_bram_oarg_15_clk1,
    input ap_bram_oarg_15_rst1,
    input [M_AXIS_BRAM_15_WIDTH/8-1:0] ap_bram_oarg_15_we1,
    input ap_bram_oarg_15_en1,
    //out BRAM to AXI-Stream interface 16
    input m_axis_bram_16_aclk,
    input m_axis_bram_16_aresetn,
    output m_axis_bram_16_tlast,
    output m_axis_bram_16_tvalid,
    output [M_AXIS_BRAM_16_DMWIDTH/8-1:0] m_axis_bram_16_tkeep,
    output [M_AXIS_BRAM_16_DMWIDTH/8-1:0] m_axis_bram_16_tstrb,
    output [M_AXIS_BRAM_16_DMWIDTH-1:0] m_axis_bram_16_tdata,
    input m_axis_bram_16_tready,
    input [M_AXIS_BRAM_16_ADDR_WIDTH-1:0] ap_bram_oarg_16_addr0,
    input [M_AXIS_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_din0,
    output [M_AXIS_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_dout0,
    input ap_bram_oarg_16_clk0,
    input ap_bram_oarg_16_rst0,
    input [M_AXIS_BRAM_16_WIDTH/8-1:0] ap_bram_oarg_16_we0,
    input ap_bram_oarg_16_en0,
    input [M_AXIS_BRAM_16_ADDR_WIDTH-1:0] ap_bram_oarg_16_addr1,
    input [M_AXIS_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_din1,
    output [M_AXIS_BRAM_16_WIDTH-1:0] ap_bram_oarg_16_dout1,
    input ap_bram_oarg_16_clk1,
    input ap_bram_oarg_16_rst1,
    input [M_AXIS_BRAM_16_WIDTH/8-1:0] ap_bram_oarg_16_we1,
    input ap_bram_oarg_16_en1,
    //out BRAM to AXI-Stream interface 17
    input m_axis_bram_17_aclk,
    input m_axis_bram_17_aresetn,
    output m_axis_bram_17_tlast,
    output m_axis_bram_17_tvalid,
    output [M_AXIS_BRAM_17_DMWIDTH/8-1:0] m_axis_bram_17_tkeep,
    output [M_AXIS_BRAM_17_DMWIDTH/8-1:0] m_axis_bram_17_tstrb,
    output [M_AXIS_BRAM_17_DMWIDTH-1:0] m_axis_bram_17_tdata,
    input m_axis_bram_17_tready,
    input [M_AXIS_BRAM_17_ADDR_WIDTH-1:0] ap_bram_oarg_17_addr0,
    input [M_AXIS_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_din0,
    output [M_AXIS_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_dout0,
    input ap_bram_oarg_17_clk0,
    input ap_bram_oarg_17_rst0,
    input [M_AXIS_BRAM_17_WIDTH/8-1:0] ap_bram_oarg_17_we0,
    input ap_bram_oarg_17_en0,
    input [M_AXIS_BRAM_17_ADDR_WIDTH-1:0] ap_bram_oarg_17_addr1,
    input [M_AXIS_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_din1,
    output [M_AXIS_BRAM_17_WIDTH-1:0] ap_bram_oarg_17_dout1,
    input ap_bram_oarg_17_clk1,
    input ap_bram_oarg_17_rst1,
    input [M_AXIS_BRAM_17_WIDTH/8-1:0] ap_bram_oarg_17_we1,
    input ap_bram_oarg_17_en1,
    //out BRAM to AXI-Stream interface 18
    input m_axis_bram_18_aclk,
    input m_axis_bram_18_aresetn,
    output m_axis_bram_18_tlast,
    output m_axis_bram_18_tvalid,
    output [M_AXIS_BRAM_18_DMWIDTH/8-1:0] m_axis_bram_18_tkeep,
    output [M_AXIS_BRAM_18_DMWIDTH/8-1:0] m_axis_bram_18_tstrb,
    output [M_AXIS_BRAM_18_DMWIDTH-1:0] m_axis_bram_18_tdata,
    input m_axis_bram_18_tready,
    input [M_AXIS_BRAM_18_ADDR_WIDTH-1:0] ap_bram_oarg_18_addr0,
    input [M_AXIS_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_din0,
    output [M_AXIS_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_dout0,
    input ap_bram_oarg_18_clk0,
    input ap_bram_oarg_18_rst0,
    input [M_AXIS_BRAM_18_WIDTH/8-1:0] ap_bram_oarg_18_we0,
    input ap_bram_oarg_18_en0,
    input [M_AXIS_BRAM_18_ADDR_WIDTH-1:0] ap_bram_oarg_18_addr1,
    input [M_AXIS_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_din1,
    output [M_AXIS_BRAM_18_WIDTH-1:0] ap_bram_oarg_18_dout1,
    input ap_bram_oarg_18_clk1,
    input ap_bram_oarg_18_rst1,
    input [M_AXIS_BRAM_18_WIDTH/8-1:0] ap_bram_oarg_18_we1,
    input ap_bram_oarg_18_en1,
    //out BRAM to AXI-Stream interface 19
    input m_axis_bram_19_aclk,
    input m_axis_bram_19_aresetn,
    output m_axis_bram_19_tlast,
    output m_axis_bram_19_tvalid,
    output [M_AXIS_BRAM_19_DMWIDTH/8-1:0] m_axis_bram_19_tkeep,
    output [M_AXIS_BRAM_19_DMWIDTH/8-1:0] m_axis_bram_19_tstrb,
    output [M_AXIS_BRAM_19_DMWIDTH-1:0] m_axis_bram_19_tdata,
    input m_axis_bram_19_tready,
    input [M_AXIS_BRAM_19_ADDR_WIDTH-1:0] ap_bram_oarg_19_addr0,
    input [M_AXIS_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_din0,
    output [M_AXIS_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_dout0,
    input ap_bram_oarg_19_clk0,
    input ap_bram_oarg_19_rst0,
    input [M_AXIS_BRAM_19_WIDTH/8-1:0] ap_bram_oarg_19_we0,
    input ap_bram_oarg_19_en0,
    input [M_AXIS_BRAM_19_ADDR_WIDTH-1:0] ap_bram_oarg_19_addr1,
    input [M_AXIS_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_din1,
    output [M_AXIS_BRAM_19_WIDTH-1:0] ap_bram_oarg_19_dout1,
    input ap_bram_oarg_19_clk1,
    input ap_bram_oarg_19_rst1,
    input [M_AXIS_BRAM_19_WIDTH/8-1:0] ap_bram_oarg_19_we1,
    input ap_bram_oarg_19_en1,
    //out BRAM to AXI-Stream interface 20
    input m_axis_bram_20_aclk,
    input m_axis_bram_20_aresetn,
    output m_axis_bram_20_tlast,
    output m_axis_bram_20_tvalid,
    output [M_AXIS_BRAM_20_DMWIDTH/8-1:0] m_axis_bram_20_tkeep,
    output [M_AXIS_BRAM_20_DMWIDTH/8-1:0] m_axis_bram_20_tstrb,
    output [M_AXIS_BRAM_20_DMWIDTH-1:0] m_axis_bram_20_tdata,
    input m_axis_bram_20_tready,
    input [M_AXIS_BRAM_20_ADDR_WIDTH-1:0] ap_bram_oarg_20_addr0,
    input [M_AXIS_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_din0,
    output [M_AXIS_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_dout0,
    input ap_bram_oarg_20_clk0,
    input ap_bram_oarg_20_rst0,
    input [M_AXIS_BRAM_20_WIDTH/8-1:0] ap_bram_oarg_20_we0,
    input ap_bram_oarg_20_en0,
    input [M_AXIS_BRAM_20_ADDR_WIDTH-1:0] ap_bram_oarg_20_addr1,
    input [M_AXIS_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_din1,
    output [M_AXIS_BRAM_20_WIDTH-1:0] ap_bram_oarg_20_dout1,
    input ap_bram_oarg_20_clk1,
    input ap_bram_oarg_20_rst1,
    input [M_AXIS_BRAM_20_WIDTH/8-1:0] ap_bram_oarg_20_we1,
    input ap_bram_oarg_20_en1,
    //out BRAM to AXI-Stream interface 21
    input m_axis_bram_21_aclk,
    input m_axis_bram_21_aresetn,
    output m_axis_bram_21_tlast,
    output m_axis_bram_21_tvalid,
    output [M_AXIS_BRAM_21_DMWIDTH/8-1:0] m_axis_bram_21_tkeep,
    output [M_AXIS_BRAM_21_DMWIDTH/8-1:0] m_axis_bram_21_tstrb,
    output [M_AXIS_BRAM_21_DMWIDTH-1:0] m_axis_bram_21_tdata,
    input m_axis_bram_21_tready,
    input [M_AXIS_BRAM_21_ADDR_WIDTH-1:0] ap_bram_oarg_21_addr0,
    input [M_AXIS_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_din0,
    output [M_AXIS_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_dout0,
    input ap_bram_oarg_21_clk0,
    input ap_bram_oarg_21_rst0,
    input [M_AXIS_BRAM_21_WIDTH/8-1:0] ap_bram_oarg_21_we0,
    input ap_bram_oarg_21_en0,
    input [M_AXIS_BRAM_21_ADDR_WIDTH-1:0] ap_bram_oarg_21_addr1,
    input [M_AXIS_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_din1,
    output [M_AXIS_BRAM_21_WIDTH-1:0] ap_bram_oarg_21_dout1,
    input ap_bram_oarg_21_clk1,
    input ap_bram_oarg_21_rst1,
    input [M_AXIS_BRAM_21_WIDTH/8-1:0] ap_bram_oarg_21_we1,
    input ap_bram_oarg_21_en1,
    //out BRAM to AXI-Stream interface 22
    input m_axis_bram_22_aclk,
    input m_axis_bram_22_aresetn,
    output m_axis_bram_22_tlast,
    output m_axis_bram_22_tvalid,
    output [M_AXIS_BRAM_22_DMWIDTH/8-1:0] m_axis_bram_22_tkeep,
    output [M_AXIS_BRAM_22_DMWIDTH/8-1:0] m_axis_bram_22_tstrb,
    output [M_AXIS_BRAM_22_DMWIDTH-1:0] m_axis_bram_22_tdata,
    input m_axis_bram_22_tready,
    input [M_AXIS_BRAM_22_ADDR_WIDTH-1:0] ap_bram_oarg_22_addr0,
    input [M_AXIS_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_din0,
    output [M_AXIS_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_dout0,
    input ap_bram_oarg_22_clk0,
    input ap_bram_oarg_22_rst0,
    input [M_AXIS_BRAM_22_WIDTH/8-1:0] ap_bram_oarg_22_we0,
    input ap_bram_oarg_22_en0,
    input [M_AXIS_BRAM_22_ADDR_WIDTH-1:0] ap_bram_oarg_22_addr1,
    input [M_AXIS_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_din1,
    output [M_AXIS_BRAM_22_WIDTH-1:0] ap_bram_oarg_22_dout1,
    input ap_bram_oarg_22_clk1,
    input ap_bram_oarg_22_rst1,
    input [M_AXIS_BRAM_22_WIDTH/8-1:0] ap_bram_oarg_22_we1,
    input ap_bram_oarg_22_en1,
    //out BRAM to AXI-Stream interface 23
    input m_axis_bram_23_aclk,
    input m_axis_bram_23_aresetn,
    output m_axis_bram_23_tlast,
    output m_axis_bram_23_tvalid,
    output [M_AXIS_BRAM_23_DMWIDTH/8-1:0] m_axis_bram_23_tkeep,
    output [M_AXIS_BRAM_23_DMWIDTH/8-1:0] m_axis_bram_23_tstrb,
    output [M_AXIS_BRAM_23_DMWIDTH-1:0] m_axis_bram_23_tdata,
    input m_axis_bram_23_tready,
    input [M_AXIS_BRAM_23_ADDR_WIDTH-1:0] ap_bram_oarg_23_addr0,
    input [M_AXIS_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_din0,
    output [M_AXIS_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_dout0,
    input ap_bram_oarg_23_clk0,
    input ap_bram_oarg_23_rst0,
    input [M_AXIS_BRAM_23_WIDTH/8-1:0] ap_bram_oarg_23_we0,
    input ap_bram_oarg_23_en0,
    input [M_AXIS_BRAM_23_ADDR_WIDTH-1:0] ap_bram_oarg_23_addr1,
    input [M_AXIS_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_din1,
    output [M_AXIS_BRAM_23_WIDTH-1:0] ap_bram_oarg_23_dout1,
    input ap_bram_oarg_23_clk1,
    input ap_bram_oarg_23_rst1,
    input [M_AXIS_BRAM_23_WIDTH/8-1:0] ap_bram_oarg_23_we1,
    input ap_bram_oarg_23_en1,
    //out BRAM to AXI-Stream interface 24
    input m_axis_bram_24_aclk,
    input m_axis_bram_24_aresetn,
    output m_axis_bram_24_tlast,
    output m_axis_bram_24_tvalid,
    output [M_AXIS_BRAM_24_DMWIDTH/8-1:0] m_axis_bram_24_tkeep,
    output [M_AXIS_BRAM_24_DMWIDTH/8-1:0] m_axis_bram_24_tstrb,
    output [M_AXIS_BRAM_24_DMWIDTH-1:0] m_axis_bram_24_tdata,
    input m_axis_bram_24_tready,
    input [M_AXIS_BRAM_24_ADDR_WIDTH-1:0] ap_bram_oarg_24_addr0,
    input [M_AXIS_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_din0,
    output [M_AXIS_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_dout0,
    input ap_bram_oarg_24_clk0,
    input ap_bram_oarg_24_rst0,
    input [M_AXIS_BRAM_24_WIDTH/8-1:0] ap_bram_oarg_24_we0,
    input ap_bram_oarg_24_en0,
    input [M_AXIS_BRAM_24_ADDR_WIDTH-1:0] ap_bram_oarg_24_addr1,
    input [M_AXIS_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_din1,
    output [M_AXIS_BRAM_24_WIDTH-1:0] ap_bram_oarg_24_dout1,
    input ap_bram_oarg_24_clk1,
    input ap_bram_oarg_24_rst1,
    input [M_AXIS_BRAM_24_WIDTH/8-1:0] ap_bram_oarg_24_we1,
    input ap_bram_oarg_24_en1,
    //out BRAM to AXI-Stream interface 25
    input m_axis_bram_25_aclk,
    input m_axis_bram_25_aresetn,
    output m_axis_bram_25_tlast,
    output m_axis_bram_25_tvalid,
    output [M_AXIS_BRAM_25_DMWIDTH/8-1:0] m_axis_bram_25_tkeep,
    output [M_AXIS_BRAM_25_DMWIDTH/8-1:0] m_axis_bram_25_tstrb,
    output [M_AXIS_BRAM_25_DMWIDTH-1:0] m_axis_bram_25_tdata,
    input m_axis_bram_25_tready,
    input [M_AXIS_BRAM_25_ADDR_WIDTH-1:0] ap_bram_oarg_25_addr0,
    input [M_AXIS_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_din0,
    output [M_AXIS_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_dout0,
    input ap_bram_oarg_25_clk0,
    input ap_bram_oarg_25_rst0,
    input [M_AXIS_BRAM_25_WIDTH/8-1:0] ap_bram_oarg_25_we0,
    input ap_bram_oarg_25_en0,
    input [M_AXIS_BRAM_25_ADDR_WIDTH-1:0] ap_bram_oarg_25_addr1,
    input [M_AXIS_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_din1,
    output [M_AXIS_BRAM_25_WIDTH-1:0] ap_bram_oarg_25_dout1,
    input ap_bram_oarg_25_clk1,
    input ap_bram_oarg_25_rst1,
    input [M_AXIS_BRAM_25_WIDTH/8-1:0] ap_bram_oarg_25_we1,
    input ap_bram_oarg_25_en1,
    //out BRAM to AXI-Stream interface 26
    input m_axis_bram_26_aclk,
    input m_axis_bram_26_aresetn,
    output m_axis_bram_26_tlast,
    output m_axis_bram_26_tvalid,
    output [M_AXIS_BRAM_26_DMWIDTH/8-1:0] m_axis_bram_26_tkeep,
    output [M_AXIS_BRAM_26_DMWIDTH/8-1:0] m_axis_bram_26_tstrb,
    output [M_AXIS_BRAM_26_DMWIDTH-1:0] m_axis_bram_26_tdata,
    input m_axis_bram_26_tready,
    input [M_AXIS_BRAM_26_ADDR_WIDTH-1:0] ap_bram_oarg_26_addr0,
    input [M_AXIS_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_din0,
    output [M_AXIS_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_dout0,
    input ap_bram_oarg_26_clk0,
    input ap_bram_oarg_26_rst0,
    input [M_AXIS_BRAM_26_WIDTH/8-1:0] ap_bram_oarg_26_we0,
    input ap_bram_oarg_26_en0,
    input [M_AXIS_BRAM_26_ADDR_WIDTH-1:0] ap_bram_oarg_26_addr1,
    input [M_AXIS_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_din1,
    output [M_AXIS_BRAM_26_WIDTH-1:0] ap_bram_oarg_26_dout1,
    input ap_bram_oarg_26_clk1,
    input ap_bram_oarg_26_rst1,
    input [M_AXIS_BRAM_26_WIDTH/8-1:0] ap_bram_oarg_26_we1,
    input ap_bram_oarg_26_en1,
    //out BRAM to AXI-Stream interface 27
    input m_axis_bram_27_aclk,
    input m_axis_bram_27_aresetn,
    output m_axis_bram_27_tlast,
    output m_axis_bram_27_tvalid,
    output [M_AXIS_BRAM_27_DMWIDTH/8-1:0] m_axis_bram_27_tkeep,
    output [M_AXIS_BRAM_27_DMWIDTH/8-1:0] m_axis_bram_27_tstrb,
    output [M_AXIS_BRAM_27_DMWIDTH-1:0] m_axis_bram_27_tdata,
    input m_axis_bram_27_tready,
    input [M_AXIS_BRAM_27_ADDR_WIDTH-1:0] ap_bram_oarg_27_addr0,
    input [M_AXIS_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_din0,
    output [M_AXIS_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_dout0,
    input ap_bram_oarg_27_clk0,
    input ap_bram_oarg_27_rst0,
    input [M_AXIS_BRAM_27_WIDTH/8-1:0] ap_bram_oarg_27_we0,
    input ap_bram_oarg_27_en0,
    input [M_AXIS_BRAM_27_ADDR_WIDTH-1:0] ap_bram_oarg_27_addr1,
    input [M_AXIS_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_din1,
    output [M_AXIS_BRAM_27_WIDTH-1:0] ap_bram_oarg_27_dout1,
    input ap_bram_oarg_27_clk1,
    input ap_bram_oarg_27_rst1,
    input [M_AXIS_BRAM_27_WIDTH/8-1:0] ap_bram_oarg_27_we1,
    input ap_bram_oarg_27_en1,
    //out BRAM to AXI-Stream interface 28
    input m_axis_bram_28_aclk,
    input m_axis_bram_28_aresetn,
    output m_axis_bram_28_tlast,
    output m_axis_bram_28_tvalid,
    output [M_AXIS_BRAM_28_DMWIDTH/8-1:0] m_axis_bram_28_tkeep,
    output [M_AXIS_BRAM_28_DMWIDTH/8-1:0] m_axis_bram_28_tstrb,
    output [M_AXIS_BRAM_28_DMWIDTH-1:0] m_axis_bram_28_tdata,
    input m_axis_bram_28_tready,
    input [M_AXIS_BRAM_28_ADDR_WIDTH-1:0] ap_bram_oarg_28_addr0,
    input [M_AXIS_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_din0,
    output [M_AXIS_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_dout0,
    input ap_bram_oarg_28_clk0,
    input ap_bram_oarg_28_rst0,
    input [M_AXIS_BRAM_28_WIDTH/8-1:0] ap_bram_oarg_28_we0,
    input ap_bram_oarg_28_en0,
    input [M_AXIS_BRAM_28_ADDR_WIDTH-1:0] ap_bram_oarg_28_addr1,
    input [M_AXIS_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_din1,
    output [M_AXIS_BRAM_28_WIDTH-1:0] ap_bram_oarg_28_dout1,
    input ap_bram_oarg_28_clk1,
    input ap_bram_oarg_28_rst1,
    input [M_AXIS_BRAM_28_WIDTH/8-1:0] ap_bram_oarg_28_we1,
    input ap_bram_oarg_28_en1,
    //out BRAM to AXI-Stream interface 29
    input m_axis_bram_29_aclk,
    input m_axis_bram_29_aresetn,
    output m_axis_bram_29_tlast,
    output m_axis_bram_29_tvalid,
    output [M_AXIS_BRAM_29_DMWIDTH/8-1:0] m_axis_bram_29_tkeep,
    output [M_AXIS_BRAM_29_DMWIDTH/8-1:0] m_axis_bram_29_tstrb,
    output [M_AXIS_BRAM_29_DMWIDTH-1:0] m_axis_bram_29_tdata,
    input m_axis_bram_29_tready,
    input [M_AXIS_BRAM_29_ADDR_WIDTH-1:0] ap_bram_oarg_29_addr0,
    input [M_AXIS_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_din0,
    output [M_AXIS_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_dout0,
    input ap_bram_oarg_29_clk0,
    input ap_bram_oarg_29_rst0,
    input [M_AXIS_BRAM_29_WIDTH/8-1:0] ap_bram_oarg_29_we0,
    input ap_bram_oarg_29_en0,
    input [M_AXIS_BRAM_29_ADDR_WIDTH-1:0] ap_bram_oarg_29_addr1,
    input [M_AXIS_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_din1,
    output [M_AXIS_BRAM_29_WIDTH-1:0] ap_bram_oarg_29_dout1,
    input ap_bram_oarg_29_clk1,
    input ap_bram_oarg_29_rst1,
    input [M_AXIS_BRAM_29_WIDTH/8-1:0] ap_bram_oarg_29_we1,
    input ap_bram_oarg_29_en1,
    //out BRAM to AXI-Stream interface 30
    input m_axis_bram_30_aclk,
    input m_axis_bram_30_aresetn,
    output m_axis_bram_30_tlast,
    output m_axis_bram_30_tvalid,
    output [M_AXIS_BRAM_30_DMWIDTH/8-1:0] m_axis_bram_30_tkeep,
    output [M_AXIS_BRAM_30_DMWIDTH/8-1:0] m_axis_bram_30_tstrb,
    output [M_AXIS_BRAM_30_DMWIDTH-1:0] m_axis_bram_30_tdata,
    input m_axis_bram_30_tready,
    input [M_AXIS_BRAM_30_ADDR_WIDTH-1:0] ap_bram_oarg_30_addr0,
    input [M_AXIS_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_din0,
    output [M_AXIS_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_dout0,
    input ap_bram_oarg_30_clk0,
    input ap_bram_oarg_30_rst0,
    input [M_AXIS_BRAM_30_WIDTH/8-1:0] ap_bram_oarg_30_we0,
    input ap_bram_oarg_30_en0,
    input [M_AXIS_BRAM_30_ADDR_WIDTH-1:0] ap_bram_oarg_30_addr1,
    input [M_AXIS_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_din1,
    output [M_AXIS_BRAM_30_WIDTH-1:0] ap_bram_oarg_30_dout1,
    input ap_bram_oarg_30_clk1,
    input ap_bram_oarg_30_rst1,
    input [M_AXIS_BRAM_30_WIDTH/8-1:0] ap_bram_oarg_30_we1,
    input ap_bram_oarg_30_en1,
    //out BRAM to AXI-Stream interface 31
    input m_axis_bram_31_aclk,
    input m_axis_bram_31_aresetn,
    output m_axis_bram_31_tlast,
    output m_axis_bram_31_tvalid,
    output [M_AXIS_BRAM_31_DMWIDTH/8-1:0] m_axis_bram_31_tkeep,
    output [M_AXIS_BRAM_31_DMWIDTH/8-1:0] m_axis_bram_31_tstrb,
    output [M_AXIS_BRAM_31_DMWIDTH-1:0] m_axis_bram_31_tdata,
    input m_axis_bram_31_tready,
    input [M_AXIS_BRAM_31_ADDR_WIDTH-1:0] ap_bram_oarg_31_addr0,
    input [M_AXIS_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_din0,
    output [M_AXIS_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_dout0,
    input ap_bram_oarg_31_clk0,
    input ap_bram_oarg_31_rst0,
    input [M_AXIS_BRAM_31_WIDTH/8-1:0] ap_bram_oarg_31_we0,
    input ap_bram_oarg_31_en0,
    input [M_AXIS_BRAM_31_ADDR_WIDTH-1:0] ap_bram_oarg_31_addr1,
    input [M_AXIS_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_din1,
    output [M_AXIS_BRAM_31_WIDTH-1:0] ap_bram_oarg_31_dout1,
    input ap_bram_oarg_31_clk1,
    input ap_bram_oarg_31_rst1,
    input [M_AXIS_BRAM_31_WIDTH/8-1:0] ap_bram_oarg_31_we1,
    input ap_bram_oarg_31_en1,
    //out BRAM to AXI-Stream interface 32
    input m_axis_bram_32_aclk,
    input m_axis_bram_32_aresetn,
    output m_axis_bram_32_tlast,
    output m_axis_bram_32_tvalid,
    output [M_AXIS_BRAM_32_DMWIDTH/8-1:0] m_axis_bram_32_tkeep,
    output [M_AXIS_BRAM_32_DMWIDTH/8-1:0] m_axis_bram_32_tstrb,
    output [M_AXIS_BRAM_32_DMWIDTH-1:0] m_axis_bram_32_tdata,
    input m_axis_bram_32_tready,
    input [M_AXIS_BRAM_32_ADDR_WIDTH-1:0] ap_bram_oarg_32_addr0,
    input [M_AXIS_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_din0,
    output [M_AXIS_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_dout0,
    input ap_bram_oarg_32_clk0,
    input ap_bram_oarg_32_rst0,
    input [M_AXIS_BRAM_32_WIDTH/8-1:0] ap_bram_oarg_32_we0,
    input ap_bram_oarg_32_en0,
    input [M_AXIS_BRAM_32_ADDR_WIDTH-1:0] ap_bram_oarg_32_addr1,
    input [M_AXIS_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_din1,
    output [M_AXIS_BRAM_32_WIDTH-1:0] ap_bram_oarg_32_dout1,
    input ap_bram_oarg_32_clk1,
    input ap_bram_oarg_32_rst1,
    input [M_AXIS_BRAM_32_WIDTH/8-1:0] ap_bram_oarg_32_we1,
    input ap_bram_oarg_32_en1,
    //out BRAM to AXI-Stream interface 33
    input m_axis_bram_33_aclk,
    input m_axis_bram_33_aresetn,
    output m_axis_bram_33_tlast,
    output m_axis_bram_33_tvalid,
    output [M_AXIS_BRAM_33_DMWIDTH/8-1:0] m_axis_bram_33_tkeep,
    output [M_AXIS_BRAM_33_DMWIDTH/8-1:0] m_axis_bram_33_tstrb,
    output [M_AXIS_BRAM_33_DMWIDTH-1:0] m_axis_bram_33_tdata,
    input m_axis_bram_33_tready,
    input [M_AXIS_BRAM_33_ADDR_WIDTH-1:0] ap_bram_oarg_33_addr0,
    input [M_AXIS_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_din0,
    output [M_AXIS_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_dout0,
    input ap_bram_oarg_33_clk0,
    input ap_bram_oarg_33_rst0,
    input [M_AXIS_BRAM_33_WIDTH/8-1:0] ap_bram_oarg_33_we0,
    input ap_bram_oarg_33_en0,
    input [M_AXIS_BRAM_33_ADDR_WIDTH-1:0] ap_bram_oarg_33_addr1,
    input [M_AXIS_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_din1,
    output [M_AXIS_BRAM_33_WIDTH-1:0] ap_bram_oarg_33_dout1,
    input ap_bram_oarg_33_clk1,
    input ap_bram_oarg_33_rst1,
    input [M_AXIS_BRAM_33_WIDTH/8-1:0] ap_bram_oarg_33_we1,
    input ap_bram_oarg_33_en1,
    //out BRAM to AXI-Stream interface 34
    input m_axis_bram_34_aclk,
    input m_axis_bram_34_aresetn,
    output m_axis_bram_34_tlast,
    output m_axis_bram_34_tvalid,
    output [M_AXIS_BRAM_34_DMWIDTH/8-1:0] m_axis_bram_34_tkeep,
    output [M_AXIS_BRAM_34_DMWIDTH/8-1:0] m_axis_bram_34_tstrb,
    output [M_AXIS_BRAM_34_DMWIDTH-1:0] m_axis_bram_34_tdata,
    input m_axis_bram_34_tready,
    input [M_AXIS_BRAM_34_ADDR_WIDTH-1:0] ap_bram_oarg_34_addr0,
    input [M_AXIS_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_din0,
    output [M_AXIS_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_dout0,
    input ap_bram_oarg_34_clk0,
    input ap_bram_oarg_34_rst0,
    input [M_AXIS_BRAM_34_WIDTH/8-1:0] ap_bram_oarg_34_we0,
    input ap_bram_oarg_34_en0,
    input [M_AXIS_BRAM_34_ADDR_WIDTH-1:0] ap_bram_oarg_34_addr1,
    input [M_AXIS_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_din1,
    output [M_AXIS_BRAM_34_WIDTH-1:0] ap_bram_oarg_34_dout1,
    input ap_bram_oarg_34_clk1,
    input ap_bram_oarg_34_rst1,
    input [M_AXIS_BRAM_34_WIDTH/8-1:0] ap_bram_oarg_34_we1,
    input ap_bram_oarg_34_en1,
    //out BRAM to AXI-Stream interface 35
    input m_axis_bram_35_aclk,
    input m_axis_bram_35_aresetn,
    output m_axis_bram_35_tlast,
    output m_axis_bram_35_tvalid,
    output [M_AXIS_BRAM_35_DMWIDTH/8-1:0] m_axis_bram_35_tkeep,
    output [M_AXIS_BRAM_35_DMWIDTH/8-1:0] m_axis_bram_35_tstrb,
    output [M_AXIS_BRAM_35_DMWIDTH-1:0] m_axis_bram_35_tdata,
    input m_axis_bram_35_tready,
    input [M_AXIS_BRAM_35_ADDR_WIDTH-1:0] ap_bram_oarg_35_addr0,
    input [M_AXIS_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_din0,
    output [M_AXIS_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_dout0,
    input ap_bram_oarg_35_clk0,
    input ap_bram_oarg_35_rst0,
    input [M_AXIS_BRAM_35_WIDTH/8-1:0] ap_bram_oarg_35_we0,
    input ap_bram_oarg_35_en0,
    input [M_AXIS_BRAM_35_ADDR_WIDTH-1:0] ap_bram_oarg_35_addr1,
    input [M_AXIS_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_din1,
    output [M_AXIS_BRAM_35_WIDTH-1:0] ap_bram_oarg_35_dout1,
    input ap_bram_oarg_35_clk1,
    input ap_bram_oarg_35_rst1,
    input [M_AXIS_BRAM_35_WIDTH/8-1:0] ap_bram_oarg_35_we1,
    input ap_bram_oarg_35_en1,
    //out BRAM to AXI-Stream interface 36
    input m_axis_bram_36_aclk,
    input m_axis_bram_36_aresetn,
    output m_axis_bram_36_tlast,
    output m_axis_bram_36_tvalid,
    output [M_AXIS_BRAM_36_DMWIDTH/8-1:0] m_axis_bram_36_tkeep,
    output [M_AXIS_BRAM_36_DMWIDTH/8-1:0] m_axis_bram_36_tstrb,
    output [M_AXIS_BRAM_36_DMWIDTH-1:0] m_axis_bram_36_tdata,
    input m_axis_bram_36_tready,
    input [M_AXIS_BRAM_36_ADDR_WIDTH-1:0] ap_bram_oarg_36_addr0,
    input [M_AXIS_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_din0,
    output [M_AXIS_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_dout0,
    input ap_bram_oarg_36_clk0,
    input ap_bram_oarg_36_rst0,
    input [M_AXIS_BRAM_36_WIDTH/8-1:0] ap_bram_oarg_36_we0,
    input ap_bram_oarg_36_en0,
    input [M_AXIS_BRAM_36_ADDR_WIDTH-1:0] ap_bram_oarg_36_addr1,
    input [M_AXIS_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_din1,
    output [M_AXIS_BRAM_36_WIDTH-1:0] ap_bram_oarg_36_dout1,
    input ap_bram_oarg_36_clk1,
    input ap_bram_oarg_36_rst1,
    input [M_AXIS_BRAM_36_WIDTH/8-1:0] ap_bram_oarg_36_we1,
    input ap_bram_oarg_36_en1,
    //out BRAM to AXI-Stream interface 37
    input m_axis_bram_37_aclk,
    input m_axis_bram_37_aresetn,
    output m_axis_bram_37_tlast,
    output m_axis_bram_37_tvalid,
    output [M_AXIS_BRAM_37_DMWIDTH/8-1:0] m_axis_bram_37_tkeep,
    output [M_AXIS_BRAM_37_DMWIDTH/8-1:0] m_axis_bram_37_tstrb,
    output [M_AXIS_BRAM_37_DMWIDTH-1:0] m_axis_bram_37_tdata,
    input m_axis_bram_37_tready,
    input [M_AXIS_BRAM_37_ADDR_WIDTH-1:0] ap_bram_oarg_37_addr0,
    input [M_AXIS_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_din0,
    output [M_AXIS_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_dout0,
    input ap_bram_oarg_37_clk0,
    input ap_bram_oarg_37_rst0,
    input [M_AXIS_BRAM_37_WIDTH/8-1:0] ap_bram_oarg_37_we0,
    input ap_bram_oarg_37_en0,
    input [M_AXIS_BRAM_37_ADDR_WIDTH-1:0] ap_bram_oarg_37_addr1,
    input [M_AXIS_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_din1,
    output [M_AXIS_BRAM_37_WIDTH-1:0] ap_bram_oarg_37_dout1,
    input ap_bram_oarg_37_clk1,
    input ap_bram_oarg_37_rst1,
    input [M_AXIS_BRAM_37_WIDTH/8-1:0] ap_bram_oarg_37_we1,
    input ap_bram_oarg_37_en1,
    //out BRAM to AXI-Stream interface 38
    input m_axis_bram_38_aclk,
    input m_axis_bram_38_aresetn,
    output m_axis_bram_38_tlast,
    output m_axis_bram_38_tvalid,
    output [M_AXIS_BRAM_38_DMWIDTH/8-1:0] m_axis_bram_38_tkeep,
    output [M_AXIS_BRAM_38_DMWIDTH/8-1:0] m_axis_bram_38_tstrb,
    output [M_AXIS_BRAM_38_DMWIDTH-1:0] m_axis_bram_38_tdata,
    input m_axis_bram_38_tready,
    input [M_AXIS_BRAM_38_ADDR_WIDTH-1:0] ap_bram_oarg_38_addr0,
    input [M_AXIS_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_din0,
    output [M_AXIS_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_dout0,
    input ap_bram_oarg_38_clk0,
    input ap_bram_oarg_38_rst0,
    input [M_AXIS_BRAM_38_WIDTH/8-1:0] ap_bram_oarg_38_we0,
    input ap_bram_oarg_38_en0,
    input [M_AXIS_BRAM_38_ADDR_WIDTH-1:0] ap_bram_oarg_38_addr1,
    input [M_AXIS_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_din1,
    output [M_AXIS_BRAM_38_WIDTH-1:0] ap_bram_oarg_38_dout1,
    input ap_bram_oarg_38_clk1,
    input ap_bram_oarg_38_rst1,
    input [M_AXIS_BRAM_38_WIDTH/8-1:0] ap_bram_oarg_38_we1,
    input ap_bram_oarg_38_en1,
    //out BRAM to AXI-Stream interface 39
    input m_axis_bram_39_aclk,
    input m_axis_bram_39_aresetn,
    output m_axis_bram_39_tlast,
    output m_axis_bram_39_tvalid,
    output [M_AXIS_BRAM_39_DMWIDTH/8-1:0] m_axis_bram_39_tkeep,
    output [M_AXIS_BRAM_39_DMWIDTH/8-1:0] m_axis_bram_39_tstrb,
    output [M_AXIS_BRAM_39_DMWIDTH-1:0] m_axis_bram_39_tdata,
    input m_axis_bram_39_tready,
    input [M_AXIS_BRAM_39_ADDR_WIDTH-1:0] ap_bram_oarg_39_addr0,
    input [M_AXIS_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_din0,
    output [M_AXIS_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_dout0,
    input ap_bram_oarg_39_clk0,
    input ap_bram_oarg_39_rst0,
    input [M_AXIS_BRAM_39_WIDTH/8-1:0] ap_bram_oarg_39_we0,
    input ap_bram_oarg_39_en0,
    input [M_AXIS_BRAM_39_ADDR_WIDTH-1:0] ap_bram_oarg_39_addr1,
    input [M_AXIS_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_din1,
    output [M_AXIS_BRAM_39_WIDTH-1:0] ap_bram_oarg_39_dout1,
    input ap_bram_oarg_39_clk1,
    input ap_bram_oarg_39_rst1,
    input [M_AXIS_BRAM_39_WIDTH/8-1:0] ap_bram_oarg_39_we1,
    input ap_bram_oarg_39_en1,
    //out BRAM to AXI-Stream interface 40
    input m_axis_bram_40_aclk,
    input m_axis_bram_40_aresetn,
    output m_axis_bram_40_tlast,
    output m_axis_bram_40_tvalid,
    output [M_AXIS_BRAM_40_DMWIDTH/8-1:0] m_axis_bram_40_tkeep,
    output [M_AXIS_BRAM_40_DMWIDTH/8-1:0] m_axis_bram_40_tstrb,
    output [M_AXIS_BRAM_40_DMWIDTH-1:0] m_axis_bram_40_tdata,
    input m_axis_bram_40_tready,
    input [M_AXIS_BRAM_40_ADDR_WIDTH-1:0] ap_bram_oarg_40_addr0,
    input [M_AXIS_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_din0,
    output [M_AXIS_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_dout0,
    input ap_bram_oarg_40_clk0,
    input ap_bram_oarg_40_rst0,
    input [M_AXIS_BRAM_40_WIDTH/8-1:0] ap_bram_oarg_40_we0,
    input ap_bram_oarg_40_en0,
    input [M_AXIS_BRAM_40_ADDR_WIDTH-1:0] ap_bram_oarg_40_addr1,
    input [M_AXIS_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_din1,
    output [M_AXIS_BRAM_40_WIDTH-1:0] ap_bram_oarg_40_dout1,
    input ap_bram_oarg_40_clk1,
    input ap_bram_oarg_40_rst1,
    input [M_AXIS_BRAM_40_WIDTH/8-1:0] ap_bram_oarg_40_we1,
    input ap_bram_oarg_40_en1,
    //out BRAM to AXI-Stream interface 41
    input m_axis_bram_41_aclk,
    input m_axis_bram_41_aresetn,
    output m_axis_bram_41_tlast,
    output m_axis_bram_41_tvalid,
    output [M_AXIS_BRAM_41_DMWIDTH/8-1:0] m_axis_bram_41_tkeep,
    output [M_AXIS_BRAM_41_DMWIDTH/8-1:0] m_axis_bram_41_tstrb,
    output [M_AXIS_BRAM_41_DMWIDTH-1:0] m_axis_bram_41_tdata,
    input m_axis_bram_41_tready,
    input [M_AXIS_BRAM_41_ADDR_WIDTH-1:0] ap_bram_oarg_41_addr0,
    input [M_AXIS_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_din0,
    output [M_AXIS_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_dout0,
    input ap_bram_oarg_41_clk0,
    input ap_bram_oarg_41_rst0,
    input [M_AXIS_BRAM_41_WIDTH/8-1:0] ap_bram_oarg_41_we0,
    input ap_bram_oarg_41_en0,
    input [M_AXIS_BRAM_41_ADDR_WIDTH-1:0] ap_bram_oarg_41_addr1,
    input [M_AXIS_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_din1,
    output [M_AXIS_BRAM_41_WIDTH-1:0] ap_bram_oarg_41_dout1,
    input ap_bram_oarg_41_clk1,
    input ap_bram_oarg_41_rst1,
    input [M_AXIS_BRAM_41_WIDTH/8-1:0] ap_bram_oarg_41_we1,
    input ap_bram_oarg_41_en1,
    //out BRAM to AXI-Stream interface 42
    input m_axis_bram_42_aclk,
    input m_axis_bram_42_aresetn,
    output m_axis_bram_42_tlast,
    output m_axis_bram_42_tvalid,
    output [M_AXIS_BRAM_42_DMWIDTH/8-1:0] m_axis_bram_42_tkeep,
    output [M_AXIS_BRAM_42_DMWIDTH/8-1:0] m_axis_bram_42_tstrb,
    output [M_AXIS_BRAM_42_DMWIDTH-1:0] m_axis_bram_42_tdata,
    input m_axis_bram_42_tready,
    input [M_AXIS_BRAM_42_ADDR_WIDTH-1:0] ap_bram_oarg_42_addr0,
    input [M_AXIS_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_din0,
    output [M_AXIS_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_dout0,
    input ap_bram_oarg_42_clk0,
    input ap_bram_oarg_42_rst0,
    input [M_AXIS_BRAM_42_WIDTH/8-1:0] ap_bram_oarg_42_we0,
    input ap_bram_oarg_42_en0,
    input [M_AXIS_BRAM_42_ADDR_WIDTH-1:0] ap_bram_oarg_42_addr1,
    input [M_AXIS_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_din1,
    output [M_AXIS_BRAM_42_WIDTH-1:0] ap_bram_oarg_42_dout1,
    input ap_bram_oarg_42_clk1,
    input ap_bram_oarg_42_rst1,
    input [M_AXIS_BRAM_42_WIDTH/8-1:0] ap_bram_oarg_42_we1,
    input ap_bram_oarg_42_en1,
    //out BRAM to AXI-Stream interface 43
    input m_axis_bram_43_aclk,
    input m_axis_bram_43_aresetn,
    output m_axis_bram_43_tlast,
    output m_axis_bram_43_tvalid,
    output [M_AXIS_BRAM_43_DMWIDTH/8-1:0] m_axis_bram_43_tkeep,
    output [M_AXIS_BRAM_43_DMWIDTH/8-1:0] m_axis_bram_43_tstrb,
    output [M_AXIS_BRAM_43_DMWIDTH-1:0] m_axis_bram_43_tdata,
    input m_axis_bram_43_tready,
    input [M_AXIS_BRAM_43_ADDR_WIDTH-1:0] ap_bram_oarg_43_addr0,
    input [M_AXIS_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_din0,
    output [M_AXIS_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_dout0,
    input ap_bram_oarg_43_clk0,
    input ap_bram_oarg_43_rst0,
    input [M_AXIS_BRAM_43_WIDTH/8-1:0] ap_bram_oarg_43_we0,
    input ap_bram_oarg_43_en0,
    input [M_AXIS_BRAM_43_ADDR_WIDTH-1:0] ap_bram_oarg_43_addr1,
    input [M_AXIS_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_din1,
    output [M_AXIS_BRAM_43_WIDTH-1:0] ap_bram_oarg_43_dout1,
    input ap_bram_oarg_43_clk1,
    input ap_bram_oarg_43_rst1,
    input [M_AXIS_BRAM_43_WIDTH/8-1:0] ap_bram_oarg_43_we1,
    input ap_bram_oarg_43_en1,
    //out BRAM to AXI-Stream interface 44
    input m_axis_bram_44_aclk,
    input m_axis_bram_44_aresetn,
    output m_axis_bram_44_tlast,
    output m_axis_bram_44_tvalid,
    output [M_AXIS_BRAM_44_DMWIDTH/8-1:0] m_axis_bram_44_tkeep,
    output [M_AXIS_BRAM_44_DMWIDTH/8-1:0] m_axis_bram_44_tstrb,
    output [M_AXIS_BRAM_44_DMWIDTH-1:0] m_axis_bram_44_tdata,
    input m_axis_bram_44_tready,
    input [M_AXIS_BRAM_44_ADDR_WIDTH-1:0] ap_bram_oarg_44_addr0,
    input [M_AXIS_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_din0,
    output [M_AXIS_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_dout0,
    input ap_bram_oarg_44_clk0,
    input ap_bram_oarg_44_rst0,
    input [M_AXIS_BRAM_44_WIDTH/8-1:0] ap_bram_oarg_44_we0,
    input ap_bram_oarg_44_en0,
    input [M_AXIS_BRAM_44_ADDR_WIDTH-1:0] ap_bram_oarg_44_addr1,
    input [M_AXIS_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_din1,
    output [M_AXIS_BRAM_44_WIDTH-1:0] ap_bram_oarg_44_dout1,
    input ap_bram_oarg_44_clk1,
    input ap_bram_oarg_44_rst1,
    input [M_AXIS_BRAM_44_WIDTH/8-1:0] ap_bram_oarg_44_we1,
    input ap_bram_oarg_44_en1,
    //out BRAM to AXI-Stream interface 45
    input m_axis_bram_45_aclk,
    input m_axis_bram_45_aresetn,
    output m_axis_bram_45_tlast,
    output m_axis_bram_45_tvalid,
    output [M_AXIS_BRAM_45_DMWIDTH/8-1:0] m_axis_bram_45_tkeep,
    output [M_AXIS_BRAM_45_DMWIDTH/8-1:0] m_axis_bram_45_tstrb,
    output [M_AXIS_BRAM_45_DMWIDTH-1:0] m_axis_bram_45_tdata,
    input m_axis_bram_45_tready,
    input [M_AXIS_BRAM_45_ADDR_WIDTH-1:0] ap_bram_oarg_45_addr0,
    input [M_AXIS_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_din0,
    output [M_AXIS_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_dout0,
    input ap_bram_oarg_45_clk0,
    input ap_bram_oarg_45_rst0,
    input [M_AXIS_BRAM_45_WIDTH/8-1:0] ap_bram_oarg_45_we0,
    input ap_bram_oarg_45_en0,
    input [M_AXIS_BRAM_45_ADDR_WIDTH-1:0] ap_bram_oarg_45_addr1,
    input [M_AXIS_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_din1,
    output [M_AXIS_BRAM_45_WIDTH-1:0] ap_bram_oarg_45_dout1,
    input ap_bram_oarg_45_clk1,
    input ap_bram_oarg_45_rst1,
    input [M_AXIS_BRAM_45_WIDTH/8-1:0] ap_bram_oarg_45_we1,
    input ap_bram_oarg_45_en1,
    //out BRAM to AXI-Stream interface 46
    input m_axis_bram_46_aclk,
    input m_axis_bram_46_aresetn,
    output m_axis_bram_46_tlast,
    output m_axis_bram_46_tvalid,
    output [M_AXIS_BRAM_46_DMWIDTH/8-1:0] m_axis_bram_46_tkeep,
    output [M_AXIS_BRAM_46_DMWIDTH/8-1:0] m_axis_bram_46_tstrb,
    output [M_AXIS_BRAM_46_DMWIDTH-1:0] m_axis_bram_46_tdata,
    input m_axis_bram_46_tready,
    input [M_AXIS_BRAM_46_ADDR_WIDTH-1:0] ap_bram_oarg_46_addr0,
    input [M_AXIS_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_din0,
    output [M_AXIS_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_dout0,
    input ap_bram_oarg_46_clk0,
    input ap_bram_oarg_46_rst0,
    input [M_AXIS_BRAM_46_WIDTH/8-1:0] ap_bram_oarg_46_we0,
    input ap_bram_oarg_46_en0,
    input [M_AXIS_BRAM_46_ADDR_WIDTH-1:0] ap_bram_oarg_46_addr1,
    input [M_AXIS_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_din1,
    output [M_AXIS_BRAM_46_WIDTH-1:0] ap_bram_oarg_46_dout1,
    input ap_bram_oarg_46_clk1,
    input ap_bram_oarg_46_rst1,
    input [M_AXIS_BRAM_46_WIDTH/8-1:0] ap_bram_oarg_46_we1,
    input ap_bram_oarg_46_en1,
    //out BRAM to AXI-Stream interface 47
    input m_axis_bram_47_aclk,
    input m_axis_bram_47_aresetn,
    output m_axis_bram_47_tlast,
    output m_axis_bram_47_tvalid,
    output [M_AXIS_BRAM_47_DMWIDTH/8-1:0] m_axis_bram_47_tkeep,
    output [M_AXIS_BRAM_47_DMWIDTH/8-1:0] m_axis_bram_47_tstrb,
    output [M_AXIS_BRAM_47_DMWIDTH-1:0] m_axis_bram_47_tdata,
    input m_axis_bram_47_tready,
    input [M_AXIS_BRAM_47_ADDR_WIDTH-1:0] ap_bram_oarg_47_addr0,
    input [M_AXIS_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_din0,
    output [M_AXIS_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_dout0,
    input ap_bram_oarg_47_clk0,
    input ap_bram_oarg_47_rst0,
    input [M_AXIS_BRAM_47_WIDTH/8-1:0] ap_bram_oarg_47_we0,
    input ap_bram_oarg_47_en0,
    input [M_AXIS_BRAM_47_ADDR_WIDTH-1:0] ap_bram_oarg_47_addr1,
    input [M_AXIS_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_din1,
    output [M_AXIS_BRAM_47_WIDTH-1:0] ap_bram_oarg_47_dout1,
    input ap_bram_oarg_47_clk1,
    input ap_bram_oarg_47_rst1,
    input [M_AXIS_BRAM_47_WIDTH/8-1:0] ap_bram_oarg_47_we1,
    input ap_bram_oarg_47_en1,
    //out BRAM to AXI-Stream interface 48
    input m_axis_bram_48_aclk,
    input m_axis_bram_48_aresetn,
    output m_axis_bram_48_tlast,
    output m_axis_bram_48_tvalid,
    output [M_AXIS_BRAM_48_DMWIDTH/8-1:0] m_axis_bram_48_tkeep,
    output [M_AXIS_BRAM_48_DMWIDTH/8-1:0] m_axis_bram_48_tstrb,
    output [M_AXIS_BRAM_48_DMWIDTH-1:0] m_axis_bram_48_tdata,
    input m_axis_bram_48_tready,
    input [M_AXIS_BRAM_48_ADDR_WIDTH-1:0] ap_bram_oarg_48_addr0,
    input [M_AXIS_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_din0,
    output [M_AXIS_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_dout0,
    input ap_bram_oarg_48_clk0,
    input ap_bram_oarg_48_rst0,
    input [M_AXIS_BRAM_48_WIDTH/8-1:0] ap_bram_oarg_48_we0,
    input ap_bram_oarg_48_en0,
    input [M_AXIS_BRAM_48_ADDR_WIDTH-1:0] ap_bram_oarg_48_addr1,
    input [M_AXIS_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_din1,
    output [M_AXIS_BRAM_48_WIDTH-1:0] ap_bram_oarg_48_dout1,
    input ap_bram_oarg_48_clk1,
    input ap_bram_oarg_48_rst1,
    input [M_AXIS_BRAM_48_WIDTH/8-1:0] ap_bram_oarg_48_we1,
    input ap_bram_oarg_48_en1,
    //out BRAM to AXI-Stream interface 49
    input m_axis_bram_49_aclk,
    input m_axis_bram_49_aresetn,
    output m_axis_bram_49_tlast,
    output m_axis_bram_49_tvalid,
    output [M_AXIS_BRAM_49_DMWIDTH/8-1:0] m_axis_bram_49_tkeep,
    output [M_AXIS_BRAM_49_DMWIDTH/8-1:0] m_axis_bram_49_tstrb,
    output [M_AXIS_BRAM_49_DMWIDTH-1:0] m_axis_bram_49_tdata,
    input m_axis_bram_49_tready,
    input [M_AXIS_BRAM_49_ADDR_WIDTH-1:0] ap_bram_oarg_49_addr0,
    input [M_AXIS_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_din0,
    output [M_AXIS_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_dout0,
    input ap_bram_oarg_49_clk0,
    input ap_bram_oarg_49_rst0,
    input [M_AXIS_BRAM_49_WIDTH/8-1:0] ap_bram_oarg_49_we0,
    input ap_bram_oarg_49_en0,
    input [M_AXIS_BRAM_49_ADDR_WIDTH-1:0] ap_bram_oarg_49_addr1,
    input [M_AXIS_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_din1,
    output [M_AXIS_BRAM_49_WIDTH-1:0] ap_bram_oarg_49_dout1,
    input ap_bram_oarg_49_clk1,
    input ap_bram_oarg_49_rst1,
    input [M_AXIS_BRAM_49_WIDTH/8-1:0] ap_bram_oarg_49_we1,
    input ap_bram_oarg_49_en1,
    //out BRAM to AXI-Stream interface 50
    input m_axis_bram_50_aclk,
    input m_axis_bram_50_aresetn,
    output m_axis_bram_50_tlast,
    output m_axis_bram_50_tvalid,
    output [M_AXIS_BRAM_50_DMWIDTH/8-1:0] m_axis_bram_50_tkeep,
    output [M_AXIS_BRAM_50_DMWIDTH/8-1:0] m_axis_bram_50_tstrb,
    output [M_AXIS_BRAM_50_DMWIDTH-1:0] m_axis_bram_50_tdata,
    input m_axis_bram_50_tready,
    input [M_AXIS_BRAM_50_ADDR_WIDTH-1:0] ap_bram_oarg_50_addr0,
    input [M_AXIS_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_din0,
    output [M_AXIS_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_dout0,
    input ap_bram_oarg_50_clk0,
    input ap_bram_oarg_50_rst0,
    input [M_AXIS_BRAM_50_WIDTH/8-1:0] ap_bram_oarg_50_we0,
    input ap_bram_oarg_50_en0,
    input [M_AXIS_BRAM_50_ADDR_WIDTH-1:0] ap_bram_oarg_50_addr1,
    input [M_AXIS_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_din1,
    output [M_AXIS_BRAM_50_WIDTH-1:0] ap_bram_oarg_50_dout1,
    input ap_bram_oarg_50_clk1,
    input ap_bram_oarg_50_rst1,
    input [M_AXIS_BRAM_50_WIDTH/8-1:0] ap_bram_oarg_50_we1,
    input ap_bram_oarg_50_en1,
    //out BRAM to AXI-Stream interface 51
    input m_axis_bram_51_aclk,
    input m_axis_bram_51_aresetn,
    output m_axis_bram_51_tlast,
    output m_axis_bram_51_tvalid,
    output [M_AXIS_BRAM_51_DMWIDTH/8-1:0] m_axis_bram_51_tkeep,
    output [M_AXIS_BRAM_51_DMWIDTH/8-1:0] m_axis_bram_51_tstrb,
    output [M_AXIS_BRAM_51_DMWIDTH-1:0] m_axis_bram_51_tdata,
    input m_axis_bram_51_tready,
    input [M_AXIS_BRAM_51_ADDR_WIDTH-1:0] ap_bram_oarg_51_addr0,
    input [M_AXIS_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_din0,
    output [M_AXIS_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_dout0,
    input ap_bram_oarg_51_clk0,
    input ap_bram_oarg_51_rst0,
    input [M_AXIS_BRAM_51_WIDTH/8-1:0] ap_bram_oarg_51_we0,
    input ap_bram_oarg_51_en0,
    input [M_AXIS_BRAM_51_ADDR_WIDTH-1:0] ap_bram_oarg_51_addr1,
    input [M_AXIS_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_din1,
    output [M_AXIS_BRAM_51_WIDTH-1:0] ap_bram_oarg_51_dout1,
    input ap_bram_oarg_51_clk1,
    input ap_bram_oarg_51_rst1,
    input [M_AXIS_BRAM_51_WIDTH/8-1:0] ap_bram_oarg_51_we1,
    input ap_bram_oarg_51_en1,
    //out BRAM to AXI-Stream interface 52
    input m_axis_bram_52_aclk,
    input m_axis_bram_52_aresetn,
    output m_axis_bram_52_tlast,
    output m_axis_bram_52_tvalid,
    output [M_AXIS_BRAM_52_DMWIDTH/8-1:0] m_axis_bram_52_tkeep,
    output [M_AXIS_BRAM_52_DMWIDTH/8-1:0] m_axis_bram_52_tstrb,
    output [M_AXIS_BRAM_52_DMWIDTH-1:0] m_axis_bram_52_tdata,
    input m_axis_bram_52_tready,
    input [M_AXIS_BRAM_52_ADDR_WIDTH-1:0] ap_bram_oarg_52_addr0,
    input [M_AXIS_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_din0,
    output [M_AXIS_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_dout0,
    input ap_bram_oarg_52_clk0,
    input ap_bram_oarg_52_rst0,
    input [M_AXIS_BRAM_52_WIDTH/8-1:0] ap_bram_oarg_52_we0,
    input ap_bram_oarg_52_en0,
    input [M_AXIS_BRAM_52_ADDR_WIDTH-1:0] ap_bram_oarg_52_addr1,
    input [M_AXIS_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_din1,
    output [M_AXIS_BRAM_52_WIDTH-1:0] ap_bram_oarg_52_dout1,
    input ap_bram_oarg_52_clk1,
    input ap_bram_oarg_52_rst1,
    input [M_AXIS_BRAM_52_WIDTH/8-1:0] ap_bram_oarg_52_we1,
    input ap_bram_oarg_52_en1,
    //out BRAM to AXI-Stream interface 53
    input m_axis_bram_53_aclk,
    input m_axis_bram_53_aresetn,
    output m_axis_bram_53_tlast,
    output m_axis_bram_53_tvalid,
    output [M_AXIS_BRAM_53_DMWIDTH/8-1:0] m_axis_bram_53_tkeep,
    output [M_AXIS_BRAM_53_DMWIDTH/8-1:0] m_axis_bram_53_tstrb,
    output [M_AXIS_BRAM_53_DMWIDTH-1:0] m_axis_bram_53_tdata,
    input m_axis_bram_53_tready,
    input [M_AXIS_BRAM_53_ADDR_WIDTH-1:0] ap_bram_oarg_53_addr0,
    input [M_AXIS_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_din0,
    output [M_AXIS_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_dout0,
    input ap_bram_oarg_53_clk0,
    input ap_bram_oarg_53_rst0,
    input [M_AXIS_BRAM_53_WIDTH/8-1:0] ap_bram_oarg_53_we0,
    input ap_bram_oarg_53_en0,
    input [M_AXIS_BRAM_53_ADDR_WIDTH-1:0] ap_bram_oarg_53_addr1,
    input [M_AXIS_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_din1,
    output [M_AXIS_BRAM_53_WIDTH-1:0] ap_bram_oarg_53_dout1,
    input ap_bram_oarg_53_clk1,
    input ap_bram_oarg_53_rst1,
    input [M_AXIS_BRAM_53_WIDTH/8-1:0] ap_bram_oarg_53_we1,
    input ap_bram_oarg_53_en1,
    //out BRAM to AXI-Stream interface 54
    input m_axis_bram_54_aclk,
    input m_axis_bram_54_aresetn,
    output m_axis_bram_54_tlast,
    output m_axis_bram_54_tvalid,
    output [M_AXIS_BRAM_54_DMWIDTH/8-1:0] m_axis_bram_54_tkeep,
    output [M_AXIS_BRAM_54_DMWIDTH/8-1:0] m_axis_bram_54_tstrb,
    output [M_AXIS_BRAM_54_DMWIDTH-1:0] m_axis_bram_54_tdata,
    input m_axis_bram_54_tready,
    input [M_AXIS_BRAM_54_ADDR_WIDTH-1:0] ap_bram_oarg_54_addr0,
    input [M_AXIS_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_din0,
    output [M_AXIS_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_dout0,
    input ap_bram_oarg_54_clk0,
    input ap_bram_oarg_54_rst0,
    input [M_AXIS_BRAM_54_WIDTH/8-1:0] ap_bram_oarg_54_we0,
    input ap_bram_oarg_54_en0,
    input [M_AXIS_BRAM_54_ADDR_WIDTH-1:0] ap_bram_oarg_54_addr1,
    input [M_AXIS_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_din1,
    output [M_AXIS_BRAM_54_WIDTH-1:0] ap_bram_oarg_54_dout1,
    input ap_bram_oarg_54_clk1,
    input ap_bram_oarg_54_rst1,
    input [M_AXIS_BRAM_54_WIDTH/8-1:0] ap_bram_oarg_54_we1,
    input ap_bram_oarg_54_en1,
    //out BRAM to AXI-Stream interface 55
    input m_axis_bram_55_aclk,
    input m_axis_bram_55_aresetn,
    output m_axis_bram_55_tlast,
    output m_axis_bram_55_tvalid,
    output [M_AXIS_BRAM_55_DMWIDTH/8-1:0] m_axis_bram_55_tkeep,
    output [M_AXIS_BRAM_55_DMWIDTH/8-1:0] m_axis_bram_55_tstrb,
    output [M_AXIS_BRAM_55_DMWIDTH-1:0] m_axis_bram_55_tdata,
    input m_axis_bram_55_tready,
    input [M_AXIS_BRAM_55_ADDR_WIDTH-1:0] ap_bram_oarg_55_addr0,
    input [M_AXIS_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_din0,
    output [M_AXIS_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_dout0,
    input ap_bram_oarg_55_clk0,
    input ap_bram_oarg_55_rst0,
    input [M_AXIS_BRAM_55_WIDTH/8-1:0] ap_bram_oarg_55_we0,
    input ap_bram_oarg_55_en0,
    input [M_AXIS_BRAM_55_ADDR_WIDTH-1:0] ap_bram_oarg_55_addr1,
    input [M_AXIS_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_din1,
    output [M_AXIS_BRAM_55_WIDTH-1:0] ap_bram_oarg_55_dout1,
    input ap_bram_oarg_55_clk1,
    input ap_bram_oarg_55_rst1,
    input [M_AXIS_BRAM_55_WIDTH/8-1:0] ap_bram_oarg_55_we1,
    input ap_bram_oarg_55_en1,
    //out BRAM to AXI-Stream interface 56
    input m_axis_bram_56_aclk,
    input m_axis_bram_56_aresetn,
    output m_axis_bram_56_tlast,
    output m_axis_bram_56_tvalid,
    output [M_AXIS_BRAM_56_DMWIDTH/8-1:0] m_axis_bram_56_tkeep,
    output [M_AXIS_BRAM_56_DMWIDTH/8-1:0] m_axis_bram_56_tstrb,
    output [M_AXIS_BRAM_56_DMWIDTH-1:0] m_axis_bram_56_tdata,
    input m_axis_bram_56_tready,
    input [M_AXIS_BRAM_56_ADDR_WIDTH-1:0] ap_bram_oarg_56_addr0,
    input [M_AXIS_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_din0,
    output [M_AXIS_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_dout0,
    input ap_bram_oarg_56_clk0,
    input ap_bram_oarg_56_rst0,
    input [M_AXIS_BRAM_56_WIDTH/8-1:0] ap_bram_oarg_56_we0,
    input ap_bram_oarg_56_en0,
    input [M_AXIS_BRAM_56_ADDR_WIDTH-1:0] ap_bram_oarg_56_addr1,
    input [M_AXIS_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_din1,
    output [M_AXIS_BRAM_56_WIDTH-1:0] ap_bram_oarg_56_dout1,
    input ap_bram_oarg_56_clk1,
    input ap_bram_oarg_56_rst1,
    input [M_AXIS_BRAM_56_WIDTH/8-1:0] ap_bram_oarg_56_we1,
    input ap_bram_oarg_56_en1,
    //out BRAM to AXI-Stream interface 57
    input m_axis_bram_57_aclk,
    input m_axis_bram_57_aresetn,
    output m_axis_bram_57_tlast,
    output m_axis_bram_57_tvalid,
    output [M_AXIS_BRAM_57_DMWIDTH/8-1:0] m_axis_bram_57_tkeep,
    output [M_AXIS_BRAM_57_DMWIDTH/8-1:0] m_axis_bram_57_tstrb,
    output [M_AXIS_BRAM_57_DMWIDTH-1:0] m_axis_bram_57_tdata,
    input m_axis_bram_57_tready,
    input [M_AXIS_BRAM_57_ADDR_WIDTH-1:0] ap_bram_oarg_57_addr0,
    input [M_AXIS_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_din0,
    output [M_AXIS_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_dout0,
    input ap_bram_oarg_57_clk0,
    input ap_bram_oarg_57_rst0,
    input [M_AXIS_BRAM_57_WIDTH/8-1:0] ap_bram_oarg_57_we0,
    input ap_bram_oarg_57_en0,
    input [M_AXIS_BRAM_57_ADDR_WIDTH-1:0] ap_bram_oarg_57_addr1,
    input [M_AXIS_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_din1,
    output [M_AXIS_BRAM_57_WIDTH-1:0] ap_bram_oarg_57_dout1,
    input ap_bram_oarg_57_clk1,
    input ap_bram_oarg_57_rst1,
    input [M_AXIS_BRAM_57_WIDTH/8-1:0] ap_bram_oarg_57_we1,
    input ap_bram_oarg_57_en1,
    //out BRAM to AXI-Stream interface 58
    input m_axis_bram_58_aclk,
    input m_axis_bram_58_aresetn,
    output m_axis_bram_58_tlast,
    output m_axis_bram_58_tvalid,
    output [M_AXIS_BRAM_58_DMWIDTH/8-1:0] m_axis_bram_58_tkeep,
    output [M_AXIS_BRAM_58_DMWIDTH/8-1:0] m_axis_bram_58_tstrb,
    output [M_AXIS_BRAM_58_DMWIDTH-1:0] m_axis_bram_58_tdata,
    input m_axis_bram_58_tready,
    input [M_AXIS_BRAM_58_ADDR_WIDTH-1:0] ap_bram_oarg_58_addr0,
    input [M_AXIS_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_din0,
    output [M_AXIS_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_dout0,
    input ap_bram_oarg_58_clk0,
    input ap_bram_oarg_58_rst0,
    input [M_AXIS_BRAM_58_WIDTH/8-1:0] ap_bram_oarg_58_we0,
    input ap_bram_oarg_58_en0,
    input [M_AXIS_BRAM_58_ADDR_WIDTH-1:0] ap_bram_oarg_58_addr1,
    input [M_AXIS_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_din1,
    output [M_AXIS_BRAM_58_WIDTH-1:0] ap_bram_oarg_58_dout1,
    input ap_bram_oarg_58_clk1,
    input ap_bram_oarg_58_rst1,
    input [M_AXIS_BRAM_58_WIDTH/8-1:0] ap_bram_oarg_58_we1,
    input ap_bram_oarg_58_en1,
    //out BRAM to AXI-Stream interface 59
    input m_axis_bram_59_aclk,
    input m_axis_bram_59_aresetn,
    output m_axis_bram_59_tlast,
    output m_axis_bram_59_tvalid,
    output [M_AXIS_BRAM_59_DMWIDTH/8-1:0] m_axis_bram_59_tkeep,
    output [M_AXIS_BRAM_59_DMWIDTH/8-1:0] m_axis_bram_59_tstrb,
    output [M_AXIS_BRAM_59_DMWIDTH-1:0] m_axis_bram_59_tdata,
    input m_axis_bram_59_tready,
    input [M_AXIS_BRAM_59_ADDR_WIDTH-1:0] ap_bram_oarg_59_addr0,
    input [M_AXIS_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_din0,
    output [M_AXIS_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_dout0,
    input ap_bram_oarg_59_clk0,
    input ap_bram_oarg_59_rst0,
    input [M_AXIS_BRAM_59_WIDTH/8-1:0] ap_bram_oarg_59_we0,
    input ap_bram_oarg_59_en0,
    input [M_AXIS_BRAM_59_ADDR_WIDTH-1:0] ap_bram_oarg_59_addr1,
    input [M_AXIS_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_din1,
    output [M_AXIS_BRAM_59_WIDTH-1:0] ap_bram_oarg_59_dout1,
    input ap_bram_oarg_59_clk1,
    input ap_bram_oarg_59_rst1,
    input [M_AXIS_BRAM_59_WIDTH/8-1:0] ap_bram_oarg_59_we1,
    input ap_bram_oarg_59_en1,
    //out BRAM to AXI-Stream interface 60
    input m_axis_bram_60_aclk,
    input m_axis_bram_60_aresetn,
    output m_axis_bram_60_tlast,
    output m_axis_bram_60_tvalid,
    output [M_AXIS_BRAM_60_DMWIDTH/8-1:0] m_axis_bram_60_tkeep,
    output [M_AXIS_BRAM_60_DMWIDTH/8-1:0] m_axis_bram_60_tstrb,
    output [M_AXIS_BRAM_60_DMWIDTH-1:0] m_axis_bram_60_tdata,
    input m_axis_bram_60_tready,
    input [M_AXIS_BRAM_60_ADDR_WIDTH-1:0] ap_bram_oarg_60_addr0,
    input [M_AXIS_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_din0,
    output [M_AXIS_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_dout0,
    input ap_bram_oarg_60_clk0,
    input ap_bram_oarg_60_rst0,
    input [M_AXIS_BRAM_60_WIDTH/8-1:0] ap_bram_oarg_60_we0,
    input ap_bram_oarg_60_en0,
    input [M_AXIS_BRAM_60_ADDR_WIDTH-1:0] ap_bram_oarg_60_addr1,
    input [M_AXIS_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_din1,
    output [M_AXIS_BRAM_60_WIDTH-1:0] ap_bram_oarg_60_dout1,
    input ap_bram_oarg_60_clk1,
    input ap_bram_oarg_60_rst1,
    input [M_AXIS_BRAM_60_WIDTH/8-1:0] ap_bram_oarg_60_we1,
    input ap_bram_oarg_60_en1,
    //out BRAM to AXI-Stream interface 61
    input m_axis_bram_61_aclk,
    input m_axis_bram_61_aresetn,
    output m_axis_bram_61_tlast,
    output m_axis_bram_61_tvalid,
    output [M_AXIS_BRAM_61_DMWIDTH/8-1:0] m_axis_bram_61_tkeep,
    output [M_AXIS_BRAM_61_DMWIDTH/8-1:0] m_axis_bram_61_tstrb,
    output [M_AXIS_BRAM_61_DMWIDTH-1:0] m_axis_bram_61_tdata,
    input m_axis_bram_61_tready,
    input [M_AXIS_BRAM_61_ADDR_WIDTH-1:0] ap_bram_oarg_61_addr0,
    input [M_AXIS_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_din0,
    output [M_AXIS_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_dout0,
    input ap_bram_oarg_61_clk0,
    input ap_bram_oarg_61_rst0,
    input [M_AXIS_BRAM_61_WIDTH/8-1:0] ap_bram_oarg_61_we0,
    input ap_bram_oarg_61_en0,
    input [M_AXIS_BRAM_61_ADDR_WIDTH-1:0] ap_bram_oarg_61_addr1,
    input [M_AXIS_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_din1,
    output [M_AXIS_BRAM_61_WIDTH-1:0] ap_bram_oarg_61_dout1,
    input ap_bram_oarg_61_clk1,
    input ap_bram_oarg_61_rst1,
    input [M_AXIS_BRAM_61_WIDTH/8-1:0] ap_bram_oarg_61_we1,
    input ap_bram_oarg_61_en1,
    //out BRAM to AXI-Stream interface 62
    input m_axis_bram_62_aclk,
    input m_axis_bram_62_aresetn,
    output m_axis_bram_62_tlast,
    output m_axis_bram_62_tvalid,
    output [M_AXIS_BRAM_62_DMWIDTH/8-1:0] m_axis_bram_62_tkeep,
    output [M_AXIS_BRAM_62_DMWIDTH/8-1:0] m_axis_bram_62_tstrb,
    output [M_AXIS_BRAM_62_DMWIDTH-1:0] m_axis_bram_62_tdata,
    input m_axis_bram_62_tready,
    input [M_AXIS_BRAM_62_ADDR_WIDTH-1:0] ap_bram_oarg_62_addr0,
    input [M_AXIS_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_din0,
    output [M_AXIS_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_dout0,
    input ap_bram_oarg_62_clk0,
    input ap_bram_oarg_62_rst0,
    input [M_AXIS_BRAM_62_WIDTH/8-1:0] ap_bram_oarg_62_we0,
    input ap_bram_oarg_62_en0,
    input [M_AXIS_BRAM_62_ADDR_WIDTH-1:0] ap_bram_oarg_62_addr1,
    input [M_AXIS_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_din1,
    output [M_AXIS_BRAM_62_WIDTH-1:0] ap_bram_oarg_62_dout1,
    input ap_bram_oarg_62_clk1,
    input ap_bram_oarg_62_rst1,
    input [M_AXIS_BRAM_62_WIDTH/8-1:0] ap_bram_oarg_62_we1,
    input ap_bram_oarg_62_en1,
    //out BRAM to AXI-Stream interface 63
    input m_axis_bram_63_aclk,
    input m_axis_bram_63_aresetn,
    output m_axis_bram_63_tlast,
    output m_axis_bram_63_tvalid,
    output [M_AXIS_BRAM_63_DMWIDTH/8-1:0] m_axis_bram_63_tkeep,
    output [M_AXIS_BRAM_63_DMWIDTH/8-1:0] m_axis_bram_63_tstrb,
    output [M_AXIS_BRAM_63_DMWIDTH-1:0] m_axis_bram_63_tdata,
    input m_axis_bram_63_tready,
    input [M_AXIS_BRAM_63_ADDR_WIDTH-1:0] ap_bram_oarg_63_addr0,
    input [M_AXIS_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_din0,
    output [M_AXIS_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_dout0,
    input ap_bram_oarg_63_clk0,
    input ap_bram_oarg_63_rst0,
    input [M_AXIS_BRAM_63_WIDTH/8-1:0] ap_bram_oarg_63_we0,
    input ap_bram_oarg_63_en0,
    input [M_AXIS_BRAM_63_ADDR_WIDTH-1:0] ap_bram_oarg_63_addr1,
    input [M_AXIS_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_din1,
    output [M_AXIS_BRAM_63_WIDTH-1:0] ap_bram_oarg_63_dout1,
    input ap_bram_oarg_63_clk1,
    input ap_bram_oarg_63_rst1,
    input [M_AXIS_BRAM_63_WIDTH/8-1:0] ap_bram_oarg_63_we1,
    input ap_bram_oarg_63_en1,
    //out BRAM to AXI-Stream interface 64
    input m_axis_bram_64_aclk,
    input m_axis_bram_64_aresetn,
    output m_axis_bram_64_tlast,
    output m_axis_bram_64_tvalid,
    output [M_AXIS_BRAM_64_DMWIDTH/8-1:0] m_axis_bram_64_tkeep,
    output [M_AXIS_BRAM_64_DMWIDTH/8-1:0] m_axis_bram_64_tstrb,
    output [M_AXIS_BRAM_64_DMWIDTH-1:0] m_axis_bram_64_tdata,
    input m_axis_bram_64_tready,
    input [M_AXIS_BRAM_64_ADDR_WIDTH-1:0] ap_bram_oarg_64_addr0,
    input [M_AXIS_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_din0,
    output [M_AXIS_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_dout0,
    input ap_bram_oarg_64_clk0,
    input ap_bram_oarg_64_rst0,
    input [M_AXIS_BRAM_64_WIDTH/8-1:0] ap_bram_oarg_64_we0,
    input ap_bram_oarg_64_en0,
    input [M_AXIS_BRAM_64_ADDR_WIDTH-1:0] ap_bram_oarg_64_addr1,
    input [M_AXIS_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_din1,
    output [M_AXIS_BRAM_64_WIDTH-1:0] ap_bram_oarg_64_dout1,
    input ap_bram_oarg_64_clk1,
    input ap_bram_oarg_64_rst1,
    input [M_AXIS_BRAM_64_WIDTH/8-1:0] ap_bram_oarg_64_we1,
    input ap_bram_oarg_64_en1,
    //out BRAM to AXI-Stream interface 65
    input m_axis_bram_65_aclk,
    input m_axis_bram_65_aresetn,
    output m_axis_bram_65_tlast,
    output m_axis_bram_65_tvalid,
    output [M_AXIS_BRAM_65_DMWIDTH/8-1:0] m_axis_bram_65_tkeep,
    output [M_AXIS_BRAM_65_DMWIDTH/8-1:0] m_axis_bram_65_tstrb,
    output [M_AXIS_BRAM_65_DMWIDTH-1:0] m_axis_bram_65_tdata,
    input m_axis_bram_65_tready,
    input [M_AXIS_BRAM_65_ADDR_WIDTH-1:0] ap_bram_oarg_65_addr0,
    input [M_AXIS_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_din0,
    output [M_AXIS_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_dout0,
    input ap_bram_oarg_65_clk0,
    input ap_bram_oarg_65_rst0,
    input [M_AXIS_BRAM_65_WIDTH/8-1:0] ap_bram_oarg_65_we0,
    input ap_bram_oarg_65_en0,
    input [M_AXIS_BRAM_65_ADDR_WIDTH-1:0] ap_bram_oarg_65_addr1,
    input [M_AXIS_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_din1,
    output [M_AXIS_BRAM_65_WIDTH-1:0] ap_bram_oarg_65_dout1,
    input ap_bram_oarg_65_clk1,
    input ap_bram_oarg_65_rst1,
    input [M_AXIS_BRAM_65_WIDTH/8-1:0] ap_bram_oarg_65_we1,
    input ap_bram_oarg_65_en1,
    //out BRAM to AXI-Stream interface 66
    input m_axis_bram_66_aclk,
    input m_axis_bram_66_aresetn,
    output m_axis_bram_66_tlast,
    output m_axis_bram_66_tvalid,
    output [M_AXIS_BRAM_66_DMWIDTH/8-1:0] m_axis_bram_66_tkeep,
    output [M_AXIS_BRAM_66_DMWIDTH/8-1:0] m_axis_bram_66_tstrb,
    output [M_AXIS_BRAM_66_DMWIDTH-1:0] m_axis_bram_66_tdata,
    input m_axis_bram_66_tready,
    input [M_AXIS_BRAM_66_ADDR_WIDTH-1:0] ap_bram_oarg_66_addr0,
    input [M_AXIS_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_din0,
    output [M_AXIS_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_dout0,
    input ap_bram_oarg_66_clk0,
    input ap_bram_oarg_66_rst0,
    input [M_AXIS_BRAM_66_WIDTH/8-1:0] ap_bram_oarg_66_we0,
    input ap_bram_oarg_66_en0,
    input [M_AXIS_BRAM_66_ADDR_WIDTH-1:0] ap_bram_oarg_66_addr1,
    input [M_AXIS_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_din1,
    output [M_AXIS_BRAM_66_WIDTH-1:0] ap_bram_oarg_66_dout1,
    input ap_bram_oarg_66_clk1,
    input ap_bram_oarg_66_rst1,
    input [M_AXIS_BRAM_66_WIDTH/8-1:0] ap_bram_oarg_66_we1,
    input ap_bram_oarg_66_en1,
    //out BRAM to AXI-Stream interface 67
    input m_axis_bram_67_aclk,
    input m_axis_bram_67_aresetn,
    output m_axis_bram_67_tlast,
    output m_axis_bram_67_tvalid,
    output [M_AXIS_BRAM_67_DMWIDTH/8-1:0] m_axis_bram_67_tkeep,
    output [M_AXIS_BRAM_67_DMWIDTH/8-1:0] m_axis_bram_67_tstrb,
    output [M_AXIS_BRAM_67_DMWIDTH-1:0] m_axis_bram_67_tdata,
    input m_axis_bram_67_tready,
    input [M_AXIS_BRAM_67_ADDR_WIDTH-1:0] ap_bram_oarg_67_addr0,
    input [M_AXIS_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_din0,
    output [M_AXIS_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_dout0,
    input ap_bram_oarg_67_clk0,
    input ap_bram_oarg_67_rst0,
    input [M_AXIS_BRAM_67_WIDTH/8-1:0] ap_bram_oarg_67_we0,
    input ap_bram_oarg_67_en0,
    input [M_AXIS_BRAM_67_ADDR_WIDTH-1:0] ap_bram_oarg_67_addr1,
    input [M_AXIS_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_din1,
    output [M_AXIS_BRAM_67_WIDTH-1:0] ap_bram_oarg_67_dout1,
    input ap_bram_oarg_67_clk1,
    input ap_bram_oarg_67_rst1,
    input [M_AXIS_BRAM_67_WIDTH/8-1:0] ap_bram_oarg_67_we1,
    input ap_bram_oarg_67_en1,
    //out BRAM to AXI-Stream interface 68
    input m_axis_bram_68_aclk,
    input m_axis_bram_68_aresetn,
    output m_axis_bram_68_tlast,
    output m_axis_bram_68_tvalid,
    output [M_AXIS_BRAM_68_DMWIDTH/8-1:0] m_axis_bram_68_tkeep,
    output [M_AXIS_BRAM_68_DMWIDTH/8-1:0] m_axis_bram_68_tstrb,
    output [M_AXIS_BRAM_68_DMWIDTH-1:0] m_axis_bram_68_tdata,
    input m_axis_bram_68_tready,
    input [M_AXIS_BRAM_68_ADDR_WIDTH-1:0] ap_bram_oarg_68_addr0,
    input [M_AXIS_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_din0,
    output [M_AXIS_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_dout0,
    input ap_bram_oarg_68_clk0,
    input ap_bram_oarg_68_rst0,
    input [M_AXIS_BRAM_68_WIDTH/8-1:0] ap_bram_oarg_68_we0,
    input ap_bram_oarg_68_en0,
    input [M_AXIS_BRAM_68_ADDR_WIDTH-1:0] ap_bram_oarg_68_addr1,
    input [M_AXIS_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_din1,
    output [M_AXIS_BRAM_68_WIDTH-1:0] ap_bram_oarg_68_dout1,
    input ap_bram_oarg_68_clk1,
    input ap_bram_oarg_68_rst1,
    input [M_AXIS_BRAM_68_WIDTH/8-1:0] ap_bram_oarg_68_we1,
    input ap_bram_oarg_68_en1,
    //out BRAM to AXI-Stream interface 69
    input m_axis_bram_69_aclk,
    input m_axis_bram_69_aresetn,
    output m_axis_bram_69_tlast,
    output m_axis_bram_69_tvalid,
    output [M_AXIS_BRAM_69_DMWIDTH/8-1:0] m_axis_bram_69_tkeep,
    output [M_AXIS_BRAM_69_DMWIDTH/8-1:0] m_axis_bram_69_tstrb,
    output [M_AXIS_BRAM_69_DMWIDTH-1:0] m_axis_bram_69_tdata,
    input m_axis_bram_69_tready,
    input [M_AXIS_BRAM_69_ADDR_WIDTH-1:0] ap_bram_oarg_69_addr0,
    input [M_AXIS_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_din0,
    output [M_AXIS_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_dout0,
    input ap_bram_oarg_69_clk0,
    input ap_bram_oarg_69_rst0,
    input [M_AXIS_BRAM_69_WIDTH/8-1:0] ap_bram_oarg_69_we0,
    input ap_bram_oarg_69_en0,
    input [M_AXIS_BRAM_69_ADDR_WIDTH-1:0] ap_bram_oarg_69_addr1,
    input [M_AXIS_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_din1,
    output [M_AXIS_BRAM_69_WIDTH-1:0] ap_bram_oarg_69_dout1,
    input ap_bram_oarg_69_clk1,
    input ap_bram_oarg_69_rst1,
    input [M_AXIS_BRAM_69_WIDTH/8-1:0] ap_bram_oarg_69_we1,
    input ap_bram_oarg_69_en1,
    //out BRAM to AXI-Stream interface 70
    input m_axis_bram_70_aclk,
    input m_axis_bram_70_aresetn,
    output m_axis_bram_70_tlast,
    output m_axis_bram_70_tvalid,
    output [M_AXIS_BRAM_70_DMWIDTH/8-1:0] m_axis_bram_70_tkeep,
    output [M_AXIS_BRAM_70_DMWIDTH/8-1:0] m_axis_bram_70_tstrb,
    output [M_AXIS_BRAM_70_DMWIDTH-1:0] m_axis_bram_70_tdata,
    input m_axis_bram_70_tready,
    input [M_AXIS_BRAM_70_ADDR_WIDTH-1:0] ap_bram_oarg_70_addr0,
    input [M_AXIS_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_din0,
    output [M_AXIS_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_dout0,
    input ap_bram_oarg_70_clk0,
    input ap_bram_oarg_70_rst0,
    input [M_AXIS_BRAM_70_WIDTH/8-1:0] ap_bram_oarg_70_we0,
    input ap_bram_oarg_70_en0,
    input [M_AXIS_BRAM_70_ADDR_WIDTH-1:0] ap_bram_oarg_70_addr1,
    input [M_AXIS_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_din1,
    output [M_AXIS_BRAM_70_WIDTH-1:0] ap_bram_oarg_70_dout1,
    input ap_bram_oarg_70_clk1,
    input ap_bram_oarg_70_rst1,
    input [M_AXIS_BRAM_70_WIDTH/8-1:0] ap_bram_oarg_70_we1,
    input ap_bram_oarg_70_en1,
    //out BRAM to AXI-Stream interface 71
    input m_axis_bram_71_aclk,
    input m_axis_bram_71_aresetn,
    output m_axis_bram_71_tlast,
    output m_axis_bram_71_tvalid,
    output [M_AXIS_BRAM_71_DMWIDTH/8-1:0] m_axis_bram_71_tkeep,
    output [M_AXIS_BRAM_71_DMWIDTH/8-1:0] m_axis_bram_71_tstrb,
    output [M_AXIS_BRAM_71_DMWIDTH-1:0] m_axis_bram_71_tdata,
    input m_axis_bram_71_tready,
    input [M_AXIS_BRAM_71_ADDR_WIDTH-1:0] ap_bram_oarg_71_addr0,
    input [M_AXIS_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_din0,
    output [M_AXIS_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_dout0,
    input ap_bram_oarg_71_clk0,
    input ap_bram_oarg_71_rst0,
    input [M_AXIS_BRAM_71_WIDTH/8-1:0] ap_bram_oarg_71_we0,
    input ap_bram_oarg_71_en0,
    input [M_AXIS_BRAM_71_ADDR_WIDTH-1:0] ap_bram_oarg_71_addr1,
    input [M_AXIS_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_din1,
    output [M_AXIS_BRAM_71_WIDTH-1:0] ap_bram_oarg_71_dout1,
    input ap_bram_oarg_71_clk1,
    input ap_bram_oarg_71_rst1,
    input [M_AXIS_BRAM_71_WIDTH/8-1:0] ap_bram_oarg_71_we1,
    input ap_bram_oarg_71_en1,
    //out BRAM to AXI-Stream interface 72
    input m_axis_bram_72_aclk,
    input m_axis_bram_72_aresetn,
    output m_axis_bram_72_tlast,
    output m_axis_bram_72_tvalid,
    output [M_AXIS_BRAM_72_DMWIDTH/8-1:0] m_axis_bram_72_tkeep,
    output [M_AXIS_BRAM_72_DMWIDTH/8-1:0] m_axis_bram_72_tstrb,
    output [M_AXIS_BRAM_72_DMWIDTH-1:0] m_axis_bram_72_tdata,
    input m_axis_bram_72_tready,
    input [M_AXIS_BRAM_72_ADDR_WIDTH-1:0] ap_bram_oarg_72_addr0,
    input [M_AXIS_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_din0,
    output [M_AXIS_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_dout0,
    input ap_bram_oarg_72_clk0,
    input ap_bram_oarg_72_rst0,
    input [M_AXIS_BRAM_72_WIDTH/8-1:0] ap_bram_oarg_72_we0,
    input ap_bram_oarg_72_en0,
    input [M_AXIS_BRAM_72_ADDR_WIDTH-1:0] ap_bram_oarg_72_addr1,
    input [M_AXIS_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_din1,
    output [M_AXIS_BRAM_72_WIDTH-1:0] ap_bram_oarg_72_dout1,
    input ap_bram_oarg_72_clk1,
    input ap_bram_oarg_72_rst1,
    input [M_AXIS_BRAM_72_WIDTH/8-1:0] ap_bram_oarg_72_we1,
    input ap_bram_oarg_72_en1,
    //out BRAM to AXI-Stream interface 73
    input m_axis_bram_73_aclk,
    input m_axis_bram_73_aresetn,
    output m_axis_bram_73_tlast,
    output m_axis_bram_73_tvalid,
    output [M_AXIS_BRAM_73_DMWIDTH/8-1:0] m_axis_bram_73_tkeep,
    output [M_AXIS_BRAM_73_DMWIDTH/8-1:0] m_axis_bram_73_tstrb,
    output [M_AXIS_BRAM_73_DMWIDTH-1:0] m_axis_bram_73_tdata,
    input m_axis_bram_73_tready,
    input [M_AXIS_BRAM_73_ADDR_WIDTH-1:0] ap_bram_oarg_73_addr0,
    input [M_AXIS_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_din0,
    output [M_AXIS_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_dout0,
    input ap_bram_oarg_73_clk0,
    input ap_bram_oarg_73_rst0,
    input [M_AXIS_BRAM_73_WIDTH/8-1:0] ap_bram_oarg_73_we0,
    input ap_bram_oarg_73_en0,
    input [M_AXIS_BRAM_73_ADDR_WIDTH-1:0] ap_bram_oarg_73_addr1,
    input [M_AXIS_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_din1,
    output [M_AXIS_BRAM_73_WIDTH-1:0] ap_bram_oarg_73_dout1,
    input ap_bram_oarg_73_clk1,
    input ap_bram_oarg_73_rst1,
    input [M_AXIS_BRAM_73_WIDTH/8-1:0] ap_bram_oarg_73_we1,
    input ap_bram_oarg_73_en1,
    //out BRAM to AXI-Stream interface 74
    input m_axis_bram_74_aclk,
    input m_axis_bram_74_aresetn,
    output m_axis_bram_74_tlast,
    output m_axis_bram_74_tvalid,
    output [M_AXIS_BRAM_74_DMWIDTH/8-1:0] m_axis_bram_74_tkeep,
    output [M_AXIS_BRAM_74_DMWIDTH/8-1:0] m_axis_bram_74_tstrb,
    output [M_AXIS_BRAM_74_DMWIDTH-1:0] m_axis_bram_74_tdata,
    input m_axis_bram_74_tready,
    input [M_AXIS_BRAM_74_ADDR_WIDTH-1:0] ap_bram_oarg_74_addr0,
    input [M_AXIS_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_din0,
    output [M_AXIS_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_dout0,
    input ap_bram_oarg_74_clk0,
    input ap_bram_oarg_74_rst0,
    input [M_AXIS_BRAM_74_WIDTH/8-1:0] ap_bram_oarg_74_we0,
    input ap_bram_oarg_74_en0,
    input [M_AXIS_BRAM_74_ADDR_WIDTH-1:0] ap_bram_oarg_74_addr1,
    input [M_AXIS_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_din1,
    output [M_AXIS_BRAM_74_WIDTH-1:0] ap_bram_oarg_74_dout1,
    input ap_bram_oarg_74_clk1,
    input ap_bram_oarg_74_rst1,
    input [M_AXIS_BRAM_74_WIDTH/8-1:0] ap_bram_oarg_74_we1,
    input ap_bram_oarg_74_en1,
    //out BRAM to AXI-Stream interface 75
    input m_axis_bram_75_aclk,
    input m_axis_bram_75_aresetn,
    output m_axis_bram_75_tlast,
    output m_axis_bram_75_tvalid,
    output [M_AXIS_BRAM_75_DMWIDTH/8-1:0] m_axis_bram_75_tkeep,
    output [M_AXIS_BRAM_75_DMWIDTH/8-1:0] m_axis_bram_75_tstrb,
    output [M_AXIS_BRAM_75_DMWIDTH-1:0] m_axis_bram_75_tdata,
    input m_axis_bram_75_tready,
    input [M_AXIS_BRAM_75_ADDR_WIDTH-1:0] ap_bram_oarg_75_addr0,
    input [M_AXIS_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_din0,
    output [M_AXIS_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_dout0,
    input ap_bram_oarg_75_clk0,
    input ap_bram_oarg_75_rst0,
    input [M_AXIS_BRAM_75_WIDTH/8-1:0] ap_bram_oarg_75_we0,
    input ap_bram_oarg_75_en0,
    input [M_AXIS_BRAM_75_ADDR_WIDTH-1:0] ap_bram_oarg_75_addr1,
    input [M_AXIS_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_din1,
    output [M_AXIS_BRAM_75_WIDTH-1:0] ap_bram_oarg_75_dout1,
    input ap_bram_oarg_75_clk1,
    input ap_bram_oarg_75_rst1,
    input [M_AXIS_BRAM_75_WIDTH/8-1:0] ap_bram_oarg_75_we1,
    input ap_bram_oarg_75_en1,
    //out BRAM to AXI-Stream interface 76
    input m_axis_bram_76_aclk,
    input m_axis_bram_76_aresetn,
    output m_axis_bram_76_tlast,
    output m_axis_bram_76_tvalid,
    output [M_AXIS_BRAM_76_DMWIDTH/8-1:0] m_axis_bram_76_tkeep,
    output [M_AXIS_BRAM_76_DMWIDTH/8-1:0] m_axis_bram_76_tstrb,
    output [M_AXIS_BRAM_76_DMWIDTH-1:0] m_axis_bram_76_tdata,
    input m_axis_bram_76_tready,
    input [M_AXIS_BRAM_76_ADDR_WIDTH-1:0] ap_bram_oarg_76_addr0,
    input [M_AXIS_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_din0,
    output [M_AXIS_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_dout0,
    input ap_bram_oarg_76_clk0,
    input ap_bram_oarg_76_rst0,
    input [M_AXIS_BRAM_76_WIDTH/8-1:0] ap_bram_oarg_76_we0,
    input ap_bram_oarg_76_en0,
    input [M_AXIS_BRAM_76_ADDR_WIDTH-1:0] ap_bram_oarg_76_addr1,
    input [M_AXIS_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_din1,
    output [M_AXIS_BRAM_76_WIDTH-1:0] ap_bram_oarg_76_dout1,
    input ap_bram_oarg_76_clk1,
    input ap_bram_oarg_76_rst1,
    input [M_AXIS_BRAM_76_WIDTH/8-1:0] ap_bram_oarg_76_we1,
    input ap_bram_oarg_76_en1,
    //out BRAM to AXI-Stream interface 77
    input m_axis_bram_77_aclk,
    input m_axis_bram_77_aresetn,
    output m_axis_bram_77_tlast,
    output m_axis_bram_77_tvalid,
    output [M_AXIS_BRAM_77_DMWIDTH/8-1:0] m_axis_bram_77_tkeep,
    output [M_AXIS_BRAM_77_DMWIDTH/8-1:0] m_axis_bram_77_tstrb,
    output [M_AXIS_BRAM_77_DMWIDTH-1:0] m_axis_bram_77_tdata,
    input m_axis_bram_77_tready,
    input [M_AXIS_BRAM_77_ADDR_WIDTH-1:0] ap_bram_oarg_77_addr0,
    input [M_AXIS_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_din0,
    output [M_AXIS_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_dout0,
    input ap_bram_oarg_77_clk0,
    input ap_bram_oarg_77_rst0,
    input [M_AXIS_BRAM_77_WIDTH/8-1:0] ap_bram_oarg_77_we0,
    input ap_bram_oarg_77_en0,
    input [M_AXIS_BRAM_77_ADDR_WIDTH-1:0] ap_bram_oarg_77_addr1,
    input [M_AXIS_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_din1,
    output [M_AXIS_BRAM_77_WIDTH-1:0] ap_bram_oarg_77_dout1,
    input ap_bram_oarg_77_clk1,
    input ap_bram_oarg_77_rst1,
    input [M_AXIS_BRAM_77_WIDTH/8-1:0] ap_bram_oarg_77_we1,
    input ap_bram_oarg_77_en1,
    //out BRAM to AXI-Stream interface 78
    input m_axis_bram_78_aclk,
    input m_axis_bram_78_aresetn,
    output m_axis_bram_78_tlast,
    output m_axis_bram_78_tvalid,
    output [M_AXIS_BRAM_78_DMWIDTH/8-1:0] m_axis_bram_78_tkeep,
    output [M_AXIS_BRAM_78_DMWIDTH/8-1:0] m_axis_bram_78_tstrb,
    output [M_AXIS_BRAM_78_DMWIDTH-1:0] m_axis_bram_78_tdata,
    input m_axis_bram_78_tready,
    input [M_AXIS_BRAM_78_ADDR_WIDTH-1:0] ap_bram_oarg_78_addr0,
    input [M_AXIS_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_din0,
    output [M_AXIS_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_dout0,
    input ap_bram_oarg_78_clk0,
    input ap_bram_oarg_78_rst0,
    input [M_AXIS_BRAM_78_WIDTH/8-1:0] ap_bram_oarg_78_we0,
    input ap_bram_oarg_78_en0,
    input [M_AXIS_BRAM_78_ADDR_WIDTH-1:0] ap_bram_oarg_78_addr1,
    input [M_AXIS_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_din1,
    output [M_AXIS_BRAM_78_WIDTH-1:0] ap_bram_oarg_78_dout1,
    input ap_bram_oarg_78_clk1,
    input ap_bram_oarg_78_rst1,
    input [M_AXIS_BRAM_78_WIDTH/8-1:0] ap_bram_oarg_78_we1,
    input ap_bram_oarg_78_en1,
    //out BRAM to AXI-Stream interface 79
    input m_axis_bram_79_aclk,
    input m_axis_bram_79_aresetn,
    output m_axis_bram_79_tlast,
    output m_axis_bram_79_tvalid,
    output [M_AXIS_BRAM_79_DMWIDTH/8-1:0] m_axis_bram_79_tkeep,
    output [M_AXIS_BRAM_79_DMWIDTH/8-1:0] m_axis_bram_79_tstrb,
    output [M_AXIS_BRAM_79_DMWIDTH-1:0] m_axis_bram_79_tdata,
    input m_axis_bram_79_tready,
    input [M_AXIS_BRAM_79_ADDR_WIDTH-1:0] ap_bram_oarg_79_addr0,
    input [M_AXIS_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_din0,
    output [M_AXIS_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_dout0,
    input ap_bram_oarg_79_clk0,
    input ap_bram_oarg_79_rst0,
    input [M_AXIS_BRAM_79_WIDTH/8-1:0] ap_bram_oarg_79_we0,
    input ap_bram_oarg_79_en0,
    input [M_AXIS_BRAM_79_ADDR_WIDTH-1:0] ap_bram_oarg_79_addr1,
    input [M_AXIS_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_din1,
    output [M_AXIS_BRAM_79_WIDTH-1:0] ap_bram_oarg_79_dout1,
    input ap_bram_oarg_79_clk1,
    input ap_bram_oarg_79_rst1,
    input [M_AXIS_BRAM_79_WIDTH/8-1:0] ap_bram_oarg_79_we1,
    input ap_bram_oarg_79_en1,
    //out BRAM to AXI-Stream interface 80
    input m_axis_bram_80_aclk,
    input m_axis_bram_80_aresetn,
    output m_axis_bram_80_tlast,
    output m_axis_bram_80_tvalid,
    output [M_AXIS_BRAM_80_DMWIDTH/8-1:0] m_axis_bram_80_tkeep,
    output [M_AXIS_BRAM_80_DMWIDTH/8-1:0] m_axis_bram_80_tstrb,
    output [M_AXIS_BRAM_80_DMWIDTH-1:0] m_axis_bram_80_tdata,
    input m_axis_bram_80_tready,
    input [M_AXIS_BRAM_80_ADDR_WIDTH-1:0] ap_bram_oarg_80_addr0,
    input [M_AXIS_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_din0,
    output [M_AXIS_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_dout0,
    input ap_bram_oarg_80_clk0,
    input ap_bram_oarg_80_rst0,
    input [M_AXIS_BRAM_80_WIDTH/8-1:0] ap_bram_oarg_80_we0,
    input ap_bram_oarg_80_en0,
    input [M_AXIS_BRAM_80_ADDR_WIDTH-1:0] ap_bram_oarg_80_addr1,
    input [M_AXIS_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_din1,
    output [M_AXIS_BRAM_80_WIDTH-1:0] ap_bram_oarg_80_dout1,
    input ap_bram_oarg_80_clk1,
    input ap_bram_oarg_80_rst1,
    input [M_AXIS_BRAM_80_WIDTH/8-1:0] ap_bram_oarg_80_we1,
    input ap_bram_oarg_80_en1,
    //out BRAM to AXI-Stream interface 81
    input m_axis_bram_81_aclk,
    input m_axis_bram_81_aresetn,
    output m_axis_bram_81_tlast,
    output m_axis_bram_81_tvalid,
    output [M_AXIS_BRAM_81_DMWIDTH/8-1:0] m_axis_bram_81_tkeep,
    output [M_AXIS_BRAM_81_DMWIDTH/8-1:0] m_axis_bram_81_tstrb,
    output [M_AXIS_BRAM_81_DMWIDTH-1:0] m_axis_bram_81_tdata,
    input m_axis_bram_81_tready,
    input [M_AXIS_BRAM_81_ADDR_WIDTH-1:0] ap_bram_oarg_81_addr0,
    input [M_AXIS_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_din0,
    output [M_AXIS_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_dout0,
    input ap_bram_oarg_81_clk0,
    input ap_bram_oarg_81_rst0,
    input [M_AXIS_BRAM_81_WIDTH/8-1:0] ap_bram_oarg_81_we0,
    input ap_bram_oarg_81_en0,
    input [M_AXIS_BRAM_81_ADDR_WIDTH-1:0] ap_bram_oarg_81_addr1,
    input [M_AXIS_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_din1,
    output [M_AXIS_BRAM_81_WIDTH-1:0] ap_bram_oarg_81_dout1,
    input ap_bram_oarg_81_clk1,
    input ap_bram_oarg_81_rst1,
    input [M_AXIS_BRAM_81_WIDTH/8-1:0] ap_bram_oarg_81_we1,
    input ap_bram_oarg_81_en1,
    //out BRAM to AXI-Stream interface 82
    input m_axis_bram_82_aclk,
    input m_axis_bram_82_aresetn,
    output m_axis_bram_82_tlast,
    output m_axis_bram_82_tvalid,
    output [M_AXIS_BRAM_82_DMWIDTH/8-1:0] m_axis_bram_82_tkeep,
    output [M_AXIS_BRAM_82_DMWIDTH/8-1:0] m_axis_bram_82_tstrb,
    output [M_AXIS_BRAM_82_DMWIDTH-1:0] m_axis_bram_82_tdata,
    input m_axis_bram_82_tready,
    input [M_AXIS_BRAM_82_ADDR_WIDTH-1:0] ap_bram_oarg_82_addr0,
    input [M_AXIS_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_din0,
    output [M_AXIS_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_dout0,
    input ap_bram_oarg_82_clk0,
    input ap_bram_oarg_82_rst0,
    input [M_AXIS_BRAM_82_WIDTH/8-1:0] ap_bram_oarg_82_we0,
    input ap_bram_oarg_82_en0,
    input [M_AXIS_BRAM_82_ADDR_WIDTH-1:0] ap_bram_oarg_82_addr1,
    input [M_AXIS_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_din1,
    output [M_AXIS_BRAM_82_WIDTH-1:0] ap_bram_oarg_82_dout1,
    input ap_bram_oarg_82_clk1,
    input ap_bram_oarg_82_rst1,
    input [M_AXIS_BRAM_82_WIDTH/8-1:0] ap_bram_oarg_82_we1,
    input ap_bram_oarg_82_en1,
    //out BRAM to AXI-Stream interface 83
    input m_axis_bram_83_aclk,
    input m_axis_bram_83_aresetn,
    output m_axis_bram_83_tlast,
    output m_axis_bram_83_tvalid,
    output [M_AXIS_BRAM_83_DMWIDTH/8-1:0] m_axis_bram_83_tkeep,
    output [M_AXIS_BRAM_83_DMWIDTH/8-1:0] m_axis_bram_83_tstrb,
    output [M_AXIS_BRAM_83_DMWIDTH-1:0] m_axis_bram_83_tdata,
    input m_axis_bram_83_tready,
    input [M_AXIS_BRAM_83_ADDR_WIDTH-1:0] ap_bram_oarg_83_addr0,
    input [M_AXIS_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_din0,
    output [M_AXIS_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_dout0,
    input ap_bram_oarg_83_clk0,
    input ap_bram_oarg_83_rst0,
    input [M_AXIS_BRAM_83_WIDTH/8-1:0] ap_bram_oarg_83_we0,
    input ap_bram_oarg_83_en0,
    input [M_AXIS_BRAM_83_ADDR_WIDTH-1:0] ap_bram_oarg_83_addr1,
    input [M_AXIS_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_din1,
    output [M_AXIS_BRAM_83_WIDTH-1:0] ap_bram_oarg_83_dout1,
    input ap_bram_oarg_83_clk1,
    input ap_bram_oarg_83_rst1,
    input [M_AXIS_BRAM_83_WIDTH/8-1:0] ap_bram_oarg_83_we1,
    input ap_bram_oarg_83_en1,
    //out BRAM to AXI-Stream interface 84
    input m_axis_bram_84_aclk,
    input m_axis_bram_84_aresetn,
    output m_axis_bram_84_tlast,
    output m_axis_bram_84_tvalid,
    output [M_AXIS_BRAM_84_DMWIDTH/8-1:0] m_axis_bram_84_tkeep,
    output [M_AXIS_BRAM_84_DMWIDTH/8-1:0] m_axis_bram_84_tstrb,
    output [M_AXIS_BRAM_84_DMWIDTH-1:0] m_axis_bram_84_tdata,
    input m_axis_bram_84_tready,
    input [M_AXIS_BRAM_84_ADDR_WIDTH-1:0] ap_bram_oarg_84_addr0,
    input [M_AXIS_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_din0,
    output [M_AXIS_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_dout0,
    input ap_bram_oarg_84_clk0,
    input ap_bram_oarg_84_rst0,
    input [M_AXIS_BRAM_84_WIDTH/8-1:0] ap_bram_oarg_84_we0,
    input ap_bram_oarg_84_en0,
    input [M_AXIS_BRAM_84_ADDR_WIDTH-1:0] ap_bram_oarg_84_addr1,
    input [M_AXIS_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_din1,
    output [M_AXIS_BRAM_84_WIDTH-1:0] ap_bram_oarg_84_dout1,
    input ap_bram_oarg_84_clk1,
    input ap_bram_oarg_84_rst1,
    input [M_AXIS_BRAM_84_WIDTH/8-1:0] ap_bram_oarg_84_we1,
    input ap_bram_oarg_84_en1,
    //out BRAM to AXI-Stream interface 85
    input m_axis_bram_85_aclk,
    input m_axis_bram_85_aresetn,
    output m_axis_bram_85_tlast,
    output m_axis_bram_85_tvalid,
    output [M_AXIS_BRAM_85_DMWIDTH/8-1:0] m_axis_bram_85_tkeep,
    output [M_AXIS_BRAM_85_DMWIDTH/8-1:0] m_axis_bram_85_tstrb,
    output [M_AXIS_BRAM_85_DMWIDTH-1:0] m_axis_bram_85_tdata,
    input m_axis_bram_85_tready,
    input [M_AXIS_BRAM_85_ADDR_WIDTH-1:0] ap_bram_oarg_85_addr0,
    input [M_AXIS_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_din0,
    output [M_AXIS_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_dout0,
    input ap_bram_oarg_85_clk0,
    input ap_bram_oarg_85_rst0,
    input [M_AXIS_BRAM_85_WIDTH/8-1:0] ap_bram_oarg_85_we0,
    input ap_bram_oarg_85_en0,
    input [M_AXIS_BRAM_85_ADDR_WIDTH-1:0] ap_bram_oarg_85_addr1,
    input [M_AXIS_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_din1,
    output [M_AXIS_BRAM_85_WIDTH-1:0] ap_bram_oarg_85_dout1,
    input ap_bram_oarg_85_clk1,
    input ap_bram_oarg_85_rst1,
    input [M_AXIS_BRAM_85_WIDTH/8-1:0] ap_bram_oarg_85_we1,
    input ap_bram_oarg_85_en1,
    //out BRAM to AXI-Stream interface 86
    input m_axis_bram_86_aclk,
    input m_axis_bram_86_aresetn,
    output m_axis_bram_86_tlast,
    output m_axis_bram_86_tvalid,
    output [M_AXIS_BRAM_86_DMWIDTH/8-1:0] m_axis_bram_86_tkeep,
    output [M_AXIS_BRAM_86_DMWIDTH/8-1:0] m_axis_bram_86_tstrb,
    output [M_AXIS_BRAM_86_DMWIDTH-1:0] m_axis_bram_86_tdata,
    input m_axis_bram_86_tready,
    input [M_AXIS_BRAM_86_ADDR_WIDTH-1:0] ap_bram_oarg_86_addr0,
    input [M_AXIS_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_din0,
    output [M_AXIS_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_dout0,
    input ap_bram_oarg_86_clk0,
    input ap_bram_oarg_86_rst0,
    input [M_AXIS_BRAM_86_WIDTH/8-1:0] ap_bram_oarg_86_we0,
    input ap_bram_oarg_86_en0,
    input [M_AXIS_BRAM_86_ADDR_WIDTH-1:0] ap_bram_oarg_86_addr1,
    input [M_AXIS_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_din1,
    output [M_AXIS_BRAM_86_WIDTH-1:0] ap_bram_oarg_86_dout1,
    input ap_bram_oarg_86_clk1,
    input ap_bram_oarg_86_rst1,
    input [M_AXIS_BRAM_86_WIDTH/8-1:0] ap_bram_oarg_86_we1,
    input ap_bram_oarg_86_en1,
    //out BRAM to AXI-Stream interface 87
    input m_axis_bram_87_aclk,
    input m_axis_bram_87_aresetn,
    output m_axis_bram_87_tlast,
    output m_axis_bram_87_tvalid,
    output [M_AXIS_BRAM_87_DMWIDTH/8-1:0] m_axis_bram_87_tkeep,
    output [M_AXIS_BRAM_87_DMWIDTH/8-1:0] m_axis_bram_87_tstrb,
    output [M_AXIS_BRAM_87_DMWIDTH-1:0] m_axis_bram_87_tdata,
    input m_axis_bram_87_tready,
    input [M_AXIS_BRAM_87_ADDR_WIDTH-1:0] ap_bram_oarg_87_addr0,
    input [M_AXIS_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_din0,
    output [M_AXIS_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_dout0,
    input ap_bram_oarg_87_clk0,
    input ap_bram_oarg_87_rst0,
    input [M_AXIS_BRAM_87_WIDTH/8-1:0] ap_bram_oarg_87_we0,
    input ap_bram_oarg_87_en0,
    input [M_AXIS_BRAM_87_ADDR_WIDTH-1:0] ap_bram_oarg_87_addr1,
    input [M_AXIS_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_din1,
    output [M_AXIS_BRAM_87_WIDTH-1:0] ap_bram_oarg_87_dout1,
    input ap_bram_oarg_87_clk1,
    input ap_bram_oarg_87_rst1,
    input [M_AXIS_BRAM_87_WIDTH/8-1:0] ap_bram_oarg_87_we1,
    input ap_bram_oarg_87_en1,
    //out BRAM to AXI-Stream interface 88
    input m_axis_bram_88_aclk,
    input m_axis_bram_88_aresetn,
    output m_axis_bram_88_tlast,
    output m_axis_bram_88_tvalid,
    output [M_AXIS_BRAM_88_DMWIDTH/8-1:0] m_axis_bram_88_tkeep,
    output [M_AXIS_BRAM_88_DMWIDTH/8-1:0] m_axis_bram_88_tstrb,
    output [M_AXIS_BRAM_88_DMWIDTH-1:0] m_axis_bram_88_tdata,
    input m_axis_bram_88_tready,
    input [M_AXIS_BRAM_88_ADDR_WIDTH-1:0] ap_bram_oarg_88_addr0,
    input [M_AXIS_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_din0,
    output [M_AXIS_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_dout0,
    input ap_bram_oarg_88_clk0,
    input ap_bram_oarg_88_rst0,
    input [M_AXIS_BRAM_88_WIDTH/8-1:0] ap_bram_oarg_88_we0,
    input ap_bram_oarg_88_en0,
    input [M_AXIS_BRAM_88_ADDR_WIDTH-1:0] ap_bram_oarg_88_addr1,
    input [M_AXIS_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_din1,
    output [M_AXIS_BRAM_88_WIDTH-1:0] ap_bram_oarg_88_dout1,
    input ap_bram_oarg_88_clk1,
    input ap_bram_oarg_88_rst1,
    input [M_AXIS_BRAM_88_WIDTH/8-1:0] ap_bram_oarg_88_we1,
    input ap_bram_oarg_88_en1,
    //out BRAM to AXI-Stream interface 89
    input m_axis_bram_89_aclk,
    input m_axis_bram_89_aresetn,
    output m_axis_bram_89_tlast,
    output m_axis_bram_89_tvalid,
    output [M_AXIS_BRAM_89_DMWIDTH/8-1:0] m_axis_bram_89_tkeep,
    output [M_AXIS_BRAM_89_DMWIDTH/8-1:0] m_axis_bram_89_tstrb,
    output [M_AXIS_BRAM_89_DMWIDTH-1:0] m_axis_bram_89_tdata,
    input m_axis_bram_89_tready,
    input [M_AXIS_BRAM_89_ADDR_WIDTH-1:0] ap_bram_oarg_89_addr0,
    input [M_AXIS_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_din0,
    output [M_AXIS_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_dout0,
    input ap_bram_oarg_89_clk0,
    input ap_bram_oarg_89_rst0,
    input [M_AXIS_BRAM_89_WIDTH/8-1:0] ap_bram_oarg_89_we0,
    input ap_bram_oarg_89_en0,
    input [M_AXIS_BRAM_89_ADDR_WIDTH-1:0] ap_bram_oarg_89_addr1,
    input [M_AXIS_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_din1,
    output [M_AXIS_BRAM_89_WIDTH-1:0] ap_bram_oarg_89_dout1,
    input ap_bram_oarg_89_clk1,
    input ap_bram_oarg_89_rst1,
    input [M_AXIS_BRAM_89_WIDTH/8-1:0] ap_bram_oarg_89_we1,
    input ap_bram_oarg_89_en1,
    //out BRAM to AXI-Stream interface 90
    input m_axis_bram_90_aclk,
    input m_axis_bram_90_aresetn,
    output m_axis_bram_90_tlast,
    output m_axis_bram_90_tvalid,
    output [M_AXIS_BRAM_90_DMWIDTH/8-1:0] m_axis_bram_90_tkeep,
    output [M_AXIS_BRAM_90_DMWIDTH/8-1:0] m_axis_bram_90_tstrb,
    output [M_AXIS_BRAM_90_DMWIDTH-1:0] m_axis_bram_90_tdata,
    input m_axis_bram_90_tready,
    input [M_AXIS_BRAM_90_ADDR_WIDTH-1:0] ap_bram_oarg_90_addr0,
    input [M_AXIS_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_din0,
    output [M_AXIS_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_dout0,
    input ap_bram_oarg_90_clk0,
    input ap_bram_oarg_90_rst0,
    input [M_AXIS_BRAM_90_WIDTH/8-1:0] ap_bram_oarg_90_we0,
    input ap_bram_oarg_90_en0,
    input [M_AXIS_BRAM_90_ADDR_WIDTH-1:0] ap_bram_oarg_90_addr1,
    input [M_AXIS_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_din1,
    output [M_AXIS_BRAM_90_WIDTH-1:0] ap_bram_oarg_90_dout1,
    input ap_bram_oarg_90_clk1,
    input ap_bram_oarg_90_rst1,
    input [M_AXIS_BRAM_90_WIDTH/8-1:0] ap_bram_oarg_90_we1,
    input ap_bram_oarg_90_en1,
    //out BRAM to AXI-Stream interface 91
    input m_axis_bram_91_aclk,
    input m_axis_bram_91_aresetn,
    output m_axis_bram_91_tlast,
    output m_axis_bram_91_tvalid,
    output [M_AXIS_BRAM_91_DMWIDTH/8-1:0] m_axis_bram_91_tkeep,
    output [M_AXIS_BRAM_91_DMWIDTH/8-1:0] m_axis_bram_91_tstrb,
    output [M_AXIS_BRAM_91_DMWIDTH-1:0] m_axis_bram_91_tdata,
    input m_axis_bram_91_tready,
    input [M_AXIS_BRAM_91_ADDR_WIDTH-1:0] ap_bram_oarg_91_addr0,
    input [M_AXIS_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_din0,
    output [M_AXIS_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_dout0,
    input ap_bram_oarg_91_clk0,
    input ap_bram_oarg_91_rst0,
    input [M_AXIS_BRAM_91_WIDTH/8-1:0] ap_bram_oarg_91_we0,
    input ap_bram_oarg_91_en0,
    input [M_AXIS_BRAM_91_ADDR_WIDTH-1:0] ap_bram_oarg_91_addr1,
    input [M_AXIS_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_din1,
    output [M_AXIS_BRAM_91_WIDTH-1:0] ap_bram_oarg_91_dout1,
    input ap_bram_oarg_91_clk1,
    input ap_bram_oarg_91_rst1,
    input [M_AXIS_BRAM_91_WIDTH/8-1:0] ap_bram_oarg_91_we1,
    input ap_bram_oarg_91_en1,
    //out BRAM to AXI-Stream interface 92
    input m_axis_bram_92_aclk,
    input m_axis_bram_92_aresetn,
    output m_axis_bram_92_tlast,
    output m_axis_bram_92_tvalid,
    output [M_AXIS_BRAM_92_DMWIDTH/8-1:0] m_axis_bram_92_tkeep,
    output [M_AXIS_BRAM_92_DMWIDTH/8-1:0] m_axis_bram_92_tstrb,
    output [M_AXIS_BRAM_92_DMWIDTH-1:0] m_axis_bram_92_tdata,
    input m_axis_bram_92_tready,
    input [M_AXIS_BRAM_92_ADDR_WIDTH-1:0] ap_bram_oarg_92_addr0,
    input [M_AXIS_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_din0,
    output [M_AXIS_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_dout0,
    input ap_bram_oarg_92_clk0,
    input ap_bram_oarg_92_rst0,
    input [M_AXIS_BRAM_92_WIDTH/8-1:0] ap_bram_oarg_92_we0,
    input ap_bram_oarg_92_en0,
    input [M_AXIS_BRAM_92_ADDR_WIDTH-1:0] ap_bram_oarg_92_addr1,
    input [M_AXIS_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_din1,
    output [M_AXIS_BRAM_92_WIDTH-1:0] ap_bram_oarg_92_dout1,
    input ap_bram_oarg_92_clk1,
    input ap_bram_oarg_92_rst1,
    input [M_AXIS_BRAM_92_WIDTH/8-1:0] ap_bram_oarg_92_we1,
    input ap_bram_oarg_92_en1,
    //out BRAM to AXI-Stream interface 93
    input m_axis_bram_93_aclk,
    input m_axis_bram_93_aresetn,
    output m_axis_bram_93_tlast,
    output m_axis_bram_93_tvalid,
    output [M_AXIS_BRAM_93_DMWIDTH/8-1:0] m_axis_bram_93_tkeep,
    output [M_AXIS_BRAM_93_DMWIDTH/8-1:0] m_axis_bram_93_tstrb,
    output [M_AXIS_BRAM_93_DMWIDTH-1:0] m_axis_bram_93_tdata,
    input m_axis_bram_93_tready,
    input [M_AXIS_BRAM_93_ADDR_WIDTH-1:0] ap_bram_oarg_93_addr0,
    input [M_AXIS_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_din0,
    output [M_AXIS_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_dout0,
    input ap_bram_oarg_93_clk0,
    input ap_bram_oarg_93_rst0,
    input [M_AXIS_BRAM_93_WIDTH/8-1:0] ap_bram_oarg_93_we0,
    input ap_bram_oarg_93_en0,
    input [M_AXIS_BRAM_93_ADDR_WIDTH-1:0] ap_bram_oarg_93_addr1,
    input [M_AXIS_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_din1,
    output [M_AXIS_BRAM_93_WIDTH-1:0] ap_bram_oarg_93_dout1,
    input ap_bram_oarg_93_clk1,
    input ap_bram_oarg_93_rst1,
    input [M_AXIS_BRAM_93_WIDTH/8-1:0] ap_bram_oarg_93_we1,
    input ap_bram_oarg_93_en1,
    //out BRAM to AXI-Stream interface 94
    input m_axis_bram_94_aclk,
    input m_axis_bram_94_aresetn,
    output m_axis_bram_94_tlast,
    output m_axis_bram_94_tvalid,
    output [M_AXIS_BRAM_94_DMWIDTH/8-1:0] m_axis_bram_94_tkeep,
    output [M_AXIS_BRAM_94_DMWIDTH/8-1:0] m_axis_bram_94_tstrb,
    output [M_AXIS_BRAM_94_DMWIDTH-1:0] m_axis_bram_94_tdata,
    input m_axis_bram_94_tready,
    input [M_AXIS_BRAM_94_ADDR_WIDTH-1:0] ap_bram_oarg_94_addr0,
    input [M_AXIS_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_din0,
    output [M_AXIS_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_dout0,
    input ap_bram_oarg_94_clk0,
    input ap_bram_oarg_94_rst0,
    input [M_AXIS_BRAM_94_WIDTH/8-1:0] ap_bram_oarg_94_we0,
    input ap_bram_oarg_94_en0,
    input [M_AXIS_BRAM_94_ADDR_WIDTH-1:0] ap_bram_oarg_94_addr1,
    input [M_AXIS_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_din1,
    output [M_AXIS_BRAM_94_WIDTH-1:0] ap_bram_oarg_94_dout1,
    input ap_bram_oarg_94_clk1,
    input ap_bram_oarg_94_rst1,
    input [M_AXIS_BRAM_94_WIDTH/8-1:0] ap_bram_oarg_94_we1,
    input ap_bram_oarg_94_en1,
    //out BRAM to AXI-Stream interface 95
    input m_axis_bram_95_aclk,
    input m_axis_bram_95_aresetn,
    output m_axis_bram_95_tlast,
    output m_axis_bram_95_tvalid,
    output [M_AXIS_BRAM_95_DMWIDTH/8-1:0] m_axis_bram_95_tkeep,
    output [M_AXIS_BRAM_95_DMWIDTH/8-1:0] m_axis_bram_95_tstrb,
    output [M_AXIS_BRAM_95_DMWIDTH-1:0] m_axis_bram_95_tdata,
    input m_axis_bram_95_tready,
    input [M_AXIS_BRAM_95_ADDR_WIDTH-1:0] ap_bram_oarg_95_addr0,
    input [M_AXIS_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_din0,
    output [M_AXIS_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_dout0,
    input ap_bram_oarg_95_clk0,
    input ap_bram_oarg_95_rst0,
    input [M_AXIS_BRAM_95_WIDTH/8-1:0] ap_bram_oarg_95_we0,
    input ap_bram_oarg_95_en0,
    input [M_AXIS_BRAM_95_ADDR_WIDTH-1:0] ap_bram_oarg_95_addr1,
    input [M_AXIS_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_din1,
    output [M_AXIS_BRAM_95_WIDTH-1:0] ap_bram_oarg_95_dout1,
    input ap_bram_oarg_95_clk1,
    input ap_bram_oarg_95_rst1,
    input [M_AXIS_BRAM_95_WIDTH/8-1:0] ap_bram_oarg_95_we1,
    input ap_bram_oarg_95_en1,
    //out BRAM to AXI-Stream interface 96
    input m_axis_bram_96_aclk,
    input m_axis_bram_96_aresetn,
    output m_axis_bram_96_tlast,
    output m_axis_bram_96_tvalid,
    output [M_AXIS_BRAM_96_DMWIDTH/8-1:0] m_axis_bram_96_tkeep,
    output [M_AXIS_BRAM_96_DMWIDTH/8-1:0] m_axis_bram_96_tstrb,
    output [M_AXIS_BRAM_96_DMWIDTH-1:0] m_axis_bram_96_tdata,
    input m_axis_bram_96_tready,
    input [M_AXIS_BRAM_96_ADDR_WIDTH-1:0] ap_bram_oarg_96_addr0,
    input [M_AXIS_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_din0,
    output [M_AXIS_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_dout0,
    input ap_bram_oarg_96_clk0,
    input ap_bram_oarg_96_rst0,
    input [M_AXIS_BRAM_96_WIDTH/8-1:0] ap_bram_oarg_96_we0,
    input ap_bram_oarg_96_en0,
    input [M_AXIS_BRAM_96_ADDR_WIDTH-1:0] ap_bram_oarg_96_addr1,
    input [M_AXIS_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_din1,
    output [M_AXIS_BRAM_96_WIDTH-1:0] ap_bram_oarg_96_dout1,
    input ap_bram_oarg_96_clk1,
    input ap_bram_oarg_96_rst1,
    input [M_AXIS_BRAM_96_WIDTH/8-1:0] ap_bram_oarg_96_we1,
    input ap_bram_oarg_96_en1,
    //out BRAM to AXI-Stream interface 97
    input m_axis_bram_97_aclk,
    input m_axis_bram_97_aresetn,
    output m_axis_bram_97_tlast,
    output m_axis_bram_97_tvalid,
    output [M_AXIS_BRAM_97_DMWIDTH/8-1:0] m_axis_bram_97_tkeep,
    output [M_AXIS_BRAM_97_DMWIDTH/8-1:0] m_axis_bram_97_tstrb,
    output [M_AXIS_BRAM_97_DMWIDTH-1:0] m_axis_bram_97_tdata,
    input m_axis_bram_97_tready,
    input [M_AXIS_BRAM_97_ADDR_WIDTH-1:0] ap_bram_oarg_97_addr0,
    input [M_AXIS_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_din0,
    output [M_AXIS_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_dout0,
    input ap_bram_oarg_97_clk0,
    input ap_bram_oarg_97_rst0,
    input [M_AXIS_BRAM_97_WIDTH/8-1:0] ap_bram_oarg_97_we0,
    input ap_bram_oarg_97_en0,
    input [M_AXIS_BRAM_97_ADDR_WIDTH-1:0] ap_bram_oarg_97_addr1,
    input [M_AXIS_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_din1,
    output [M_AXIS_BRAM_97_WIDTH-1:0] ap_bram_oarg_97_dout1,
    input ap_bram_oarg_97_clk1,
    input ap_bram_oarg_97_rst1,
    input [M_AXIS_BRAM_97_WIDTH/8-1:0] ap_bram_oarg_97_we1,
    input ap_bram_oarg_97_en1,
    //out BRAM to AXI-Stream interface 98
    input m_axis_bram_98_aclk,
    input m_axis_bram_98_aresetn,
    output m_axis_bram_98_tlast,
    output m_axis_bram_98_tvalid,
    output [M_AXIS_BRAM_98_DMWIDTH/8-1:0] m_axis_bram_98_tkeep,
    output [M_AXIS_BRAM_98_DMWIDTH/8-1:0] m_axis_bram_98_tstrb,
    output [M_AXIS_BRAM_98_DMWIDTH-1:0] m_axis_bram_98_tdata,
    input m_axis_bram_98_tready,
    input [M_AXIS_BRAM_98_ADDR_WIDTH-1:0] ap_bram_oarg_98_addr0,
    input [M_AXIS_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_din0,
    output [M_AXIS_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_dout0,
    input ap_bram_oarg_98_clk0,
    input ap_bram_oarg_98_rst0,
    input [M_AXIS_BRAM_98_WIDTH/8-1:0] ap_bram_oarg_98_we0,
    input ap_bram_oarg_98_en0,
    input [M_AXIS_BRAM_98_ADDR_WIDTH-1:0] ap_bram_oarg_98_addr1,
    input [M_AXIS_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_din1,
    output [M_AXIS_BRAM_98_WIDTH-1:0] ap_bram_oarg_98_dout1,
    input ap_bram_oarg_98_clk1,
    input ap_bram_oarg_98_rst1,
    input [M_AXIS_BRAM_98_WIDTH/8-1:0] ap_bram_oarg_98_we1,
    input ap_bram_oarg_98_en1,
    //out BRAM to AXI-Stream interface 99
    input m_axis_bram_99_aclk,
    input m_axis_bram_99_aresetn,
    output m_axis_bram_99_tlast,
    output m_axis_bram_99_tvalid,
    output [M_AXIS_BRAM_99_DMWIDTH/8-1:0] m_axis_bram_99_tkeep,
    output [M_AXIS_BRAM_99_DMWIDTH/8-1:0] m_axis_bram_99_tstrb,
    output [M_AXIS_BRAM_99_DMWIDTH-1:0] m_axis_bram_99_tdata,
    input m_axis_bram_99_tready,
    input [M_AXIS_BRAM_99_ADDR_WIDTH-1:0] ap_bram_oarg_99_addr0,
    input [M_AXIS_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_din0,
    output [M_AXIS_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_dout0,
    input ap_bram_oarg_99_clk0,
    input ap_bram_oarg_99_rst0,
    input [M_AXIS_BRAM_99_WIDTH/8-1:0] ap_bram_oarg_99_we0,
    input ap_bram_oarg_99_en0,
    input [M_AXIS_BRAM_99_ADDR_WIDTH-1:0] ap_bram_oarg_99_addr1,
    input [M_AXIS_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_din1,
    output [M_AXIS_BRAM_99_WIDTH-1:0] ap_bram_oarg_99_dout1,
    input ap_bram_oarg_99_clk1,
    input ap_bram_oarg_99_rst1,
    input [M_AXIS_BRAM_99_WIDTH/8-1:0] ap_bram_oarg_99_we1,
    input ap_bram_oarg_99_en1,
    //out BRAM to AXI-Stream interface 100
    input m_axis_bram_100_aclk,
    input m_axis_bram_100_aresetn,
    output m_axis_bram_100_tlast,
    output m_axis_bram_100_tvalid,
    output [M_AXIS_BRAM_100_DMWIDTH/8-1:0] m_axis_bram_100_tkeep,
    output [M_AXIS_BRAM_100_DMWIDTH/8-1:0] m_axis_bram_100_tstrb,
    output [M_AXIS_BRAM_100_DMWIDTH-1:0] m_axis_bram_100_tdata,
    input m_axis_bram_100_tready,
    input [M_AXIS_BRAM_100_ADDR_WIDTH-1:0] ap_bram_oarg_100_addr0,
    input [M_AXIS_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_din0,
    output [M_AXIS_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_dout0,
    input ap_bram_oarg_100_clk0,
    input ap_bram_oarg_100_rst0,
    input [M_AXIS_BRAM_100_WIDTH/8-1:0] ap_bram_oarg_100_we0,
    input ap_bram_oarg_100_en0,
    input [M_AXIS_BRAM_100_ADDR_WIDTH-1:0] ap_bram_oarg_100_addr1,
    input [M_AXIS_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_din1,
    output [M_AXIS_BRAM_100_WIDTH-1:0] ap_bram_oarg_100_dout1,
    input ap_bram_oarg_100_clk1,
    input ap_bram_oarg_100_rst1,
    input [M_AXIS_BRAM_100_WIDTH/8-1:0] ap_bram_oarg_100_we1,
    input ap_bram_oarg_100_en1,
    //out BRAM to AXI-Stream interface 101
    input m_axis_bram_101_aclk,
    input m_axis_bram_101_aresetn,
    output m_axis_bram_101_tlast,
    output m_axis_bram_101_tvalid,
    output [M_AXIS_BRAM_101_DMWIDTH/8-1:0] m_axis_bram_101_tkeep,
    output [M_AXIS_BRAM_101_DMWIDTH/8-1:0] m_axis_bram_101_tstrb,
    output [M_AXIS_BRAM_101_DMWIDTH-1:0] m_axis_bram_101_tdata,
    input m_axis_bram_101_tready,
    input [M_AXIS_BRAM_101_ADDR_WIDTH-1:0] ap_bram_oarg_101_addr0,
    input [M_AXIS_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_din0,
    output [M_AXIS_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_dout0,
    input ap_bram_oarg_101_clk0,
    input ap_bram_oarg_101_rst0,
    input [M_AXIS_BRAM_101_WIDTH/8-1:0] ap_bram_oarg_101_we0,
    input ap_bram_oarg_101_en0,
    input [M_AXIS_BRAM_101_ADDR_WIDTH-1:0] ap_bram_oarg_101_addr1,
    input [M_AXIS_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_din1,
    output [M_AXIS_BRAM_101_WIDTH-1:0] ap_bram_oarg_101_dout1,
    input ap_bram_oarg_101_clk1,
    input ap_bram_oarg_101_rst1,
    input [M_AXIS_BRAM_101_WIDTH/8-1:0] ap_bram_oarg_101_we1,
    input ap_bram_oarg_101_en1,
    //out BRAM to AXI-Stream interface 102
    input m_axis_bram_102_aclk,
    input m_axis_bram_102_aresetn,
    output m_axis_bram_102_tlast,
    output m_axis_bram_102_tvalid,
    output [M_AXIS_BRAM_102_DMWIDTH/8-1:0] m_axis_bram_102_tkeep,
    output [M_AXIS_BRAM_102_DMWIDTH/8-1:0] m_axis_bram_102_tstrb,
    output [M_AXIS_BRAM_102_DMWIDTH-1:0] m_axis_bram_102_tdata,
    input m_axis_bram_102_tready,
    input [M_AXIS_BRAM_102_ADDR_WIDTH-1:0] ap_bram_oarg_102_addr0,
    input [M_AXIS_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_din0,
    output [M_AXIS_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_dout0,
    input ap_bram_oarg_102_clk0,
    input ap_bram_oarg_102_rst0,
    input [M_AXIS_BRAM_102_WIDTH/8-1:0] ap_bram_oarg_102_we0,
    input ap_bram_oarg_102_en0,
    input [M_AXIS_BRAM_102_ADDR_WIDTH-1:0] ap_bram_oarg_102_addr1,
    input [M_AXIS_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_din1,
    output [M_AXIS_BRAM_102_WIDTH-1:0] ap_bram_oarg_102_dout1,
    input ap_bram_oarg_102_clk1,
    input ap_bram_oarg_102_rst1,
    input [M_AXIS_BRAM_102_WIDTH/8-1:0] ap_bram_oarg_102_we1,
    input ap_bram_oarg_102_en1,
    //out BRAM to AXI-Stream interface 103
    input m_axis_bram_103_aclk,
    input m_axis_bram_103_aresetn,
    output m_axis_bram_103_tlast,
    output m_axis_bram_103_tvalid,
    output [M_AXIS_BRAM_103_DMWIDTH/8-1:0] m_axis_bram_103_tkeep,
    output [M_AXIS_BRAM_103_DMWIDTH/8-1:0] m_axis_bram_103_tstrb,
    output [M_AXIS_BRAM_103_DMWIDTH-1:0] m_axis_bram_103_tdata,
    input m_axis_bram_103_tready,
    input [M_AXIS_BRAM_103_ADDR_WIDTH-1:0] ap_bram_oarg_103_addr0,
    input [M_AXIS_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_din0,
    output [M_AXIS_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_dout0,
    input ap_bram_oarg_103_clk0,
    input ap_bram_oarg_103_rst0,
    input [M_AXIS_BRAM_103_WIDTH/8-1:0] ap_bram_oarg_103_we0,
    input ap_bram_oarg_103_en0,
    input [M_AXIS_BRAM_103_ADDR_WIDTH-1:0] ap_bram_oarg_103_addr1,
    input [M_AXIS_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_din1,
    output [M_AXIS_BRAM_103_WIDTH-1:0] ap_bram_oarg_103_dout1,
    input ap_bram_oarg_103_clk1,
    input ap_bram_oarg_103_rst1,
    input [M_AXIS_BRAM_103_WIDTH/8-1:0] ap_bram_oarg_103_we1,
    input ap_bram_oarg_103_en1,
    //out BRAM to AXI-Stream interface 104
    input m_axis_bram_104_aclk,
    input m_axis_bram_104_aresetn,
    output m_axis_bram_104_tlast,
    output m_axis_bram_104_tvalid,
    output [M_AXIS_BRAM_104_DMWIDTH/8-1:0] m_axis_bram_104_tkeep,
    output [M_AXIS_BRAM_104_DMWIDTH/8-1:0] m_axis_bram_104_tstrb,
    output [M_AXIS_BRAM_104_DMWIDTH-1:0] m_axis_bram_104_tdata,
    input m_axis_bram_104_tready,
    input [M_AXIS_BRAM_104_ADDR_WIDTH-1:0] ap_bram_oarg_104_addr0,
    input [M_AXIS_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_din0,
    output [M_AXIS_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_dout0,
    input ap_bram_oarg_104_clk0,
    input ap_bram_oarg_104_rst0,
    input [M_AXIS_BRAM_104_WIDTH/8-1:0] ap_bram_oarg_104_we0,
    input ap_bram_oarg_104_en0,
    input [M_AXIS_BRAM_104_ADDR_WIDTH-1:0] ap_bram_oarg_104_addr1,
    input [M_AXIS_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_din1,
    output [M_AXIS_BRAM_104_WIDTH-1:0] ap_bram_oarg_104_dout1,
    input ap_bram_oarg_104_clk1,
    input ap_bram_oarg_104_rst1,
    input [M_AXIS_BRAM_104_WIDTH/8-1:0] ap_bram_oarg_104_we1,
    input ap_bram_oarg_104_en1,
    //out BRAM to AXI-Stream interface 105
    input m_axis_bram_105_aclk,
    input m_axis_bram_105_aresetn,
    output m_axis_bram_105_tlast,
    output m_axis_bram_105_tvalid,
    output [M_AXIS_BRAM_105_DMWIDTH/8-1:0] m_axis_bram_105_tkeep,
    output [M_AXIS_BRAM_105_DMWIDTH/8-1:0] m_axis_bram_105_tstrb,
    output [M_AXIS_BRAM_105_DMWIDTH-1:0] m_axis_bram_105_tdata,
    input m_axis_bram_105_tready,
    input [M_AXIS_BRAM_105_ADDR_WIDTH-1:0] ap_bram_oarg_105_addr0,
    input [M_AXIS_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_din0,
    output [M_AXIS_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_dout0,
    input ap_bram_oarg_105_clk0,
    input ap_bram_oarg_105_rst0,
    input [M_AXIS_BRAM_105_WIDTH/8-1:0] ap_bram_oarg_105_we0,
    input ap_bram_oarg_105_en0,
    input [M_AXIS_BRAM_105_ADDR_WIDTH-1:0] ap_bram_oarg_105_addr1,
    input [M_AXIS_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_din1,
    output [M_AXIS_BRAM_105_WIDTH-1:0] ap_bram_oarg_105_dout1,
    input ap_bram_oarg_105_clk1,
    input ap_bram_oarg_105_rst1,
    input [M_AXIS_BRAM_105_WIDTH/8-1:0] ap_bram_oarg_105_we1,
    input ap_bram_oarg_105_en1,
    //out BRAM to AXI-Stream interface 106
    input m_axis_bram_106_aclk,
    input m_axis_bram_106_aresetn,
    output m_axis_bram_106_tlast,
    output m_axis_bram_106_tvalid,
    output [M_AXIS_BRAM_106_DMWIDTH/8-1:0] m_axis_bram_106_tkeep,
    output [M_AXIS_BRAM_106_DMWIDTH/8-1:0] m_axis_bram_106_tstrb,
    output [M_AXIS_BRAM_106_DMWIDTH-1:0] m_axis_bram_106_tdata,
    input m_axis_bram_106_tready,
    input [M_AXIS_BRAM_106_ADDR_WIDTH-1:0] ap_bram_oarg_106_addr0,
    input [M_AXIS_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_din0,
    output [M_AXIS_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_dout0,
    input ap_bram_oarg_106_clk0,
    input ap_bram_oarg_106_rst0,
    input [M_AXIS_BRAM_106_WIDTH/8-1:0] ap_bram_oarg_106_we0,
    input ap_bram_oarg_106_en0,
    input [M_AXIS_BRAM_106_ADDR_WIDTH-1:0] ap_bram_oarg_106_addr1,
    input [M_AXIS_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_din1,
    output [M_AXIS_BRAM_106_WIDTH-1:0] ap_bram_oarg_106_dout1,
    input ap_bram_oarg_106_clk1,
    input ap_bram_oarg_106_rst1,
    input [M_AXIS_BRAM_106_WIDTH/8-1:0] ap_bram_oarg_106_we1,
    input ap_bram_oarg_106_en1,
    //out BRAM to AXI-Stream interface 107
    input m_axis_bram_107_aclk,
    input m_axis_bram_107_aresetn,
    output m_axis_bram_107_tlast,
    output m_axis_bram_107_tvalid,
    output [M_AXIS_BRAM_107_DMWIDTH/8-1:0] m_axis_bram_107_tkeep,
    output [M_AXIS_BRAM_107_DMWIDTH/8-1:0] m_axis_bram_107_tstrb,
    output [M_AXIS_BRAM_107_DMWIDTH-1:0] m_axis_bram_107_tdata,
    input m_axis_bram_107_tready,
    input [M_AXIS_BRAM_107_ADDR_WIDTH-1:0] ap_bram_oarg_107_addr0,
    input [M_AXIS_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_din0,
    output [M_AXIS_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_dout0,
    input ap_bram_oarg_107_clk0,
    input ap_bram_oarg_107_rst0,
    input [M_AXIS_BRAM_107_WIDTH/8-1:0] ap_bram_oarg_107_we0,
    input ap_bram_oarg_107_en0,
    input [M_AXIS_BRAM_107_ADDR_WIDTH-1:0] ap_bram_oarg_107_addr1,
    input [M_AXIS_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_din1,
    output [M_AXIS_BRAM_107_WIDTH-1:0] ap_bram_oarg_107_dout1,
    input ap_bram_oarg_107_clk1,
    input ap_bram_oarg_107_rst1,
    input [M_AXIS_BRAM_107_WIDTH/8-1:0] ap_bram_oarg_107_we1,
    input ap_bram_oarg_107_en1,
    //out BRAM to AXI-Stream interface 108
    input m_axis_bram_108_aclk,
    input m_axis_bram_108_aresetn,
    output m_axis_bram_108_tlast,
    output m_axis_bram_108_tvalid,
    output [M_AXIS_BRAM_108_DMWIDTH/8-1:0] m_axis_bram_108_tkeep,
    output [M_AXIS_BRAM_108_DMWIDTH/8-1:0] m_axis_bram_108_tstrb,
    output [M_AXIS_BRAM_108_DMWIDTH-1:0] m_axis_bram_108_tdata,
    input m_axis_bram_108_tready,
    input [M_AXIS_BRAM_108_ADDR_WIDTH-1:0] ap_bram_oarg_108_addr0,
    input [M_AXIS_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_din0,
    output [M_AXIS_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_dout0,
    input ap_bram_oarg_108_clk0,
    input ap_bram_oarg_108_rst0,
    input [M_AXIS_BRAM_108_WIDTH/8-1:0] ap_bram_oarg_108_we0,
    input ap_bram_oarg_108_en0,
    input [M_AXIS_BRAM_108_ADDR_WIDTH-1:0] ap_bram_oarg_108_addr1,
    input [M_AXIS_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_din1,
    output [M_AXIS_BRAM_108_WIDTH-1:0] ap_bram_oarg_108_dout1,
    input ap_bram_oarg_108_clk1,
    input ap_bram_oarg_108_rst1,
    input [M_AXIS_BRAM_108_WIDTH/8-1:0] ap_bram_oarg_108_we1,
    input ap_bram_oarg_108_en1,
    //out BRAM to AXI-Stream interface 109
    input m_axis_bram_109_aclk,
    input m_axis_bram_109_aresetn,
    output m_axis_bram_109_tlast,
    output m_axis_bram_109_tvalid,
    output [M_AXIS_BRAM_109_DMWIDTH/8-1:0] m_axis_bram_109_tkeep,
    output [M_AXIS_BRAM_109_DMWIDTH/8-1:0] m_axis_bram_109_tstrb,
    output [M_AXIS_BRAM_109_DMWIDTH-1:0] m_axis_bram_109_tdata,
    input m_axis_bram_109_tready,
    input [M_AXIS_BRAM_109_ADDR_WIDTH-1:0] ap_bram_oarg_109_addr0,
    input [M_AXIS_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_din0,
    output [M_AXIS_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_dout0,
    input ap_bram_oarg_109_clk0,
    input ap_bram_oarg_109_rst0,
    input [M_AXIS_BRAM_109_WIDTH/8-1:0] ap_bram_oarg_109_we0,
    input ap_bram_oarg_109_en0,
    input [M_AXIS_BRAM_109_ADDR_WIDTH-1:0] ap_bram_oarg_109_addr1,
    input [M_AXIS_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_din1,
    output [M_AXIS_BRAM_109_WIDTH-1:0] ap_bram_oarg_109_dout1,
    input ap_bram_oarg_109_clk1,
    input ap_bram_oarg_109_rst1,
    input [M_AXIS_BRAM_109_WIDTH/8-1:0] ap_bram_oarg_109_we1,
    input ap_bram_oarg_109_en1,
    //out BRAM to AXI-Stream interface 110
    input m_axis_bram_110_aclk,
    input m_axis_bram_110_aresetn,
    output m_axis_bram_110_tlast,
    output m_axis_bram_110_tvalid,
    output [M_AXIS_BRAM_110_DMWIDTH/8-1:0] m_axis_bram_110_tkeep,
    output [M_AXIS_BRAM_110_DMWIDTH/8-1:0] m_axis_bram_110_tstrb,
    output [M_AXIS_BRAM_110_DMWIDTH-1:0] m_axis_bram_110_tdata,
    input m_axis_bram_110_tready,
    input [M_AXIS_BRAM_110_ADDR_WIDTH-1:0] ap_bram_oarg_110_addr0,
    input [M_AXIS_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_din0,
    output [M_AXIS_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_dout0,
    input ap_bram_oarg_110_clk0,
    input ap_bram_oarg_110_rst0,
    input [M_AXIS_BRAM_110_WIDTH/8-1:0] ap_bram_oarg_110_we0,
    input ap_bram_oarg_110_en0,
    input [M_AXIS_BRAM_110_ADDR_WIDTH-1:0] ap_bram_oarg_110_addr1,
    input [M_AXIS_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_din1,
    output [M_AXIS_BRAM_110_WIDTH-1:0] ap_bram_oarg_110_dout1,
    input ap_bram_oarg_110_clk1,
    input ap_bram_oarg_110_rst1,
    input [M_AXIS_BRAM_110_WIDTH/8-1:0] ap_bram_oarg_110_we1,
    input ap_bram_oarg_110_en1,
    //out BRAM to AXI-Stream interface 111
    input m_axis_bram_111_aclk,
    input m_axis_bram_111_aresetn,
    output m_axis_bram_111_tlast,
    output m_axis_bram_111_tvalid,
    output [M_AXIS_BRAM_111_DMWIDTH/8-1:0] m_axis_bram_111_tkeep,
    output [M_AXIS_BRAM_111_DMWIDTH/8-1:0] m_axis_bram_111_tstrb,
    output [M_AXIS_BRAM_111_DMWIDTH-1:0] m_axis_bram_111_tdata,
    input m_axis_bram_111_tready,
    input [M_AXIS_BRAM_111_ADDR_WIDTH-1:0] ap_bram_oarg_111_addr0,
    input [M_AXIS_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_din0,
    output [M_AXIS_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_dout0,
    input ap_bram_oarg_111_clk0,
    input ap_bram_oarg_111_rst0,
    input [M_AXIS_BRAM_111_WIDTH/8-1:0] ap_bram_oarg_111_we0,
    input ap_bram_oarg_111_en0,
    input [M_AXIS_BRAM_111_ADDR_WIDTH-1:0] ap_bram_oarg_111_addr1,
    input [M_AXIS_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_din1,
    output [M_AXIS_BRAM_111_WIDTH-1:0] ap_bram_oarg_111_dout1,
    input ap_bram_oarg_111_clk1,
    input ap_bram_oarg_111_rst1,
    input [M_AXIS_BRAM_111_WIDTH/8-1:0] ap_bram_oarg_111_we1,
    input ap_bram_oarg_111_en1,
    //out BRAM to AXI-Stream interface 112
    input m_axis_bram_112_aclk,
    input m_axis_bram_112_aresetn,
    output m_axis_bram_112_tlast,
    output m_axis_bram_112_tvalid,
    output [M_AXIS_BRAM_112_DMWIDTH/8-1:0] m_axis_bram_112_tkeep,
    output [M_AXIS_BRAM_112_DMWIDTH/8-1:0] m_axis_bram_112_tstrb,
    output [M_AXIS_BRAM_112_DMWIDTH-1:0] m_axis_bram_112_tdata,
    input m_axis_bram_112_tready,
    input [M_AXIS_BRAM_112_ADDR_WIDTH-1:0] ap_bram_oarg_112_addr0,
    input [M_AXIS_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_din0,
    output [M_AXIS_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_dout0,
    input ap_bram_oarg_112_clk0,
    input ap_bram_oarg_112_rst0,
    input [M_AXIS_BRAM_112_WIDTH/8-1:0] ap_bram_oarg_112_we0,
    input ap_bram_oarg_112_en0,
    input [M_AXIS_BRAM_112_ADDR_WIDTH-1:0] ap_bram_oarg_112_addr1,
    input [M_AXIS_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_din1,
    output [M_AXIS_BRAM_112_WIDTH-1:0] ap_bram_oarg_112_dout1,
    input ap_bram_oarg_112_clk1,
    input ap_bram_oarg_112_rst1,
    input [M_AXIS_BRAM_112_WIDTH/8-1:0] ap_bram_oarg_112_we1,
    input ap_bram_oarg_112_en1,
    //out BRAM to AXI-Stream interface 113
    input m_axis_bram_113_aclk,
    input m_axis_bram_113_aresetn,
    output m_axis_bram_113_tlast,
    output m_axis_bram_113_tvalid,
    output [M_AXIS_BRAM_113_DMWIDTH/8-1:0] m_axis_bram_113_tkeep,
    output [M_AXIS_BRAM_113_DMWIDTH/8-1:0] m_axis_bram_113_tstrb,
    output [M_AXIS_BRAM_113_DMWIDTH-1:0] m_axis_bram_113_tdata,
    input m_axis_bram_113_tready,
    input [M_AXIS_BRAM_113_ADDR_WIDTH-1:0] ap_bram_oarg_113_addr0,
    input [M_AXIS_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_din0,
    output [M_AXIS_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_dout0,
    input ap_bram_oarg_113_clk0,
    input ap_bram_oarg_113_rst0,
    input [M_AXIS_BRAM_113_WIDTH/8-1:0] ap_bram_oarg_113_we0,
    input ap_bram_oarg_113_en0,
    input [M_AXIS_BRAM_113_ADDR_WIDTH-1:0] ap_bram_oarg_113_addr1,
    input [M_AXIS_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_din1,
    output [M_AXIS_BRAM_113_WIDTH-1:0] ap_bram_oarg_113_dout1,
    input ap_bram_oarg_113_clk1,
    input ap_bram_oarg_113_rst1,
    input [M_AXIS_BRAM_113_WIDTH/8-1:0] ap_bram_oarg_113_we1,
    input ap_bram_oarg_113_en1,
    //out BRAM to AXI-Stream interface 114
    input m_axis_bram_114_aclk,
    input m_axis_bram_114_aresetn,
    output m_axis_bram_114_tlast,
    output m_axis_bram_114_tvalid,
    output [M_AXIS_BRAM_114_DMWIDTH/8-1:0] m_axis_bram_114_tkeep,
    output [M_AXIS_BRAM_114_DMWIDTH/8-1:0] m_axis_bram_114_tstrb,
    output [M_AXIS_BRAM_114_DMWIDTH-1:0] m_axis_bram_114_tdata,
    input m_axis_bram_114_tready,
    input [M_AXIS_BRAM_114_ADDR_WIDTH-1:0] ap_bram_oarg_114_addr0,
    input [M_AXIS_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_din0,
    output [M_AXIS_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_dout0,
    input ap_bram_oarg_114_clk0,
    input ap_bram_oarg_114_rst0,
    input [M_AXIS_BRAM_114_WIDTH/8-1:0] ap_bram_oarg_114_we0,
    input ap_bram_oarg_114_en0,
    input [M_AXIS_BRAM_114_ADDR_WIDTH-1:0] ap_bram_oarg_114_addr1,
    input [M_AXIS_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_din1,
    output [M_AXIS_BRAM_114_WIDTH-1:0] ap_bram_oarg_114_dout1,
    input ap_bram_oarg_114_clk1,
    input ap_bram_oarg_114_rst1,
    input [M_AXIS_BRAM_114_WIDTH/8-1:0] ap_bram_oarg_114_we1,
    input ap_bram_oarg_114_en1,
    //out BRAM to AXI-Stream interface 115
    input m_axis_bram_115_aclk,
    input m_axis_bram_115_aresetn,
    output m_axis_bram_115_tlast,
    output m_axis_bram_115_tvalid,
    output [M_AXIS_BRAM_115_DMWIDTH/8-1:0] m_axis_bram_115_tkeep,
    output [M_AXIS_BRAM_115_DMWIDTH/8-1:0] m_axis_bram_115_tstrb,
    output [M_AXIS_BRAM_115_DMWIDTH-1:0] m_axis_bram_115_tdata,
    input m_axis_bram_115_tready,
    input [M_AXIS_BRAM_115_ADDR_WIDTH-1:0] ap_bram_oarg_115_addr0,
    input [M_AXIS_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_din0,
    output [M_AXIS_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_dout0,
    input ap_bram_oarg_115_clk0,
    input ap_bram_oarg_115_rst0,
    input [M_AXIS_BRAM_115_WIDTH/8-1:0] ap_bram_oarg_115_we0,
    input ap_bram_oarg_115_en0,
    input [M_AXIS_BRAM_115_ADDR_WIDTH-1:0] ap_bram_oarg_115_addr1,
    input [M_AXIS_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_din1,
    output [M_AXIS_BRAM_115_WIDTH-1:0] ap_bram_oarg_115_dout1,
    input ap_bram_oarg_115_clk1,
    input ap_bram_oarg_115_rst1,
    input [M_AXIS_BRAM_115_WIDTH/8-1:0] ap_bram_oarg_115_we1,
    input ap_bram_oarg_115_en1,
    //out BRAM to AXI-Stream interface 116
    input m_axis_bram_116_aclk,
    input m_axis_bram_116_aresetn,
    output m_axis_bram_116_tlast,
    output m_axis_bram_116_tvalid,
    output [M_AXIS_BRAM_116_DMWIDTH/8-1:0] m_axis_bram_116_tkeep,
    output [M_AXIS_BRAM_116_DMWIDTH/8-1:0] m_axis_bram_116_tstrb,
    output [M_AXIS_BRAM_116_DMWIDTH-1:0] m_axis_bram_116_tdata,
    input m_axis_bram_116_tready,
    input [M_AXIS_BRAM_116_ADDR_WIDTH-1:0] ap_bram_oarg_116_addr0,
    input [M_AXIS_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_din0,
    output [M_AXIS_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_dout0,
    input ap_bram_oarg_116_clk0,
    input ap_bram_oarg_116_rst0,
    input [M_AXIS_BRAM_116_WIDTH/8-1:0] ap_bram_oarg_116_we0,
    input ap_bram_oarg_116_en0,
    input [M_AXIS_BRAM_116_ADDR_WIDTH-1:0] ap_bram_oarg_116_addr1,
    input [M_AXIS_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_din1,
    output [M_AXIS_BRAM_116_WIDTH-1:0] ap_bram_oarg_116_dout1,
    input ap_bram_oarg_116_clk1,
    input ap_bram_oarg_116_rst1,
    input [M_AXIS_BRAM_116_WIDTH/8-1:0] ap_bram_oarg_116_we1,
    input ap_bram_oarg_116_en1,
    //out BRAM to AXI-Stream interface 117
    input m_axis_bram_117_aclk,
    input m_axis_bram_117_aresetn,
    output m_axis_bram_117_tlast,
    output m_axis_bram_117_tvalid,
    output [M_AXIS_BRAM_117_DMWIDTH/8-1:0] m_axis_bram_117_tkeep,
    output [M_AXIS_BRAM_117_DMWIDTH/8-1:0] m_axis_bram_117_tstrb,
    output [M_AXIS_BRAM_117_DMWIDTH-1:0] m_axis_bram_117_tdata,
    input m_axis_bram_117_tready,
    input [M_AXIS_BRAM_117_ADDR_WIDTH-1:0] ap_bram_oarg_117_addr0,
    input [M_AXIS_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_din0,
    output [M_AXIS_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_dout0,
    input ap_bram_oarg_117_clk0,
    input ap_bram_oarg_117_rst0,
    input [M_AXIS_BRAM_117_WIDTH/8-1:0] ap_bram_oarg_117_we0,
    input ap_bram_oarg_117_en0,
    input [M_AXIS_BRAM_117_ADDR_WIDTH-1:0] ap_bram_oarg_117_addr1,
    input [M_AXIS_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_din1,
    output [M_AXIS_BRAM_117_WIDTH-1:0] ap_bram_oarg_117_dout1,
    input ap_bram_oarg_117_clk1,
    input ap_bram_oarg_117_rst1,
    input [M_AXIS_BRAM_117_WIDTH/8-1:0] ap_bram_oarg_117_we1,
    input ap_bram_oarg_117_en1,
    //out BRAM to AXI-Stream interface 118
    input m_axis_bram_118_aclk,
    input m_axis_bram_118_aresetn,
    output m_axis_bram_118_tlast,
    output m_axis_bram_118_tvalid,
    output [M_AXIS_BRAM_118_DMWIDTH/8-1:0] m_axis_bram_118_tkeep,
    output [M_AXIS_BRAM_118_DMWIDTH/8-1:0] m_axis_bram_118_tstrb,
    output [M_AXIS_BRAM_118_DMWIDTH-1:0] m_axis_bram_118_tdata,
    input m_axis_bram_118_tready,
    input [M_AXIS_BRAM_118_ADDR_WIDTH-1:0] ap_bram_oarg_118_addr0,
    input [M_AXIS_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_din0,
    output [M_AXIS_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_dout0,
    input ap_bram_oarg_118_clk0,
    input ap_bram_oarg_118_rst0,
    input [M_AXIS_BRAM_118_WIDTH/8-1:0] ap_bram_oarg_118_we0,
    input ap_bram_oarg_118_en0,
    input [M_AXIS_BRAM_118_ADDR_WIDTH-1:0] ap_bram_oarg_118_addr1,
    input [M_AXIS_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_din1,
    output [M_AXIS_BRAM_118_WIDTH-1:0] ap_bram_oarg_118_dout1,
    input ap_bram_oarg_118_clk1,
    input ap_bram_oarg_118_rst1,
    input [M_AXIS_BRAM_118_WIDTH/8-1:0] ap_bram_oarg_118_we1,
    input ap_bram_oarg_118_en1,
    //out BRAM to AXI-Stream interface 119
    input m_axis_bram_119_aclk,
    input m_axis_bram_119_aresetn,
    output m_axis_bram_119_tlast,
    output m_axis_bram_119_tvalid,
    output [M_AXIS_BRAM_119_DMWIDTH/8-1:0] m_axis_bram_119_tkeep,
    output [M_AXIS_BRAM_119_DMWIDTH/8-1:0] m_axis_bram_119_tstrb,
    output [M_AXIS_BRAM_119_DMWIDTH-1:0] m_axis_bram_119_tdata,
    input m_axis_bram_119_tready,
    input [M_AXIS_BRAM_119_ADDR_WIDTH-1:0] ap_bram_oarg_119_addr0,
    input [M_AXIS_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_din0,
    output [M_AXIS_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_dout0,
    input ap_bram_oarg_119_clk0,
    input ap_bram_oarg_119_rst0,
    input [M_AXIS_BRAM_119_WIDTH/8-1:0] ap_bram_oarg_119_we0,
    input ap_bram_oarg_119_en0,
    input [M_AXIS_BRAM_119_ADDR_WIDTH-1:0] ap_bram_oarg_119_addr1,
    input [M_AXIS_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_din1,
    output [M_AXIS_BRAM_119_WIDTH-1:0] ap_bram_oarg_119_dout1,
    input ap_bram_oarg_119_clk1,
    input ap_bram_oarg_119_rst1,
    input [M_AXIS_BRAM_119_WIDTH/8-1:0] ap_bram_oarg_119_we1,
    input ap_bram_oarg_119_en1,
    //out BRAM to AXI-Stream interface 120
    input m_axis_bram_120_aclk,
    input m_axis_bram_120_aresetn,
    output m_axis_bram_120_tlast,
    output m_axis_bram_120_tvalid,
    output [M_AXIS_BRAM_120_DMWIDTH/8-1:0] m_axis_bram_120_tkeep,
    output [M_AXIS_BRAM_120_DMWIDTH/8-1:0] m_axis_bram_120_tstrb,
    output [M_AXIS_BRAM_120_DMWIDTH-1:0] m_axis_bram_120_tdata,
    input m_axis_bram_120_tready,
    input [M_AXIS_BRAM_120_ADDR_WIDTH-1:0] ap_bram_oarg_120_addr0,
    input [M_AXIS_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_din0,
    output [M_AXIS_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_dout0,
    input ap_bram_oarg_120_clk0,
    input ap_bram_oarg_120_rst0,
    input [M_AXIS_BRAM_120_WIDTH/8-1:0] ap_bram_oarg_120_we0,
    input ap_bram_oarg_120_en0,
    input [M_AXIS_BRAM_120_ADDR_WIDTH-1:0] ap_bram_oarg_120_addr1,
    input [M_AXIS_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_din1,
    output [M_AXIS_BRAM_120_WIDTH-1:0] ap_bram_oarg_120_dout1,
    input ap_bram_oarg_120_clk1,
    input ap_bram_oarg_120_rst1,
    input [M_AXIS_BRAM_120_WIDTH/8-1:0] ap_bram_oarg_120_we1,
    input ap_bram_oarg_120_en1,
    //out BRAM to AXI-Stream interface 121
    input m_axis_bram_121_aclk,
    input m_axis_bram_121_aresetn,
    output m_axis_bram_121_tlast,
    output m_axis_bram_121_tvalid,
    output [M_AXIS_BRAM_121_DMWIDTH/8-1:0] m_axis_bram_121_tkeep,
    output [M_AXIS_BRAM_121_DMWIDTH/8-1:0] m_axis_bram_121_tstrb,
    output [M_AXIS_BRAM_121_DMWIDTH-1:0] m_axis_bram_121_tdata,
    input m_axis_bram_121_tready,
    input [M_AXIS_BRAM_121_ADDR_WIDTH-1:0] ap_bram_oarg_121_addr0,
    input [M_AXIS_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_din0,
    output [M_AXIS_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_dout0,
    input ap_bram_oarg_121_clk0,
    input ap_bram_oarg_121_rst0,
    input [M_AXIS_BRAM_121_WIDTH/8-1:0] ap_bram_oarg_121_we0,
    input ap_bram_oarg_121_en0,
    input [M_AXIS_BRAM_121_ADDR_WIDTH-1:0] ap_bram_oarg_121_addr1,
    input [M_AXIS_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_din1,
    output [M_AXIS_BRAM_121_WIDTH-1:0] ap_bram_oarg_121_dout1,
    input ap_bram_oarg_121_clk1,
    input ap_bram_oarg_121_rst1,
    input [M_AXIS_BRAM_121_WIDTH/8-1:0] ap_bram_oarg_121_we1,
    input ap_bram_oarg_121_en1,
    //out BRAM to AXI-Stream interface 122
    input m_axis_bram_122_aclk,
    input m_axis_bram_122_aresetn,
    output m_axis_bram_122_tlast,
    output m_axis_bram_122_tvalid,
    output [M_AXIS_BRAM_122_DMWIDTH/8-1:0] m_axis_bram_122_tkeep,
    output [M_AXIS_BRAM_122_DMWIDTH/8-1:0] m_axis_bram_122_tstrb,
    output [M_AXIS_BRAM_122_DMWIDTH-1:0] m_axis_bram_122_tdata,
    input m_axis_bram_122_tready,
    input [M_AXIS_BRAM_122_ADDR_WIDTH-1:0] ap_bram_oarg_122_addr0,
    input [M_AXIS_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_din0,
    output [M_AXIS_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_dout0,
    input ap_bram_oarg_122_clk0,
    input ap_bram_oarg_122_rst0,
    input [M_AXIS_BRAM_122_WIDTH/8-1:0] ap_bram_oarg_122_we0,
    input ap_bram_oarg_122_en0,
    input [M_AXIS_BRAM_122_ADDR_WIDTH-1:0] ap_bram_oarg_122_addr1,
    input [M_AXIS_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_din1,
    output [M_AXIS_BRAM_122_WIDTH-1:0] ap_bram_oarg_122_dout1,
    input ap_bram_oarg_122_clk1,
    input ap_bram_oarg_122_rst1,
    input [M_AXIS_BRAM_122_WIDTH/8-1:0] ap_bram_oarg_122_we1,
    input ap_bram_oarg_122_en1,
    //out BRAM to AXI-Stream interface 123
    input m_axis_bram_123_aclk,
    input m_axis_bram_123_aresetn,
    output m_axis_bram_123_tlast,
    output m_axis_bram_123_tvalid,
    output [M_AXIS_BRAM_123_DMWIDTH/8-1:0] m_axis_bram_123_tkeep,
    output [M_AXIS_BRAM_123_DMWIDTH/8-1:0] m_axis_bram_123_tstrb,
    output [M_AXIS_BRAM_123_DMWIDTH-1:0] m_axis_bram_123_tdata,
    input m_axis_bram_123_tready,
    input [M_AXIS_BRAM_123_ADDR_WIDTH-1:0] ap_bram_oarg_123_addr0,
    input [M_AXIS_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_din0,
    output [M_AXIS_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_dout0,
    input ap_bram_oarg_123_clk0,
    input ap_bram_oarg_123_rst0,
    input [M_AXIS_BRAM_123_WIDTH/8-1:0] ap_bram_oarg_123_we0,
    input ap_bram_oarg_123_en0,
    input [M_AXIS_BRAM_123_ADDR_WIDTH-1:0] ap_bram_oarg_123_addr1,
    input [M_AXIS_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_din1,
    output [M_AXIS_BRAM_123_WIDTH-1:0] ap_bram_oarg_123_dout1,
    input ap_bram_oarg_123_clk1,
    input ap_bram_oarg_123_rst1,
    input [M_AXIS_BRAM_123_WIDTH/8-1:0] ap_bram_oarg_123_we1,
    input ap_bram_oarg_123_en1,
    //out BRAM to AXI-Stream interface 124
    input m_axis_bram_124_aclk,
    input m_axis_bram_124_aresetn,
    output m_axis_bram_124_tlast,
    output m_axis_bram_124_tvalid,
    output [M_AXIS_BRAM_124_DMWIDTH/8-1:0] m_axis_bram_124_tkeep,
    output [M_AXIS_BRAM_124_DMWIDTH/8-1:0] m_axis_bram_124_tstrb,
    output [M_AXIS_BRAM_124_DMWIDTH-1:0] m_axis_bram_124_tdata,
    input m_axis_bram_124_tready,
    input [M_AXIS_BRAM_124_ADDR_WIDTH-1:0] ap_bram_oarg_124_addr0,
    input [M_AXIS_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_din0,
    output [M_AXIS_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_dout0,
    input ap_bram_oarg_124_clk0,
    input ap_bram_oarg_124_rst0,
    input [M_AXIS_BRAM_124_WIDTH/8-1:0] ap_bram_oarg_124_we0,
    input ap_bram_oarg_124_en0,
    input [M_AXIS_BRAM_124_ADDR_WIDTH-1:0] ap_bram_oarg_124_addr1,
    input [M_AXIS_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_din1,
    output [M_AXIS_BRAM_124_WIDTH-1:0] ap_bram_oarg_124_dout1,
    input ap_bram_oarg_124_clk1,
    input ap_bram_oarg_124_rst1,
    input [M_AXIS_BRAM_124_WIDTH/8-1:0] ap_bram_oarg_124_we1,
    input ap_bram_oarg_124_en1,
    //out BRAM to AXI-Stream interface 125
    input m_axis_bram_125_aclk,
    input m_axis_bram_125_aresetn,
    output m_axis_bram_125_tlast,
    output m_axis_bram_125_tvalid,
    output [M_AXIS_BRAM_125_DMWIDTH/8-1:0] m_axis_bram_125_tkeep,
    output [M_AXIS_BRAM_125_DMWIDTH/8-1:0] m_axis_bram_125_tstrb,
    output [M_AXIS_BRAM_125_DMWIDTH-1:0] m_axis_bram_125_tdata,
    input m_axis_bram_125_tready,
    input [M_AXIS_BRAM_125_ADDR_WIDTH-1:0] ap_bram_oarg_125_addr0,
    input [M_AXIS_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_din0,
    output [M_AXIS_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_dout0,
    input ap_bram_oarg_125_clk0,
    input ap_bram_oarg_125_rst0,
    input [M_AXIS_BRAM_125_WIDTH/8-1:0] ap_bram_oarg_125_we0,
    input ap_bram_oarg_125_en0,
    input [M_AXIS_BRAM_125_ADDR_WIDTH-1:0] ap_bram_oarg_125_addr1,
    input [M_AXIS_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_din1,
    output [M_AXIS_BRAM_125_WIDTH-1:0] ap_bram_oarg_125_dout1,
    input ap_bram_oarg_125_clk1,
    input ap_bram_oarg_125_rst1,
    input [M_AXIS_BRAM_125_WIDTH/8-1:0] ap_bram_oarg_125_we1,
    input ap_bram_oarg_125_en1,
    //out BRAM to AXI-Stream interface 126
    input m_axis_bram_126_aclk,
    input m_axis_bram_126_aresetn,
    output m_axis_bram_126_tlast,
    output m_axis_bram_126_tvalid,
    output [M_AXIS_BRAM_126_DMWIDTH/8-1:0] m_axis_bram_126_tkeep,
    output [M_AXIS_BRAM_126_DMWIDTH/8-1:0] m_axis_bram_126_tstrb,
    output [M_AXIS_BRAM_126_DMWIDTH-1:0] m_axis_bram_126_tdata,
    input m_axis_bram_126_tready,
    input [M_AXIS_BRAM_126_ADDR_WIDTH-1:0] ap_bram_oarg_126_addr0,
    input [M_AXIS_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_din0,
    output [M_AXIS_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_dout0,
    input ap_bram_oarg_126_clk0,
    input ap_bram_oarg_126_rst0,
    input [M_AXIS_BRAM_126_WIDTH/8-1:0] ap_bram_oarg_126_we0,
    input ap_bram_oarg_126_en0,
    input [M_AXIS_BRAM_126_ADDR_WIDTH-1:0] ap_bram_oarg_126_addr1,
    input [M_AXIS_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_din1,
    output [M_AXIS_BRAM_126_WIDTH-1:0] ap_bram_oarg_126_dout1,
    input ap_bram_oarg_126_clk1,
    input ap_bram_oarg_126_rst1,
    input [M_AXIS_BRAM_126_WIDTH/8-1:0] ap_bram_oarg_126_we1,
    input ap_bram_oarg_126_en1,
    //out BRAM to AXI-Stream interface 127
    input m_axis_bram_127_aclk,
    input m_axis_bram_127_aresetn,
    output m_axis_bram_127_tlast,
    output m_axis_bram_127_tvalid,
    output [M_AXIS_BRAM_127_DMWIDTH/8-1:0] m_axis_bram_127_tkeep,
    output [M_AXIS_BRAM_127_DMWIDTH/8-1:0] m_axis_bram_127_tstrb,
    output [M_AXIS_BRAM_127_DMWIDTH-1:0] m_axis_bram_127_tdata,
    input m_axis_bram_127_tready,
    input [M_AXIS_BRAM_127_ADDR_WIDTH-1:0] ap_bram_oarg_127_addr0,
    input [M_AXIS_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_din0,
    output [M_AXIS_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_dout0,
    input ap_bram_oarg_127_clk0,
    input ap_bram_oarg_127_rst0,
    input [M_AXIS_BRAM_127_WIDTH/8-1:0] ap_bram_oarg_127_we0,
    input ap_bram_oarg_127_en0,
    input [M_AXIS_BRAM_127_ADDR_WIDTH-1:0] ap_bram_oarg_127_addr1,
    input [M_AXIS_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_din1,
    output [M_AXIS_BRAM_127_WIDTH-1:0] ap_bram_oarg_127_dout1,
    input ap_bram_oarg_127_clk1,
    input ap_bram_oarg_127_rst1,
    input [M_AXIS_BRAM_127_WIDTH/8-1:0] ap_bram_oarg_127_we1,
    input ap_bram_oarg_127_en1,
    //-----------------------------------------------------
    //input AXI-Stream pass-through interface 0
    input s_axis_iarg_0_aclk,
    input s_axis_iarg_0_aresetn,
    input s_axis_iarg_0_tlast,
    input s_axis_iarg_0_tvalid,
    input [S_AXIS_IARG_0_DMWIDTH/8-1:0] s_axis_iarg_0_tkeep,
    input [S_AXIS_IARG_0_DMWIDTH/8-1:0] s_axis_iarg_0_tstrb,
    input [S_AXIS_IARG_0_DMWIDTH-1:0] s_axis_iarg_0_tdata,
    output s_axis_iarg_0_tready,
    input ap_axis_iarg_0_tready,
    output ap_axis_iarg_0_tlast,
    output ap_axis_iarg_0_tvalid,
    output [S_AXIS_IARG_0_WIDTH/8-1:0] ap_axis_iarg_0_tkeep,
    output [S_AXIS_IARG_0_WIDTH/8-1:0] ap_axis_iarg_0_tstrb,
    output [S_AXIS_IARG_0_WIDTH-1:0] ap_axis_iarg_0_tdata,
    //input AXI-Stream pass-through interface 1
    input s_axis_iarg_1_aclk,
    input s_axis_iarg_1_aresetn,
    input s_axis_iarg_1_tlast,
    input s_axis_iarg_1_tvalid,
    input [S_AXIS_IARG_1_DMWIDTH/8-1:0] s_axis_iarg_1_tkeep,
    input [S_AXIS_IARG_1_DMWIDTH/8-1:0] s_axis_iarg_1_tstrb,
    input [S_AXIS_IARG_1_DMWIDTH-1:0] s_axis_iarg_1_tdata,
    output s_axis_iarg_1_tready,
    input ap_axis_iarg_1_tready,
    output ap_axis_iarg_1_tlast,
    output ap_axis_iarg_1_tvalid,
    output [S_AXIS_IARG_1_WIDTH/8-1:0] ap_axis_iarg_1_tkeep,
    output [S_AXIS_IARG_1_WIDTH/8-1:0] ap_axis_iarg_1_tstrb,
    output [S_AXIS_IARG_1_WIDTH-1:0] ap_axis_iarg_1_tdata,
    //input AXI-Stream pass-through interface 2
    input s_axis_iarg_2_aclk,
    input s_axis_iarg_2_aresetn,
    input s_axis_iarg_2_tlast,
    input s_axis_iarg_2_tvalid,
    input [S_AXIS_IARG_2_DMWIDTH/8-1:0] s_axis_iarg_2_tkeep,
    input [S_AXIS_IARG_2_DMWIDTH/8-1:0] s_axis_iarg_2_tstrb,
    input [S_AXIS_IARG_2_DMWIDTH-1:0] s_axis_iarg_2_tdata,
    output s_axis_iarg_2_tready,
    input ap_axis_iarg_2_tready,
    output ap_axis_iarg_2_tlast,
    output ap_axis_iarg_2_tvalid,
    output [S_AXIS_IARG_2_WIDTH/8-1:0] ap_axis_iarg_2_tkeep,
    output [S_AXIS_IARG_2_WIDTH/8-1:0] ap_axis_iarg_2_tstrb,
    output [S_AXIS_IARG_2_WIDTH-1:0] ap_axis_iarg_2_tdata,
    //input AXI-Stream pass-through interface 3
    input s_axis_iarg_3_aclk,
    input s_axis_iarg_3_aresetn,
    input s_axis_iarg_3_tlast,
    input s_axis_iarg_3_tvalid,
    input [S_AXIS_IARG_3_DMWIDTH/8-1:0] s_axis_iarg_3_tkeep,
    input [S_AXIS_IARG_3_DMWIDTH/8-1:0] s_axis_iarg_3_tstrb,
    input [S_AXIS_IARG_3_DMWIDTH-1:0] s_axis_iarg_3_tdata,
    output s_axis_iarg_3_tready,
    input ap_axis_iarg_3_tready,
    output ap_axis_iarg_3_tlast,
    output ap_axis_iarg_3_tvalid,
    output [S_AXIS_IARG_3_WIDTH/8-1:0] ap_axis_iarg_3_tkeep,
    output [S_AXIS_IARG_3_WIDTH/8-1:0] ap_axis_iarg_3_tstrb,
    output [S_AXIS_IARG_3_WIDTH-1:0] ap_axis_iarg_3_tdata,
    //input AXI-Stream pass-through interface 4
    input s_axis_iarg_4_aclk,
    input s_axis_iarg_4_aresetn,
    input s_axis_iarg_4_tlast,
    input s_axis_iarg_4_tvalid,
    input [S_AXIS_IARG_4_DMWIDTH/8-1:0] s_axis_iarg_4_tkeep,
    input [S_AXIS_IARG_4_DMWIDTH/8-1:0] s_axis_iarg_4_tstrb,
    input [S_AXIS_IARG_4_DMWIDTH-1:0] s_axis_iarg_4_tdata,
    output s_axis_iarg_4_tready,
    input ap_axis_iarg_4_tready,
    output ap_axis_iarg_4_tlast,
    output ap_axis_iarg_4_tvalid,
    output [S_AXIS_IARG_4_WIDTH/8-1:0] ap_axis_iarg_4_tkeep,
    output [S_AXIS_IARG_4_WIDTH/8-1:0] ap_axis_iarg_4_tstrb,
    output [S_AXIS_IARG_4_WIDTH-1:0] ap_axis_iarg_4_tdata,
    //input AXI-Stream pass-through interface 5
    input s_axis_iarg_5_aclk,
    input s_axis_iarg_5_aresetn,
    input s_axis_iarg_5_tlast,
    input s_axis_iarg_5_tvalid,
    input [S_AXIS_IARG_5_DMWIDTH/8-1:0] s_axis_iarg_5_tkeep,
    input [S_AXIS_IARG_5_DMWIDTH/8-1:0] s_axis_iarg_5_tstrb,
    input [S_AXIS_IARG_5_DMWIDTH-1:0] s_axis_iarg_5_tdata,
    output s_axis_iarg_5_tready,
    input ap_axis_iarg_5_tready,
    output ap_axis_iarg_5_tlast,
    output ap_axis_iarg_5_tvalid,
    output [S_AXIS_IARG_5_WIDTH/8-1:0] ap_axis_iarg_5_tkeep,
    output [S_AXIS_IARG_5_WIDTH/8-1:0] ap_axis_iarg_5_tstrb,
    output [S_AXIS_IARG_5_WIDTH-1:0] ap_axis_iarg_5_tdata,
    //input AXI-Stream pass-through interface 6
    input s_axis_iarg_6_aclk,
    input s_axis_iarg_6_aresetn,
    input s_axis_iarg_6_tlast,
    input s_axis_iarg_6_tvalid,
    input [S_AXIS_IARG_6_DMWIDTH/8-1:0] s_axis_iarg_6_tkeep,
    input [S_AXIS_IARG_6_DMWIDTH/8-1:0] s_axis_iarg_6_tstrb,
    input [S_AXIS_IARG_6_DMWIDTH-1:0] s_axis_iarg_6_tdata,
    output s_axis_iarg_6_tready,
    input ap_axis_iarg_6_tready,
    output ap_axis_iarg_6_tlast,
    output ap_axis_iarg_6_tvalid,
    output [S_AXIS_IARG_6_WIDTH/8-1:0] ap_axis_iarg_6_tkeep,
    output [S_AXIS_IARG_6_WIDTH/8-1:0] ap_axis_iarg_6_tstrb,
    output [S_AXIS_IARG_6_WIDTH-1:0] ap_axis_iarg_6_tdata,
    //input AXI-Stream pass-through interface 7
    input s_axis_iarg_7_aclk,
    input s_axis_iarg_7_aresetn,
    input s_axis_iarg_7_tlast,
    input s_axis_iarg_7_tvalid,
    input [S_AXIS_IARG_7_DMWIDTH/8-1:0] s_axis_iarg_7_tkeep,
    input [S_AXIS_IARG_7_DMWIDTH/8-1:0] s_axis_iarg_7_tstrb,
    input [S_AXIS_IARG_7_DMWIDTH-1:0] s_axis_iarg_7_tdata,
    output s_axis_iarg_7_tready,
    input ap_axis_iarg_7_tready,
    output ap_axis_iarg_7_tlast,
    output ap_axis_iarg_7_tvalid,
    output [S_AXIS_IARG_7_WIDTH/8-1:0] ap_axis_iarg_7_tkeep,
    output [S_AXIS_IARG_7_WIDTH/8-1:0] ap_axis_iarg_7_tstrb,
    output [S_AXIS_IARG_7_WIDTH-1:0] ap_axis_iarg_7_tdata,
    //input AXI-Stream pass-through interface 8
    input s_axis_iarg_8_aclk,
    input s_axis_iarg_8_aresetn,
    input s_axis_iarg_8_tlast,
    input s_axis_iarg_8_tvalid,
    input [S_AXIS_IARG_8_DMWIDTH/8-1:0] s_axis_iarg_8_tkeep,
    input [S_AXIS_IARG_8_DMWIDTH/8-1:0] s_axis_iarg_8_tstrb,
    input [S_AXIS_IARG_8_DMWIDTH-1:0] s_axis_iarg_8_tdata,
    output s_axis_iarg_8_tready,
    input ap_axis_iarg_8_tready,
    output ap_axis_iarg_8_tlast,
    output ap_axis_iarg_8_tvalid,
    output [S_AXIS_IARG_8_WIDTH/8-1:0] ap_axis_iarg_8_tkeep,
    output [S_AXIS_IARG_8_WIDTH/8-1:0] ap_axis_iarg_8_tstrb,
    output [S_AXIS_IARG_8_WIDTH-1:0] ap_axis_iarg_8_tdata,
    //input AXI-Stream pass-through interface 9
    input s_axis_iarg_9_aclk,
    input s_axis_iarg_9_aresetn,
    input s_axis_iarg_9_tlast,
    input s_axis_iarg_9_tvalid,
    input [S_AXIS_IARG_9_DMWIDTH/8-1:0] s_axis_iarg_9_tkeep,
    input [S_AXIS_IARG_9_DMWIDTH/8-1:0] s_axis_iarg_9_tstrb,
    input [S_AXIS_IARG_9_DMWIDTH-1:0] s_axis_iarg_9_tdata,
    output s_axis_iarg_9_tready,
    input ap_axis_iarg_9_tready,
    output ap_axis_iarg_9_tlast,
    output ap_axis_iarg_9_tvalid,
    output [S_AXIS_IARG_9_WIDTH/8-1:0] ap_axis_iarg_9_tkeep,
    output [S_AXIS_IARG_9_WIDTH/8-1:0] ap_axis_iarg_9_tstrb,
    output [S_AXIS_IARG_9_WIDTH-1:0] ap_axis_iarg_9_tdata,
    //input AXI-Stream pass-through interface 10
    input s_axis_iarg_10_aclk,
    input s_axis_iarg_10_aresetn,
    input s_axis_iarg_10_tlast,
    input s_axis_iarg_10_tvalid,
    input [S_AXIS_IARG_10_DMWIDTH/8-1:0] s_axis_iarg_10_tkeep,
    input [S_AXIS_IARG_10_DMWIDTH/8-1:0] s_axis_iarg_10_tstrb,
    input [S_AXIS_IARG_10_DMWIDTH-1:0] s_axis_iarg_10_tdata,
    output s_axis_iarg_10_tready,
    input ap_axis_iarg_10_tready,
    output ap_axis_iarg_10_tlast,
    output ap_axis_iarg_10_tvalid,
    output [S_AXIS_IARG_10_WIDTH/8-1:0] ap_axis_iarg_10_tkeep,
    output [S_AXIS_IARG_10_WIDTH/8-1:0] ap_axis_iarg_10_tstrb,
    output [S_AXIS_IARG_10_WIDTH-1:0] ap_axis_iarg_10_tdata,
    //input AXI-Stream pass-through interface 11
    input s_axis_iarg_11_aclk,
    input s_axis_iarg_11_aresetn,
    input s_axis_iarg_11_tlast,
    input s_axis_iarg_11_tvalid,
    input [S_AXIS_IARG_11_DMWIDTH/8-1:0] s_axis_iarg_11_tkeep,
    input [S_AXIS_IARG_11_DMWIDTH/8-1:0] s_axis_iarg_11_tstrb,
    input [S_AXIS_IARG_11_DMWIDTH-1:0] s_axis_iarg_11_tdata,
    output s_axis_iarg_11_tready,
    input ap_axis_iarg_11_tready,
    output ap_axis_iarg_11_tlast,
    output ap_axis_iarg_11_tvalid,
    output [S_AXIS_IARG_11_WIDTH/8-1:0] ap_axis_iarg_11_tkeep,
    output [S_AXIS_IARG_11_WIDTH/8-1:0] ap_axis_iarg_11_tstrb,
    output [S_AXIS_IARG_11_WIDTH-1:0] ap_axis_iarg_11_tdata,
    //input AXI-Stream pass-through interface 12
    input s_axis_iarg_12_aclk,
    input s_axis_iarg_12_aresetn,
    input s_axis_iarg_12_tlast,
    input s_axis_iarg_12_tvalid,
    input [S_AXIS_IARG_12_DMWIDTH/8-1:0] s_axis_iarg_12_tkeep,
    input [S_AXIS_IARG_12_DMWIDTH/8-1:0] s_axis_iarg_12_tstrb,
    input [S_AXIS_IARG_12_DMWIDTH-1:0] s_axis_iarg_12_tdata,
    output s_axis_iarg_12_tready,
    input ap_axis_iarg_12_tready,
    output ap_axis_iarg_12_tlast,
    output ap_axis_iarg_12_tvalid,
    output [S_AXIS_IARG_12_WIDTH/8-1:0] ap_axis_iarg_12_tkeep,
    output [S_AXIS_IARG_12_WIDTH/8-1:0] ap_axis_iarg_12_tstrb,
    output [S_AXIS_IARG_12_WIDTH-1:0] ap_axis_iarg_12_tdata,
    //input AXI-Stream pass-through interface 13
    input s_axis_iarg_13_aclk,
    input s_axis_iarg_13_aresetn,
    input s_axis_iarg_13_tlast,
    input s_axis_iarg_13_tvalid,
    input [S_AXIS_IARG_13_DMWIDTH/8-1:0] s_axis_iarg_13_tkeep,
    input [S_AXIS_IARG_13_DMWIDTH/8-1:0] s_axis_iarg_13_tstrb,
    input [S_AXIS_IARG_13_DMWIDTH-1:0] s_axis_iarg_13_tdata,
    output s_axis_iarg_13_tready,
    input ap_axis_iarg_13_tready,
    output ap_axis_iarg_13_tlast,
    output ap_axis_iarg_13_tvalid,
    output [S_AXIS_IARG_13_WIDTH/8-1:0] ap_axis_iarg_13_tkeep,
    output [S_AXIS_IARG_13_WIDTH/8-1:0] ap_axis_iarg_13_tstrb,
    output [S_AXIS_IARG_13_WIDTH-1:0] ap_axis_iarg_13_tdata,
    //input AXI-Stream pass-through interface 14
    input s_axis_iarg_14_aclk,
    input s_axis_iarg_14_aresetn,
    input s_axis_iarg_14_tlast,
    input s_axis_iarg_14_tvalid,
    input [S_AXIS_IARG_14_DMWIDTH/8-1:0] s_axis_iarg_14_tkeep,
    input [S_AXIS_IARG_14_DMWIDTH/8-1:0] s_axis_iarg_14_tstrb,
    input [S_AXIS_IARG_14_DMWIDTH-1:0] s_axis_iarg_14_tdata,
    output s_axis_iarg_14_tready,
    input ap_axis_iarg_14_tready,
    output ap_axis_iarg_14_tlast,
    output ap_axis_iarg_14_tvalid,
    output [S_AXIS_IARG_14_WIDTH/8-1:0] ap_axis_iarg_14_tkeep,
    output [S_AXIS_IARG_14_WIDTH/8-1:0] ap_axis_iarg_14_tstrb,
    output [S_AXIS_IARG_14_WIDTH-1:0] ap_axis_iarg_14_tdata,
    //input AXI-Stream pass-through interface 15
    input s_axis_iarg_15_aclk,
    input s_axis_iarg_15_aresetn,
    input s_axis_iarg_15_tlast,
    input s_axis_iarg_15_tvalid,
    input [S_AXIS_IARG_15_DMWIDTH/8-1:0] s_axis_iarg_15_tkeep,
    input [S_AXIS_IARG_15_DMWIDTH/8-1:0] s_axis_iarg_15_tstrb,
    input [S_AXIS_IARG_15_DMWIDTH-1:0] s_axis_iarg_15_tdata,
    output s_axis_iarg_15_tready,
    input ap_axis_iarg_15_tready,
    output ap_axis_iarg_15_tlast,
    output ap_axis_iarg_15_tvalid,
    output [S_AXIS_IARG_15_WIDTH/8-1:0] ap_axis_iarg_15_tkeep,
    output [S_AXIS_IARG_15_WIDTH/8-1:0] ap_axis_iarg_15_tstrb,
    output [S_AXIS_IARG_15_WIDTH-1:0] ap_axis_iarg_15_tdata,
    //input AXI-Stream pass-through interface 16
    input s_axis_iarg_16_aclk,
    input s_axis_iarg_16_aresetn,
    input s_axis_iarg_16_tlast,
    input s_axis_iarg_16_tvalid,
    input [S_AXIS_IARG_16_DMWIDTH/8-1:0] s_axis_iarg_16_tkeep,
    input [S_AXIS_IARG_16_DMWIDTH/8-1:0] s_axis_iarg_16_tstrb,
    input [S_AXIS_IARG_16_DMWIDTH-1:0] s_axis_iarg_16_tdata,
    output s_axis_iarg_16_tready,
    input ap_axis_iarg_16_tready,
    output ap_axis_iarg_16_tlast,
    output ap_axis_iarg_16_tvalid,
    output [S_AXIS_IARG_16_WIDTH/8-1:0] ap_axis_iarg_16_tkeep,
    output [S_AXIS_IARG_16_WIDTH/8-1:0] ap_axis_iarg_16_tstrb,
    output [S_AXIS_IARG_16_WIDTH-1:0] ap_axis_iarg_16_tdata,
    //input AXI-Stream pass-through interface 17
    input s_axis_iarg_17_aclk,
    input s_axis_iarg_17_aresetn,
    input s_axis_iarg_17_tlast,
    input s_axis_iarg_17_tvalid,
    input [S_AXIS_IARG_17_DMWIDTH/8-1:0] s_axis_iarg_17_tkeep,
    input [S_AXIS_IARG_17_DMWIDTH/8-1:0] s_axis_iarg_17_tstrb,
    input [S_AXIS_IARG_17_DMWIDTH-1:0] s_axis_iarg_17_tdata,
    output s_axis_iarg_17_tready,
    input ap_axis_iarg_17_tready,
    output ap_axis_iarg_17_tlast,
    output ap_axis_iarg_17_tvalid,
    output [S_AXIS_IARG_17_WIDTH/8-1:0] ap_axis_iarg_17_tkeep,
    output [S_AXIS_IARG_17_WIDTH/8-1:0] ap_axis_iarg_17_tstrb,
    output [S_AXIS_IARG_17_WIDTH-1:0] ap_axis_iarg_17_tdata,
    //input AXI-Stream pass-through interface 18
    input s_axis_iarg_18_aclk,
    input s_axis_iarg_18_aresetn,
    input s_axis_iarg_18_tlast,
    input s_axis_iarg_18_tvalid,
    input [S_AXIS_IARG_18_DMWIDTH/8-1:0] s_axis_iarg_18_tkeep,
    input [S_AXIS_IARG_18_DMWIDTH/8-1:0] s_axis_iarg_18_tstrb,
    input [S_AXIS_IARG_18_DMWIDTH-1:0] s_axis_iarg_18_tdata,
    output s_axis_iarg_18_tready,
    input ap_axis_iarg_18_tready,
    output ap_axis_iarg_18_tlast,
    output ap_axis_iarg_18_tvalid,
    output [S_AXIS_IARG_18_WIDTH/8-1:0] ap_axis_iarg_18_tkeep,
    output [S_AXIS_IARG_18_WIDTH/8-1:0] ap_axis_iarg_18_tstrb,
    output [S_AXIS_IARG_18_WIDTH-1:0] ap_axis_iarg_18_tdata,
    //input AXI-Stream pass-through interface 19
    input s_axis_iarg_19_aclk,
    input s_axis_iarg_19_aresetn,
    input s_axis_iarg_19_tlast,
    input s_axis_iarg_19_tvalid,
    input [S_AXIS_IARG_19_DMWIDTH/8-1:0] s_axis_iarg_19_tkeep,
    input [S_AXIS_IARG_19_DMWIDTH/8-1:0] s_axis_iarg_19_tstrb,
    input [S_AXIS_IARG_19_DMWIDTH-1:0] s_axis_iarg_19_tdata,
    output s_axis_iarg_19_tready,
    input ap_axis_iarg_19_tready,
    output ap_axis_iarg_19_tlast,
    output ap_axis_iarg_19_tvalid,
    output [S_AXIS_IARG_19_WIDTH/8-1:0] ap_axis_iarg_19_tkeep,
    output [S_AXIS_IARG_19_WIDTH/8-1:0] ap_axis_iarg_19_tstrb,
    output [S_AXIS_IARG_19_WIDTH-1:0] ap_axis_iarg_19_tdata,
    //input AXI-Stream pass-through interface 20
    input s_axis_iarg_20_aclk,
    input s_axis_iarg_20_aresetn,
    input s_axis_iarg_20_tlast,
    input s_axis_iarg_20_tvalid,
    input [S_AXIS_IARG_20_DMWIDTH/8-1:0] s_axis_iarg_20_tkeep,
    input [S_AXIS_IARG_20_DMWIDTH/8-1:0] s_axis_iarg_20_tstrb,
    input [S_AXIS_IARG_20_DMWIDTH-1:0] s_axis_iarg_20_tdata,
    output s_axis_iarg_20_tready,
    input ap_axis_iarg_20_tready,
    output ap_axis_iarg_20_tlast,
    output ap_axis_iarg_20_tvalid,
    output [S_AXIS_IARG_20_WIDTH/8-1:0] ap_axis_iarg_20_tkeep,
    output [S_AXIS_IARG_20_WIDTH/8-1:0] ap_axis_iarg_20_tstrb,
    output [S_AXIS_IARG_20_WIDTH-1:0] ap_axis_iarg_20_tdata,
    //input AXI-Stream pass-through interface 21
    input s_axis_iarg_21_aclk,
    input s_axis_iarg_21_aresetn,
    input s_axis_iarg_21_tlast,
    input s_axis_iarg_21_tvalid,
    input [S_AXIS_IARG_21_DMWIDTH/8-1:0] s_axis_iarg_21_tkeep,
    input [S_AXIS_IARG_21_DMWIDTH/8-1:0] s_axis_iarg_21_tstrb,
    input [S_AXIS_IARG_21_DMWIDTH-1:0] s_axis_iarg_21_tdata,
    output s_axis_iarg_21_tready,
    input ap_axis_iarg_21_tready,
    output ap_axis_iarg_21_tlast,
    output ap_axis_iarg_21_tvalid,
    output [S_AXIS_IARG_21_WIDTH/8-1:0] ap_axis_iarg_21_tkeep,
    output [S_AXIS_IARG_21_WIDTH/8-1:0] ap_axis_iarg_21_tstrb,
    output [S_AXIS_IARG_21_WIDTH-1:0] ap_axis_iarg_21_tdata,
    //input AXI-Stream pass-through interface 22
    input s_axis_iarg_22_aclk,
    input s_axis_iarg_22_aresetn,
    input s_axis_iarg_22_tlast,
    input s_axis_iarg_22_tvalid,
    input [S_AXIS_IARG_22_DMWIDTH/8-1:0] s_axis_iarg_22_tkeep,
    input [S_AXIS_IARG_22_DMWIDTH/8-1:0] s_axis_iarg_22_tstrb,
    input [S_AXIS_IARG_22_DMWIDTH-1:0] s_axis_iarg_22_tdata,
    output s_axis_iarg_22_tready,
    input ap_axis_iarg_22_tready,
    output ap_axis_iarg_22_tlast,
    output ap_axis_iarg_22_tvalid,
    output [S_AXIS_IARG_22_WIDTH/8-1:0] ap_axis_iarg_22_tkeep,
    output [S_AXIS_IARG_22_WIDTH/8-1:0] ap_axis_iarg_22_tstrb,
    output [S_AXIS_IARG_22_WIDTH-1:0] ap_axis_iarg_22_tdata,
    //input AXI-Stream pass-through interface 23
    input s_axis_iarg_23_aclk,
    input s_axis_iarg_23_aresetn,
    input s_axis_iarg_23_tlast,
    input s_axis_iarg_23_tvalid,
    input [S_AXIS_IARG_23_DMWIDTH/8-1:0] s_axis_iarg_23_tkeep,
    input [S_AXIS_IARG_23_DMWIDTH/8-1:0] s_axis_iarg_23_tstrb,
    input [S_AXIS_IARG_23_DMWIDTH-1:0] s_axis_iarg_23_tdata,
    output s_axis_iarg_23_tready,
    input ap_axis_iarg_23_tready,
    output ap_axis_iarg_23_tlast,
    output ap_axis_iarg_23_tvalid,
    output [S_AXIS_IARG_23_WIDTH/8-1:0] ap_axis_iarg_23_tkeep,
    output [S_AXIS_IARG_23_WIDTH/8-1:0] ap_axis_iarg_23_tstrb,
    output [S_AXIS_IARG_23_WIDTH-1:0] ap_axis_iarg_23_tdata,
    //input AXI-Stream pass-through interface 24
    input s_axis_iarg_24_aclk,
    input s_axis_iarg_24_aresetn,
    input s_axis_iarg_24_tlast,
    input s_axis_iarg_24_tvalid,
    input [S_AXIS_IARG_24_DMWIDTH/8-1:0] s_axis_iarg_24_tkeep,
    input [S_AXIS_IARG_24_DMWIDTH/8-1:0] s_axis_iarg_24_tstrb,
    input [S_AXIS_IARG_24_DMWIDTH-1:0] s_axis_iarg_24_tdata,
    output s_axis_iarg_24_tready,
    input ap_axis_iarg_24_tready,
    output ap_axis_iarg_24_tlast,
    output ap_axis_iarg_24_tvalid,
    output [S_AXIS_IARG_24_WIDTH/8-1:0] ap_axis_iarg_24_tkeep,
    output [S_AXIS_IARG_24_WIDTH/8-1:0] ap_axis_iarg_24_tstrb,
    output [S_AXIS_IARG_24_WIDTH-1:0] ap_axis_iarg_24_tdata,
    //input AXI-Stream pass-through interface 25
    input s_axis_iarg_25_aclk,
    input s_axis_iarg_25_aresetn,
    input s_axis_iarg_25_tlast,
    input s_axis_iarg_25_tvalid,
    input [S_AXIS_IARG_25_DMWIDTH/8-1:0] s_axis_iarg_25_tkeep,
    input [S_AXIS_IARG_25_DMWIDTH/8-1:0] s_axis_iarg_25_tstrb,
    input [S_AXIS_IARG_25_DMWIDTH-1:0] s_axis_iarg_25_tdata,
    output s_axis_iarg_25_tready,
    input ap_axis_iarg_25_tready,
    output ap_axis_iarg_25_tlast,
    output ap_axis_iarg_25_tvalid,
    output [S_AXIS_IARG_25_WIDTH/8-1:0] ap_axis_iarg_25_tkeep,
    output [S_AXIS_IARG_25_WIDTH/8-1:0] ap_axis_iarg_25_tstrb,
    output [S_AXIS_IARG_25_WIDTH-1:0] ap_axis_iarg_25_tdata,
    //input AXI-Stream pass-through interface 26
    input s_axis_iarg_26_aclk,
    input s_axis_iarg_26_aresetn,
    input s_axis_iarg_26_tlast,
    input s_axis_iarg_26_tvalid,
    input [S_AXIS_IARG_26_DMWIDTH/8-1:0] s_axis_iarg_26_tkeep,
    input [S_AXIS_IARG_26_DMWIDTH/8-1:0] s_axis_iarg_26_tstrb,
    input [S_AXIS_IARG_26_DMWIDTH-1:0] s_axis_iarg_26_tdata,
    output s_axis_iarg_26_tready,
    input ap_axis_iarg_26_tready,
    output ap_axis_iarg_26_tlast,
    output ap_axis_iarg_26_tvalid,
    output [S_AXIS_IARG_26_WIDTH/8-1:0] ap_axis_iarg_26_tkeep,
    output [S_AXIS_IARG_26_WIDTH/8-1:0] ap_axis_iarg_26_tstrb,
    output [S_AXIS_IARG_26_WIDTH-1:0] ap_axis_iarg_26_tdata,
    //input AXI-Stream pass-through interface 27
    input s_axis_iarg_27_aclk,
    input s_axis_iarg_27_aresetn,
    input s_axis_iarg_27_tlast,
    input s_axis_iarg_27_tvalid,
    input [S_AXIS_IARG_27_DMWIDTH/8-1:0] s_axis_iarg_27_tkeep,
    input [S_AXIS_IARG_27_DMWIDTH/8-1:0] s_axis_iarg_27_tstrb,
    input [S_AXIS_IARG_27_DMWIDTH-1:0] s_axis_iarg_27_tdata,
    output s_axis_iarg_27_tready,
    input ap_axis_iarg_27_tready,
    output ap_axis_iarg_27_tlast,
    output ap_axis_iarg_27_tvalid,
    output [S_AXIS_IARG_27_WIDTH/8-1:0] ap_axis_iarg_27_tkeep,
    output [S_AXIS_IARG_27_WIDTH/8-1:0] ap_axis_iarg_27_tstrb,
    output [S_AXIS_IARG_27_WIDTH-1:0] ap_axis_iarg_27_tdata,
    //input AXI-Stream pass-through interface 28
    input s_axis_iarg_28_aclk,
    input s_axis_iarg_28_aresetn,
    input s_axis_iarg_28_tlast,
    input s_axis_iarg_28_tvalid,
    input [S_AXIS_IARG_28_DMWIDTH/8-1:0] s_axis_iarg_28_tkeep,
    input [S_AXIS_IARG_28_DMWIDTH/8-1:0] s_axis_iarg_28_tstrb,
    input [S_AXIS_IARG_28_DMWIDTH-1:0] s_axis_iarg_28_tdata,
    output s_axis_iarg_28_tready,
    input ap_axis_iarg_28_tready,
    output ap_axis_iarg_28_tlast,
    output ap_axis_iarg_28_tvalid,
    output [S_AXIS_IARG_28_WIDTH/8-1:0] ap_axis_iarg_28_tkeep,
    output [S_AXIS_IARG_28_WIDTH/8-1:0] ap_axis_iarg_28_tstrb,
    output [S_AXIS_IARG_28_WIDTH-1:0] ap_axis_iarg_28_tdata,
    //input AXI-Stream pass-through interface 29
    input s_axis_iarg_29_aclk,
    input s_axis_iarg_29_aresetn,
    input s_axis_iarg_29_tlast,
    input s_axis_iarg_29_tvalid,
    input [S_AXIS_IARG_29_DMWIDTH/8-1:0] s_axis_iarg_29_tkeep,
    input [S_AXIS_IARG_29_DMWIDTH/8-1:0] s_axis_iarg_29_tstrb,
    input [S_AXIS_IARG_29_DMWIDTH-1:0] s_axis_iarg_29_tdata,
    output s_axis_iarg_29_tready,
    input ap_axis_iarg_29_tready,
    output ap_axis_iarg_29_tlast,
    output ap_axis_iarg_29_tvalid,
    output [S_AXIS_IARG_29_WIDTH/8-1:0] ap_axis_iarg_29_tkeep,
    output [S_AXIS_IARG_29_WIDTH/8-1:0] ap_axis_iarg_29_tstrb,
    output [S_AXIS_IARG_29_WIDTH-1:0] ap_axis_iarg_29_tdata,
    //input AXI-Stream pass-through interface 30
    input s_axis_iarg_30_aclk,
    input s_axis_iarg_30_aresetn,
    input s_axis_iarg_30_tlast,
    input s_axis_iarg_30_tvalid,
    input [S_AXIS_IARG_30_DMWIDTH/8-1:0] s_axis_iarg_30_tkeep,
    input [S_AXIS_IARG_30_DMWIDTH/8-1:0] s_axis_iarg_30_tstrb,
    input [S_AXIS_IARG_30_DMWIDTH-1:0] s_axis_iarg_30_tdata,
    output s_axis_iarg_30_tready,
    input ap_axis_iarg_30_tready,
    output ap_axis_iarg_30_tlast,
    output ap_axis_iarg_30_tvalid,
    output [S_AXIS_IARG_30_WIDTH/8-1:0] ap_axis_iarg_30_tkeep,
    output [S_AXIS_IARG_30_WIDTH/8-1:0] ap_axis_iarg_30_tstrb,
    output [S_AXIS_IARG_30_WIDTH-1:0] ap_axis_iarg_30_tdata,
    //input AXI-Stream pass-through interface 31
    input s_axis_iarg_31_aclk,
    input s_axis_iarg_31_aresetn,
    input s_axis_iarg_31_tlast,
    input s_axis_iarg_31_tvalid,
    input [S_AXIS_IARG_31_DMWIDTH/8-1:0] s_axis_iarg_31_tkeep,
    input [S_AXIS_IARG_31_DMWIDTH/8-1:0] s_axis_iarg_31_tstrb,
    input [S_AXIS_IARG_31_DMWIDTH-1:0] s_axis_iarg_31_tdata,
    output s_axis_iarg_31_tready,
    input ap_axis_iarg_31_tready,
    output ap_axis_iarg_31_tlast,
    output ap_axis_iarg_31_tvalid,
    output [S_AXIS_IARG_31_WIDTH/8-1:0] ap_axis_iarg_31_tkeep,
    output [S_AXIS_IARG_31_WIDTH/8-1:0] ap_axis_iarg_31_tstrb,
    output [S_AXIS_IARG_31_WIDTH-1:0] ap_axis_iarg_31_tdata,
    //input AXI-Stream pass-through interface 32
    input s_axis_iarg_32_aclk,
    input s_axis_iarg_32_aresetn,
    input s_axis_iarg_32_tlast,
    input s_axis_iarg_32_tvalid,
    input [S_AXIS_IARG_32_DMWIDTH/8-1:0] s_axis_iarg_32_tkeep,
    input [S_AXIS_IARG_32_DMWIDTH/8-1:0] s_axis_iarg_32_tstrb,
    input [S_AXIS_IARG_32_DMWIDTH-1:0] s_axis_iarg_32_tdata,
    output s_axis_iarg_32_tready,
    input ap_axis_iarg_32_tready,
    output ap_axis_iarg_32_tlast,
    output ap_axis_iarg_32_tvalid,
    output [S_AXIS_IARG_32_WIDTH/8-1:0] ap_axis_iarg_32_tkeep,
    output [S_AXIS_IARG_32_WIDTH/8-1:0] ap_axis_iarg_32_tstrb,
    output [S_AXIS_IARG_32_WIDTH-1:0] ap_axis_iarg_32_tdata,
    //input AXI-Stream pass-through interface 33
    input s_axis_iarg_33_aclk,
    input s_axis_iarg_33_aresetn,
    input s_axis_iarg_33_tlast,
    input s_axis_iarg_33_tvalid,
    input [S_AXIS_IARG_33_DMWIDTH/8-1:0] s_axis_iarg_33_tkeep,
    input [S_AXIS_IARG_33_DMWIDTH/8-1:0] s_axis_iarg_33_tstrb,
    input [S_AXIS_IARG_33_DMWIDTH-1:0] s_axis_iarg_33_tdata,
    output s_axis_iarg_33_tready,
    input ap_axis_iarg_33_tready,
    output ap_axis_iarg_33_tlast,
    output ap_axis_iarg_33_tvalid,
    output [S_AXIS_IARG_33_WIDTH/8-1:0] ap_axis_iarg_33_tkeep,
    output [S_AXIS_IARG_33_WIDTH/8-1:0] ap_axis_iarg_33_tstrb,
    output [S_AXIS_IARG_33_WIDTH-1:0] ap_axis_iarg_33_tdata,
    //input AXI-Stream pass-through interface 34
    input s_axis_iarg_34_aclk,
    input s_axis_iarg_34_aresetn,
    input s_axis_iarg_34_tlast,
    input s_axis_iarg_34_tvalid,
    input [S_AXIS_IARG_34_DMWIDTH/8-1:0] s_axis_iarg_34_tkeep,
    input [S_AXIS_IARG_34_DMWIDTH/8-1:0] s_axis_iarg_34_tstrb,
    input [S_AXIS_IARG_34_DMWIDTH-1:0] s_axis_iarg_34_tdata,
    output s_axis_iarg_34_tready,
    input ap_axis_iarg_34_tready,
    output ap_axis_iarg_34_tlast,
    output ap_axis_iarg_34_tvalid,
    output [S_AXIS_IARG_34_WIDTH/8-1:0] ap_axis_iarg_34_tkeep,
    output [S_AXIS_IARG_34_WIDTH/8-1:0] ap_axis_iarg_34_tstrb,
    output [S_AXIS_IARG_34_WIDTH-1:0] ap_axis_iarg_34_tdata,
    //input AXI-Stream pass-through interface 35
    input s_axis_iarg_35_aclk,
    input s_axis_iarg_35_aresetn,
    input s_axis_iarg_35_tlast,
    input s_axis_iarg_35_tvalid,
    input [S_AXIS_IARG_35_DMWIDTH/8-1:0] s_axis_iarg_35_tkeep,
    input [S_AXIS_IARG_35_DMWIDTH/8-1:0] s_axis_iarg_35_tstrb,
    input [S_AXIS_IARG_35_DMWIDTH-1:0] s_axis_iarg_35_tdata,
    output s_axis_iarg_35_tready,
    input ap_axis_iarg_35_tready,
    output ap_axis_iarg_35_tlast,
    output ap_axis_iarg_35_tvalid,
    output [S_AXIS_IARG_35_WIDTH/8-1:0] ap_axis_iarg_35_tkeep,
    output [S_AXIS_IARG_35_WIDTH/8-1:0] ap_axis_iarg_35_tstrb,
    output [S_AXIS_IARG_35_WIDTH-1:0] ap_axis_iarg_35_tdata,
    //input AXI-Stream pass-through interface 36
    input s_axis_iarg_36_aclk,
    input s_axis_iarg_36_aresetn,
    input s_axis_iarg_36_tlast,
    input s_axis_iarg_36_tvalid,
    input [S_AXIS_IARG_36_DMWIDTH/8-1:0] s_axis_iarg_36_tkeep,
    input [S_AXIS_IARG_36_DMWIDTH/8-1:0] s_axis_iarg_36_tstrb,
    input [S_AXIS_IARG_36_DMWIDTH-1:0] s_axis_iarg_36_tdata,
    output s_axis_iarg_36_tready,
    input ap_axis_iarg_36_tready,
    output ap_axis_iarg_36_tlast,
    output ap_axis_iarg_36_tvalid,
    output [S_AXIS_IARG_36_WIDTH/8-1:0] ap_axis_iarg_36_tkeep,
    output [S_AXIS_IARG_36_WIDTH/8-1:0] ap_axis_iarg_36_tstrb,
    output [S_AXIS_IARG_36_WIDTH-1:0] ap_axis_iarg_36_tdata,
    //input AXI-Stream pass-through interface 37
    input s_axis_iarg_37_aclk,
    input s_axis_iarg_37_aresetn,
    input s_axis_iarg_37_tlast,
    input s_axis_iarg_37_tvalid,
    input [S_AXIS_IARG_37_DMWIDTH/8-1:0] s_axis_iarg_37_tkeep,
    input [S_AXIS_IARG_37_DMWIDTH/8-1:0] s_axis_iarg_37_tstrb,
    input [S_AXIS_IARG_37_DMWIDTH-1:0] s_axis_iarg_37_tdata,
    output s_axis_iarg_37_tready,
    input ap_axis_iarg_37_tready,
    output ap_axis_iarg_37_tlast,
    output ap_axis_iarg_37_tvalid,
    output [S_AXIS_IARG_37_WIDTH/8-1:0] ap_axis_iarg_37_tkeep,
    output [S_AXIS_IARG_37_WIDTH/8-1:0] ap_axis_iarg_37_tstrb,
    output [S_AXIS_IARG_37_WIDTH-1:0] ap_axis_iarg_37_tdata,
    //input AXI-Stream pass-through interface 38
    input s_axis_iarg_38_aclk,
    input s_axis_iarg_38_aresetn,
    input s_axis_iarg_38_tlast,
    input s_axis_iarg_38_tvalid,
    input [S_AXIS_IARG_38_DMWIDTH/8-1:0] s_axis_iarg_38_tkeep,
    input [S_AXIS_IARG_38_DMWIDTH/8-1:0] s_axis_iarg_38_tstrb,
    input [S_AXIS_IARG_38_DMWIDTH-1:0] s_axis_iarg_38_tdata,
    output s_axis_iarg_38_tready,
    input ap_axis_iarg_38_tready,
    output ap_axis_iarg_38_tlast,
    output ap_axis_iarg_38_tvalid,
    output [S_AXIS_IARG_38_WIDTH/8-1:0] ap_axis_iarg_38_tkeep,
    output [S_AXIS_IARG_38_WIDTH/8-1:0] ap_axis_iarg_38_tstrb,
    output [S_AXIS_IARG_38_WIDTH-1:0] ap_axis_iarg_38_tdata,
    //input AXI-Stream pass-through interface 39
    input s_axis_iarg_39_aclk,
    input s_axis_iarg_39_aresetn,
    input s_axis_iarg_39_tlast,
    input s_axis_iarg_39_tvalid,
    input [S_AXIS_IARG_39_DMWIDTH/8-1:0] s_axis_iarg_39_tkeep,
    input [S_AXIS_IARG_39_DMWIDTH/8-1:0] s_axis_iarg_39_tstrb,
    input [S_AXIS_IARG_39_DMWIDTH-1:0] s_axis_iarg_39_tdata,
    output s_axis_iarg_39_tready,
    input ap_axis_iarg_39_tready,
    output ap_axis_iarg_39_tlast,
    output ap_axis_iarg_39_tvalid,
    output [S_AXIS_IARG_39_WIDTH/8-1:0] ap_axis_iarg_39_tkeep,
    output [S_AXIS_IARG_39_WIDTH/8-1:0] ap_axis_iarg_39_tstrb,
    output [S_AXIS_IARG_39_WIDTH-1:0] ap_axis_iarg_39_tdata,
    //input AXI-Stream pass-through interface 40
    input s_axis_iarg_40_aclk,
    input s_axis_iarg_40_aresetn,
    input s_axis_iarg_40_tlast,
    input s_axis_iarg_40_tvalid,
    input [S_AXIS_IARG_40_DMWIDTH/8-1:0] s_axis_iarg_40_tkeep,
    input [S_AXIS_IARG_40_DMWIDTH/8-1:0] s_axis_iarg_40_tstrb,
    input [S_AXIS_IARG_40_DMWIDTH-1:0] s_axis_iarg_40_tdata,
    output s_axis_iarg_40_tready,
    input ap_axis_iarg_40_tready,
    output ap_axis_iarg_40_tlast,
    output ap_axis_iarg_40_tvalid,
    output [S_AXIS_IARG_40_WIDTH/8-1:0] ap_axis_iarg_40_tkeep,
    output [S_AXIS_IARG_40_WIDTH/8-1:0] ap_axis_iarg_40_tstrb,
    output [S_AXIS_IARG_40_WIDTH-1:0] ap_axis_iarg_40_tdata,
    //input AXI-Stream pass-through interface 41
    input s_axis_iarg_41_aclk,
    input s_axis_iarg_41_aresetn,
    input s_axis_iarg_41_tlast,
    input s_axis_iarg_41_tvalid,
    input [S_AXIS_IARG_41_DMWIDTH/8-1:0] s_axis_iarg_41_tkeep,
    input [S_AXIS_IARG_41_DMWIDTH/8-1:0] s_axis_iarg_41_tstrb,
    input [S_AXIS_IARG_41_DMWIDTH-1:0] s_axis_iarg_41_tdata,
    output s_axis_iarg_41_tready,
    input ap_axis_iarg_41_tready,
    output ap_axis_iarg_41_tlast,
    output ap_axis_iarg_41_tvalid,
    output [S_AXIS_IARG_41_WIDTH/8-1:0] ap_axis_iarg_41_tkeep,
    output [S_AXIS_IARG_41_WIDTH/8-1:0] ap_axis_iarg_41_tstrb,
    output [S_AXIS_IARG_41_WIDTH-1:0] ap_axis_iarg_41_tdata,
    //input AXI-Stream pass-through interface 42
    input s_axis_iarg_42_aclk,
    input s_axis_iarg_42_aresetn,
    input s_axis_iarg_42_tlast,
    input s_axis_iarg_42_tvalid,
    input [S_AXIS_IARG_42_DMWIDTH/8-1:0] s_axis_iarg_42_tkeep,
    input [S_AXIS_IARG_42_DMWIDTH/8-1:0] s_axis_iarg_42_tstrb,
    input [S_AXIS_IARG_42_DMWIDTH-1:0] s_axis_iarg_42_tdata,
    output s_axis_iarg_42_tready,
    input ap_axis_iarg_42_tready,
    output ap_axis_iarg_42_tlast,
    output ap_axis_iarg_42_tvalid,
    output [S_AXIS_IARG_42_WIDTH/8-1:0] ap_axis_iarg_42_tkeep,
    output [S_AXIS_IARG_42_WIDTH/8-1:0] ap_axis_iarg_42_tstrb,
    output [S_AXIS_IARG_42_WIDTH-1:0] ap_axis_iarg_42_tdata,
    //input AXI-Stream pass-through interface 43
    input s_axis_iarg_43_aclk,
    input s_axis_iarg_43_aresetn,
    input s_axis_iarg_43_tlast,
    input s_axis_iarg_43_tvalid,
    input [S_AXIS_IARG_43_DMWIDTH/8-1:0] s_axis_iarg_43_tkeep,
    input [S_AXIS_IARG_43_DMWIDTH/8-1:0] s_axis_iarg_43_tstrb,
    input [S_AXIS_IARG_43_DMWIDTH-1:0] s_axis_iarg_43_tdata,
    output s_axis_iarg_43_tready,
    input ap_axis_iarg_43_tready,
    output ap_axis_iarg_43_tlast,
    output ap_axis_iarg_43_tvalid,
    output [S_AXIS_IARG_43_WIDTH/8-1:0] ap_axis_iarg_43_tkeep,
    output [S_AXIS_IARG_43_WIDTH/8-1:0] ap_axis_iarg_43_tstrb,
    output [S_AXIS_IARG_43_WIDTH-1:0] ap_axis_iarg_43_tdata,
    //input AXI-Stream pass-through interface 44
    input s_axis_iarg_44_aclk,
    input s_axis_iarg_44_aresetn,
    input s_axis_iarg_44_tlast,
    input s_axis_iarg_44_tvalid,
    input [S_AXIS_IARG_44_DMWIDTH/8-1:0] s_axis_iarg_44_tkeep,
    input [S_AXIS_IARG_44_DMWIDTH/8-1:0] s_axis_iarg_44_tstrb,
    input [S_AXIS_IARG_44_DMWIDTH-1:0] s_axis_iarg_44_tdata,
    output s_axis_iarg_44_tready,
    input ap_axis_iarg_44_tready,
    output ap_axis_iarg_44_tlast,
    output ap_axis_iarg_44_tvalid,
    output [S_AXIS_IARG_44_WIDTH/8-1:0] ap_axis_iarg_44_tkeep,
    output [S_AXIS_IARG_44_WIDTH/8-1:0] ap_axis_iarg_44_tstrb,
    output [S_AXIS_IARG_44_WIDTH-1:0] ap_axis_iarg_44_tdata,
    //input AXI-Stream pass-through interface 45
    input s_axis_iarg_45_aclk,
    input s_axis_iarg_45_aresetn,
    input s_axis_iarg_45_tlast,
    input s_axis_iarg_45_tvalid,
    input [S_AXIS_IARG_45_DMWIDTH/8-1:0] s_axis_iarg_45_tkeep,
    input [S_AXIS_IARG_45_DMWIDTH/8-1:0] s_axis_iarg_45_tstrb,
    input [S_AXIS_IARG_45_DMWIDTH-1:0] s_axis_iarg_45_tdata,
    output s_axis_iarg_45_tready,
    input ap_axis_iarg_45_tready,
    output ap_axis_iarg_45_tlast,
    output ap_axis_iarg_45_tvalid,
    output [S_AXIS_IARG_45_WIDTH/8-1:0] ap_axis_iarg_45_tkeep,
    output [S_AXIS_IARG_45_WIDTH/8-1:0] ap_axis_iarg_45_tstrb,
    output [S_AXIS_IARG_45_WIDTH-1:0] ap_axis_iarg_45_tdata,
    //input AXI-Stream pass-through interface 46
    input s_axis_iarg_46_aclk,
    input s_axis_iarg_46_aresetn,
    input s_axis_iarg_46_tlast,
    input s_axis_iarg_46_tvalid,
    input [S_AXIS_IARG_46_DMWIDTH/8-1:0] s_axis_iarg_46_tkeep,
    input [S_AXIS_IARG_46_DMWIDTH/8-1:0] s_axis_iarg_46_tstrb,
    input [S_AXIS_IARG_46_DMWIDTH-1:0] s_axis_iarg_46_tdata,
    output s_axis_iarg_46_tready,
    input ap_axis_iarg_46_tready,
    output ap_axis_iarg_46_tlast,
    output ap_axis_iarg_46_tvalid,
    output [S_AXIS_IARG_46_WIDTH/8-1:0] ap_axis_iarg_46_tkeep,
    output [S_AXIS_IARG_46_WIDTH/8-1:0] ap_axis_iarg_46_tstrb,
    output [S_AXIS_IARG_46_WIDTH-1:0] ap_axis_iarg_46_tdata,
    //input AXI-Stream pass-through interface 47
    input s_axis_iarg_47_aclk,
    input s_axis_iarg_47_aresetn,
    input s_axis_iarg_47_tlast,
    input s_axis_iarg_47_tvalid,
    input [S_AXIS_IARG_47_DMWIDTH/8-1:0] s_axis_iarg_47_tkeep,
    input [S_AXIS_IARG_47_DMWIDTH/8-1:0] s_axis_iarg_47_tstrb,
    input [S_AXIS_IARG_47_DMWIDTH-1:0] s_axis_iarg_47_tdata,
    output s_axis_iarg_47_tready,
    input ap_axis_iarg_47_tready,
    output ap_axis_iarg_47_tlast,
    output ap_axis_iarg_47_tvalid,
    output [S_AXIS_IARG_47_WIDTH/8-1:0] ap_axis_iarg_47_tkeep,
    output [S_AXIS_IARG_47_WIDTH/8-1:0] ap_axis_iarg_47_tstrb,
    output [S_AXIS_IARG_47_WIDTH-1:0] ap_axis_iarg_47_tdata,
    //input AXI-Stream pass-through interface 48
    input s_axis_iarg_48_aclk,
    input s_axis_iarg_48_aresetn,
    input s_axis_iarg_48_tlast,
    input s_axis_iarg_48_tvalid,
    input [S_AXIS_IARG_48_DMWIDTH/8-1:0] s_axis_iarg_48_tkeep,
    input [S_AXIS_IARG_48_DMWIDTH/8-1:0] s_axis_iarg_48_tstrb,
    input [S_AXIS_IARG_48_DMWIDTH-1:0] s_axis_iarg_48_tdata,
    output s_axis_iarg_48_tready,
    input ap_axis_iarg_48_tready,
    output ap_axis_iarg_48_tlast,
    output ap_axis_iarg_48_tvalid,
    output [S_AXIS_IARG_48_WIDTH/8-1:0] ap_axis_iarg_48_tkeep,
    output [S_AXIS_IARG_48_WIDTH/8-1:0] ap_axis_iarg_48_tstrb,
    output [S_AXIS_IARG_48_WIDTH-1:0] ap_axis_iarg_48_tdata,
    //input AXI-Stream pass-through interface 49
    input s_axis_iarg_49_aclk,
    input s_axis_iarg_49_aresetn,
    input s_axis_iarg_49_tlast,
    input s_axis_iarg_49_tvalid,
    input [S_AXIS_IARG_49_DMWIDTH/8-1:0] s_axis_iarg_49_tkeep,
    input [S_AXIS_IARG_49_DMWIDTH/8-1:0] s_axis_iarg_49_tstrb,
    input [S_AXIS_IARG_49_DMWIDTH-1:0] s_axis_iarg_49_tdata,
    output s_axis_iarg_49_tready,
    input ap_axis_iarg_49_tready,
    output ap_axis_iarg_49_tlast,
    output ap_axis_iarg_49_tvalid,
    output [S_AXIS_IARG_49_WIDTH/8-1:0] ap_axis_iarg_49_tkeep,
    output [S_AXIS_IARG_49_WIDTH/8-1:0] ap_axis_iarg_49_tstrb,
    output [S_AXIS_IARG_49_WIDTH-1:0] ap_axis_iarg_49_tdata,
    //input AXI-Stream pass-through interface 50
    input s_axis_iarg_50_aclk,
    input s_axis_iarg_50_aresetn,
    input s_axis_iarg_50_tlast,
    input s_axis_iarg_50_tvalid,
    input [S_AXIS_IARG_50_DMWIDTH/8-1:0] s_axis_iarg_50_tkeep,
    input [S_AXIS_IARG_50_DMWIDTH/8-1:0] s_axis_iarg_50_tstrb,
    input [S_AXIS_IARG_50_DMWIDTH-1:0] s_axis_iarg_50_tdata,
    output s_axis_iarg_50_tready,
    input ap_axis_iarg_50_tready,
    output ap_axis_iarg_50_tlast,
    output ap_axis_iarg_50_tvalid,
    output [S_AXIS_IARG_50_WIDTH/8-1:0] ap_axis_iarg_50_tkeep,
    output [S_AXIS_IARG_50_WIDTH/8-1:0] ap_axis_iarg_50_tstrb,
    output [S_AXIS_IARG_50_WIDTH-1:0] ap_axis_iarg_50_tdata,
    //input AXI-Stream pass-through interface 51
    input s_axis_iarg_51_aclk,
    input s_axis_iarg_51_aresetn,
    input s_axis_iarg_51_tlast,
    input s_axis_iarg_51_tvalid,
    input [S_AXIS_IARG_51_DMWIDTH/8-1:0] s_axis_iarg_51_tkeep,
    input [S_AXIS_IARG_51_DMWIDTH/8-1:0] s_axis_iarg_51_tstrb,
    input [S_AXIS_IARG_51_DMWIDTH-1:0] s_axis_iarg_51_tdata,
    output s_axis_iarg_51_tready,
    input ap_axis_iarg_51_tready,
    output ap_axis_iarg_51_tlast,
    output ap_axis_iarg_51_tvalid,
    output [S_AXIS_IARG_51_WIDTH/8-1:0] ap_axis_iarg_51_tkeep,
    output [S_AXIS_IARG_51_WIDTH/8-1:0] ap_axis_iarg_51_tstrb,
    output [S_AXIS_IARG_51_WIDTH-1:0] ap_axis_iarg_51_tdata,
    //input AXI-Stream pass-through interface 52
    input s_axis_iarg_52_aclk,
    input s_axis_iarg_52_aresetn,
    input s_axis_iarg_52_tlast,
    input s_axis_iarg_52_tvalid,
    input [S_AXIS_IARG_52_DMWIDTH/8-1:0] s_axis_iarg_52_tkeep,
    input [S_AXIS_IARG_52_DMWIDTH/8-1:0] s_axis_iarg_52_tstrb,
    input [S_AXIS_IARG_52_DMWIDTH-1:0] s_axis_iarg_52_tdata,
    output s_axis_iarg_52_tready,
    input ap_axis_iarg_52_tready,
    output ap_axis_iarg_52_tlast,
    output ap_axis_iarg_52_tvalid,
    output [S_AXIS_IARG_52_WIDTH/8-1:0] ap_axis_iarg_52_tkeep,
    output [S_AXIS_IARG_52_WIDTH/8-1:0] ap_axis_iarg_52_tstrb,
    output [S_AXIS_IARG_52_WIDTH-1:0] ap_axis_iarg_52_tdata,
    //input AXI-Stream pass-through interface 53
    input s_axis_iarg_53_aclk,
    input s_axis_iarg_53_aresetn,
    input s_axis_iarg_53_tlast,
    input s_axis_iarg_53_tvalid,
    input [S_AXIS_IARG_53_DMWIDTH/8-1:0] s_axis_iarg_53_tkeep,
    input [S_AXIS_IARG_53_DMWIDTH/8-1:0] s_axis_iarg_53_tstrb,
    input [S_AXIS_IARG_53_DMWIDTH-1:0] s_axis_iarg_53_tdata,
    output s_axis_iarg_53_tready,
    input ap_axis_iarg_53_tready,
    output ap_axis_iarg_53_tlast,
    output ap_axis_iarg_53_tvalid,
    output [S_AXIS_IARG_53_WIDTH/8-1:0] ap_axis_iarg_53_tkeep,
    output [S_AXIS_IARG_53_WIDTH/8-1:0] ap_axis_iarg_53_tstrb,
    output [S_AXIS_IARG_53_WIDTH-1:0] ap_axis_iarg_53_tdata,
    //input AXI-Stream pass-through interface 54
    input s_axis_iarg_54_aclk,
    input s_axis_iarg_54_aresetn,
    input s_axis_iarg_54_tlast,
    input s_axis_iarg_54_tvalid,
    input [S_AXIS_IARG_54_DMWIDTH/8-1:0] s_axis_iarg_54_tkeep,
    input [S_AXIS_IARG_54_DMWIDTH/8-1:0] s_axis_iarg_54_tstrb,
    input [S_AXIS_IARG_54_DMWIDTH-1:0] s_axis_iarg_54_tdata,
    output s_axis_iarg_54_tready,
    input ap_axis_iarg_54_tready,
    output ap_axis_iarg_54_tlast,
    output ap_axis_iarg_54_tvalid,
    output [S_AXIS_IARG_54_WIDTH/8-1:0] ap_axis_iarg_54_tkeep,
    output [S_AXIS_IARG_54_WIDTH/8-1:0] ap_axis_iarg_54_tstrb,
    output [S_AXIS_IARG_54_WIDTH-1:0] ap_axis_iarg_54_tdata,
    //input AXI-Stream pass-through interface 55
    input s_axis_iarg_55_aclk,
    input s_axis_iarg_55_aresetn,
    input s_axis_iarg_55_tlast,
    input s_axis_iarg_55_tvalid,
    input [S_AXIS_IARG_55_DMWIDTH/8-1:0] s_axis_iarg_55_tkeep,
    input [S_AXIS_IARG_55_DMWIDTH/8-1:0] s_axis_iarg_55_tstrb,
    input [S_AXIS_IARG_55_DMWIDTH-1:0] s_axis_iarg_55_tdata,
    output s_axis_iarg_55_tready,
    input ap_axis_iarg_55_tready,
    output ap_axis_iarg_55_tlast,
    output ap_axis_iarg_55_tvalid,
    output [S_AXIS_IARG_55_WIDTH/8-1:0] ap_axis_iarg_55_tkeep,
    output [S_AXIS_IARG_55_WIDTH/8-1:0] ap_axis_iarg_55_tstrb,
    output [S_AXIS_IARG_55_WIDTH-1:0] ap_axis_iarg_55_tdata,
    //input AXI-Stream pass-through interface 56
    input s_axis_iarg_56_aclk,
    input s_axis_iarg_56_aresetn,
    input s_axis_iarg_56_tlast,
    input s_axis_iarg_56_tvalid,
    input [S_AXIS_IARG_56_DMWIDTH/8-1:0] s_axis_iarg_56_tkeep,
    input [S_AXIS_IARG_56_DMWIDTH/8-1:0] s_axis_iarg_56_tstrb,
    input [S_AXIS_IARG_56_DMWIDTH-1:0] s_axis_iarg_56_tdata,
    output s_axis_iarg_56_tready,
    input ap_axis_iarg_56_tready,
    output ap_axis_iarg_56_tlast,
    output ap_axis_iarg_56_tvalid,
    output [S_AXIS_IARG_56_WIDTH/8-1:0] ap_axis_iarg_56_tkeep,
    output [S_AXIS_IARG_56_WIDTH/8-1:0] ap_axis_iarg_56_tstrb,
    output [S_AXIS_IARG_56_WIDTH-1:0] ap_axis_iarg_56_tdata,
    //input AXI-Stream pass-through interface 57
    input s_axis_iarg_57_aclk,
    input s_axis_iarg_57_aresetn,
    input s_axis_iarg_57_tlast,
    input s_axis_iarg_57_tvalid,
    input [S_AXIS_IARG_57_DMWIDTH/8-1:0] s_axis_iarg_57_tkeep,
    input [S_AXIS_IARG_57_DMWIDTH/8-1:0] s_axis_iarg_57_tstrb,
    input [S_AXIS_IARG_57_DMWIDTH-1:0] s_axis_iarg_57_tdata,
    output s_axis_iarg_57_tready,
    input ap_axis_iarg_57_tready,
    output ap_axis_iarg_57_tlast,
    output ap_axis_iarg_57_tvalid,
    output [S_AXIS_IARG_57_WIDTH/8-1:0] ap_axis_iarg_57_tkeep,
    output [S_AXIS_IARG_57_WIDTH/8-1:0] ap_axis_iarg_57_tstrb,
    output [S_AXIS_IARG_57_WIDTH-1:0] ap_axis_iarg_57_tdata,
    //input AXI-Stream pass-through interface 58
    input s_axis_iarg_58_aclk,
    input s_axis_iarg_58_aresetn,
    input s_axis_iarg_58_tlast,
    input s_axis_iarg_58_tvalid,
    input [S_AXIS_IARG_58_DMWIDTH/8-1:0] s_axis_iarg_58_tkeep,
    input [S_AXIS_IARG_58_DMWIDTH/8-1:0] s_axis_iarg_58_tstrb,
    input [S_AXIS_IARG_58_DMWIDTH-1:0] s_axis_iarg_58_tdata,
    output s_axis_iarg_58_tready,
    input ap_axis_iarg_58_tready,
    output ap_axis_iarg_58_tlast,
    output ap_axis_iarg_58_tvalid,
    output [S_AXIS_IARG_58_WIDTH/8-1:0] ap_axis_iarg_58_tkeep,
    output [S_AXIS_IARG_58_WIDTH/8-1:0] ap_axis_iarg_58_tstrb,
    output [S_AXIS_IARG_58_WIDTH-1:0] ap_axis_iarg_58_tdata,
    //input AXI-Stream pass-through interface 59
    input s_axis_iarg_59_aclk,
    input s_axis_iarg_59_aresetn,
    input s_axis_iarg_59_tlast,
    input s_axis_iarg_59_tvalid,
    input [S_AXIS_IARG_59_DMWIDTH/8-1:0] s_axis_iarg_59_tkeep,
    input [S_AXIS_IARG_59_DMWIDTH/8-1:0] s_axis_iarg_59_tstrb,
    input [S_AXIS_IARG_59_DMWIDTH-1:0] s_axis_iarg_59_tdata,
    output s_axis_iarg_59_tready,
    input ap_axis_iarg_59_tready,
    output ap_axis_iarg_59_tlast,
    output ap_axis_iarg_59_tvalid,
    output [S_AXIS_IARG_59_WIDTH/8-1:0] ap_axis_iarg_59_tkeep,
    output [S_AXIS_IARG_59_WIDTH/8-1:0] ap_axis_iarg_59_tstrb,
    output [S_AXIS_IARG_59_WIDTH-1:0] ap_axis_iarg_59_tdata,
    //input AXI-Stream pass-through interface 60
    input s_axis_iarg_60_aclk,
    input s_axis_iarg_60_aresetn,
    input s_axis_iarg_60_tlast,
    input s_axis_iarg_60_tvalid,
    input [S_AXIS_IARG_60_DMWIDTH/8-1:0] s_axis_iarg_60_tkeep,
    input [S_AXIS_IARG_60_DMWIDTH/8-1:0] s_axis_iarg_60_tstrb,
    input [S_AXIS_IARG_60_DMWIDTH-1:0] s_axis_iarg_60_tdata,
    output s_axis_iarg_60_tready,
    input ap_axis_iarg_60_tready,
    output ap_axis_iarg_60_tlast,
    output ap_axis_iarg_60_tvalid,
    output [S_AXIS_IARG_60_WIDTH/8-1:0] ap_axis_iarg_60_tkeep,
    output [S_AXIS_IARG_60_WIDTH/8-1:0] ap_axis_iarg_60_tstrb,
    output [S_AXIS_IARG_60_WIDTH-1:0] ap_axis_iarg_60_tdata,
    //input AXI-Stream pass-through interface 61
    input s_axis_iarg_61_aclk,
    input s_axis_iarg_61_aresetn,
    input s_axis_iarg_61_tlast,
    input s_axis_iarg_61_tvalid,
    input [S_AXIS_IARG_61_DMWIDTH/8-1:0] s_axis_iarg_61_tkeep,
    input [S_AXIS_IARG_61_DMWIDTH/8-1:0] s_axis_iarg_61_tstrb,
    input [S_AXIS_IARG_61_DMWIDTH-1:0] s_axis_iarg_61_tdata,
    output s_axis_iarg_61_tready,
    input ap_axis_iarg_61_tready,
    output ap_axis_iarg_61_tlast,
    output ap_axis_iarg_61_tvalid,
    output [S_AXIS_IARG_61_WIDTH/8-1:0] ap_axis_iarg_61_tkeep,
    output [S_AXIS_IARG_61_WIDTH/8-1:0] ap_axis_iarg_61_tstrb,
    output [S_AXIS_IARG_61_WIDTH-1:0] ap_axis_iarg_61_tdata,
    //input AXI-Stream pass-through interface 62
    input s_axis_iarg_62_aclk,
    input s_axis_iarg_62_aresetn,
    input s_axis_iarg_62_tlast,
    input s_axis_iarg_62_tvalid,
    input [S_AXIS_IARG_62_DMWIDTH/8-1:0] s_axis_iarg_62_tkeep,
    input [S_AXIS_IARG_62_DMWIDTH/8-1:0] s_axis_iarg_62_tstrb,
    input [S_AXIS_IARG_62_DMWIDTH-1:0] s_axis_iarg_62_tdata,
    output s_axis_iarg_62_tready,
    input ap_axis_iarg_62_tready,
    output ap_axis_iarg_62_tlast,
    output ap_axis_iarg_62_tvalid,
    output [S_AXIS_IARG_62_WIDTH/8-1:0] ap_axis_iarg_62_tkeep,
    output [S_AXIS_IARG_62_WIDTH/8-1:0] ap_axis_iarg_62_tstrb,
    output [S_AXIS_IARG_62_WIDTH-1:0] ap_axis_iarg_62_tdata,
    //input AXI-Stream pass-through interface 63
    input s_axis_iarg_63_aclk,
    input s_axis_iarg_63_aresetn,
    input s_axis_iarg_63_tlast,
    input s_axis_iarg_63_tvalid,
    input [S_AXIS_IARG_63_DMWIDTH/8-1:0] s_axis_iarg_63_tkeep,
    input [S_AXIS_IARG_63_DMWIDTH/8-1:0] s_axis_iarg_63_tstrb,
    input [S_AXIS_IARG_63_DMWIDTH-1:0] s_axis_iarg_63_tdata,
    output s_axis_iarg_63_tready,
    input ap_axis_iarg_63_tready,
    output ap_axis_iarg_63_tlast,
    output ap_axis_iarg_63_tvalid,
    output [S_AXIS_IARG_63_WIDTH/8-1:0] ap_axis_iarg_63_tkeep,
    output [S_AXIS_IARG_63_WIDTH/8-1:0] ap_axis_iarg_63_tstrb,
    output [S_AXIS_IARG_63_WIDTH-1:0] ap_axis_iarg_63_tdata,
    //input AXI-Stream pass-through interface 64
    input s_axis_iarg_64_aclk,
    input s_axis_iarg_64_aresetn,
    input s_axis_iarg_64_tlast,
    input s_axis_iarg_64_tvalid,
    input [S_AXIS_IARG_64_DMWIDTH/8-1:0] s_axis_iarg_64_tkeep,
    input [S_AXIS_IARG_64_DMWIDTH/8-1:0] s_axis_iarg_64_tstrb,
    input [S_AXIS_IARG_64_DMWIDTH-1:0] s_axis_iarg_64_tdata,
    output s_axis_iarg_64_tready,
    input ap_axis_iarg_64_tready,
    output ap_axis_iarg_64_tlast,
    output ap_axis_iarg_64_tvalid,
    output [S_AXIS_IARG_64_WIDTH/8-1:0] ap_axis_iarg_64_tkeep,
    output [S_AXIS_IARG_64_WIDTH/8-1:0] ap_axis_iarg_64_tstrb,
    output [S_AXIS_IARG_64_WIDTH-1:0] ap_axis_iarg_64_tdata,
    //input AXI-Stream pass-through interface 65
    input s_axis_iarg_65_aclk,
    input s_axis_iarg_65_aresetn,
    input s_axis_iarg_65_tlast,
    input s_axis_iarg_65_tvalid,
    input [S_AXIS_IARG_65_DMWIDTH/8-1:0] s_axis_iarg_65_tkeep,
    input [S_AXIS_IARG_65_DMWIDTH/8-1:0] s_axis_iarg_65_tstrb,
    input [S_AXIS_IARG_65_DMWIDTH-1:0] s_axis_iarg_65_tdata,
    output s_axis_iarg_65_tready,
    input ap_axis_iarg_65_tready,
    output ap_axis_iarg_65_tlast,
    output ap_axis_iarg_65_tvalid,
    output [S_AXIS_IARG_65_WIDTH/8-1:0] ap_axis_iarg_65_tkeep,
    output [S_AXIS_IARG_65_WIDTH/8-1:0] ap_axis_iarg_65_tstrb,
    output [S_AXIS_IARG_65_WIDTH-1:0] ap_axis_iarg_65_tdata,
    //input AXI-Stream pass-through interface 66
    input s_axis_iarg_66_aclk,
    input s_axis_iarg_66_aresetn,
    input s_axis_iarg_66_tlast,
    input s_axis_iarg_66_tvalid,
    input [S_AXIS_IARG_66_DMWIDTH/8-1:0] s_axis_iarg_66_tkeep,
    input [S_AXIS_IARG_66_DMWIDTH/8-1:0] s_axis_iarg_66_tstrb,
    input [S_AXIS_IARG_66_DMWIDTH-1:0] s_axis_iarg_66_tdata,
    output s_axis_iarg_66_tready,
    input ap_axis_iarg_66_tready,
    output ap_axis_iarg_66_tlast,
    output ap_axis_iarg_66_tvalid,
    output [S_AXIS_IARG_66_WIDTH/8-1:0] ap_axis_iarg_66_tkeep,
    output [S_AXIS_IARG_66_WIDTH/8-1:0] ap_axis_iarg_66_tstrb,
    output [S_AXIS_IARG_66_WIDTH-1:0] ap_axis_iarg_66_tdata,
    //input AXI-Stream pass-through interface 67
    input s_axis_iarg_67_aclk,
    input s_axis_iarg_67_aresetn,
    input s_axis_iarg_67_tlast,
    input s_axis_iarg_67_tvalid,
    input [S_AXIS_IARG_67_DMWIDTH/8-1:0] s_axis_iarg_67_tkeep,
    input [S_AXIS_IARG_67_DMWIDTH/8-1:0] s_axis_iarg_67_tstrb,
    input [S_AXIS_IARG_67_DMWIDTH-1:0] s_axis_iarg_67_tdata,
    output s_axis_iarg_67_tready,
    input ap_axis_iarg_67_tready,
    output ap_axis_iarg_67_tlast,
    output ap_axis_iarg_67_tvalid,
    output [S_AXIS_IARG_67_WIDTH/8-1:0] ap_axis_iarg_67_tkeep,
    output [S_AXIS_IARG_67_WIDTH/8-1:0] ap_axis_iarg_67_tstrb,
    output [S_AXIS_IARG_67_WIDTH-1:0] ap_axis_iarg_67_tdata,
    //input AXI-Stream pass-through interface 68
    input s_axis_iarg_68_aclk,
    input s_axis_iarg_68_aresetn,
    input s_axis_iarg_68_tlast,
    input s_axis_iarg_68_tvalid,
    input [S_AXIS_IARG_68_DMWIDTH/8-1:0] s_axis_iarg_68_tkeep,
    input [S_AXIS_IARG_68_DMWIDTH/8-1:0] s_axis_iarg_68_tstrb,
    input [S_AXIS_IARG_68_DMWIDTH-1:0] s_axis_iarg_68_tdata,
    output s_axis_iarg_68_tready,
    input ap_axis_iarg_68_tready,
    output ap_axis_iarg_68_tlast,
    output ap_axis_iarg_68_tvalid,
    output [S_AXIS_IARG_68_WIDTH/8-1:0] ap_axis_iarg_68_tkeep,
    output [S_AXIS_IARG_68_WIDTH/8-1:0] ap_axis_iarg_68_tstrb,
    output [S_AXIS_IARG_68_WIDTH-1:0] ap_axis_iarg_68_tdata,
    //input AXI-Stream pass-through interface 69
    input s_axis_iarg_69_aclk,
    input s_axis_iarg_69_aresetn,
    input s_axis_iarg_69_tlast,
    input s_axis_iarg_69_tvalid,
    input [S_AXIS_IARG_69_DMWIDTH/8-1:0] s_axis_iarg_69_tkeep,
    input [S_AXIS_IARG_69_DMWIDTH/8-1:0] s_axis_iarg_69_tstrb,
    input [S_AXIS_IARG_69_DMWIDTH-1:0] s_axis_iarg_69_tdata,
    output s_axis_iarg_69_tready,
    input ap_axis_iarg_69_tready,
    output ap_axis_iarg_69_tlast,
    output ap_axis_iarg_69_tvalid,
    output [S_AXIS_IARG_69_WIDTH/8-1:0] ap_axis_iarg_69_tkeep,
    output [S_AXIS_IARG_69_WIDTH/8-1:0] ap_axis_iarg_69_tstrb,
    output [S_AXIS_IARG_69_WIDTH-1:0] ap_axis_iarg_69_tdata,
    //input AXI-Stream pass-through interface 70
    input s_axis_iarg_70_aclk,
    input s_axis_iarg_70_aresetn,
    input s_axis_iarg_70_tlast,
    input s_axis_iarg_70_tvalid,
    input [S_AXIS_IARG_70_DMWIDTH/8-1:0] s_axis_iarg_70_tkeep,
    input [S_AXIS_IARG_70_DMWIDTH/8-1:0] s_axis_iarg_70_tstrb,
    input [S_AXIS_IARG_70_DMWIDTH-1:0] s_axis_iarg_70_tdata,
    output s_axis_iarg_70_tready,
    input ap_axis_iarg_70_tready,
    output ap_axis_iarg_70_tlast,
    output ap_axis_iarg_70_tvalid,
    output [S_AXIS_IARG_70_WIDTH/8-1:0] ap_axis_iarg_70_tkeep,
    output [S_AXIS_IARG_70_WIDTH/8-1:0] ap_axis_iarg_70_tstrb,
    output [S_AXIS_IARG_70_WIDTH-1:0] ap_axis_iarg_70_tdata,
    //input AXI-Stream pass-through interface 71
    input s_axis_iarg_71_aclk,
    input s_axis_iarg_71_aresetn,
    input s_axis_iarg_71_tlast,
    input s_axis_iarg_71_tvalid,
    input [S_AXIS_IARG_71_DMWIDTH/8-1:0] s_axis_iarg_71_tkeep,
    input [S_AXIS_IARG_71_DMWIDTH/8-1:0] s_axis_iarg_71_tstrb,
    input [S_AXIS_IARG_71_DMWIDTH-1:0] s_axis_iarg_71_tdata,
    output s_axis_iarg_71_tready,
    input ap_axis_iarg_71_tready,
    output ap_axis_iarg_71_tlast,
    output ap_axis_iarg_71_tvalid,
    output [S_AXIS_IARG_71_WIDTH/8-1:0] ap_axis_iarg_71_tkeep,
    output [S_AXIS_IARG_71_WIDTH/8-1:0] ap_axis_iarg_71_tstrb,
    output [S_AXIS_IARG_71_WIDTH-1:0] ap_axis_iarg_71_tdata,
    //input AXI-Stream pass-through interface 72
    input s_axis_iarg_72_aclk,
    input s_axis_iarg_72_aresetn,
    input s_axis_iarg_72_tlast,
    input s_axis_iarg_72_tvalid,
    input [S_AXIS_IARG_72_DMWIDTH/8-1:0] s_axis_iarg_72_tkeep,
    input [S_AXIS_IARG_72_DMWIDTH/8-1:0] s_axis_iarg_72_tstrb,
    input [S_AXIS_IARG_72_DMWIDTH-1:0] s_axis_iarg_72_tdata,
    output s_axis_iarg_72_tready,
    input ap_axis_iarg_72_tready,
    output ap_axis_iarg_72_tlast,
    output ap_axis_iarg_72_tvalid,
    output [S_AXIS_IARG_72_WIDTH/8-1:0] ap_axis_iarg_72_tkeep,
    output [S_AXIS_IARG_72_WIDTH/8-1:0] ap_axis_iarg_72_tstrb,
    output [S_AXIS_IARG_72_WIDTH-1:0] ap_axis_iarg_72_tdata,
    //input AXI-Stream pass-through interface 73
    input s_axis_iarg_73_aclk,
    input s_axis_iarg_73_aresetn,
    input s_axis_iarg_73_tlast,
    input s_axis_iarg_73_tvalid,
    input [S_AXIS_IARG_73_DMWIDTH/8-1:0] s_axis_iarg_73_tkeep,
    input [S_AXIS_IARG_73_DMWIDTH/8-1:0] s_axis_iarg_73_tstrb,
    input [S_AXIS_IARG_73_DMWIDTH-1:0] s_axis_iarg_73_tdata,
    output s_axis_iarg_73_tready,
    input ap_axis_iarg_73_tready,
    output ap_axis_iarg_73_tlast,
    output ap_axis_iarg_73_tvalid,
    output [S_AXIS_IARG_73_WIDTH/8-1:0] ap_axis_iarg_73_tkeep,
    output [S_AXIS_IARG_73_WIDTH/8-1:0] ap_axis_iarg_73_tstrb,
    output [S_AXIS_IARG_73_WIDTH-1:0] ap_axis_iarg_73_tdata,
    //input AXI-Stream pass-through interface 74
    input s_axis_iarg_74_aclk,
    input s_axis_iarg_74_aresetn,
    input s_axis_iarg_74_tlast,
    input s_axis_iarg_74_tvalid,
    input [S_AXIS_IARG_74_DMWIDTH/8-1:0] s_axis_iarg_74_tkeep,
    input [S_AXIS_IARG_74_DMWIDTH/8-1:0] s_axis_iarg_74_tstrb,
    input [S_AXIS_IARG_74_DMWIDTH-1:0] s_axis_iarg_74_tdata,
    output s_axis_iarg_74_tready,
    input ap_axis_iarg_74_tready,
    output ap_axis_iarg_74_tlast,
    output ap_axis_iarg_74_tvalid,
    output [S_AXIS_IARG_74_WIDTH/8-1:0] ap_axis_iarg_74_tkeep,
    output [S_AXIS_IARG_74_WIDTH/8-1:0] ap_axis_iarg_74_tstrb,
    output [S_AXIS_IARG_74_WIDTH-1:0] ap_axis_iarg_74_tdata,
    //input AXI-Stream pass-through interface 75
    input s_axis_iarg_75_aclk,
    input s_axis_iarg_75_aresetn,
    input s_axis_iarg_75_tlast,
    input s_axis_iarg_75_tvalid,
    input [S_AXIS_IARG_75_DMWIDTH/8-1:0] s_axis_iarg_75_tkeep,
    input [S_AXIS_IARG_75_DMWIDTH/8-1:0] s_axis_iarg_75_tstrb,
    input [S_AXIS_IARG_75_DMWIDTH-1:0] s_axis_iarg_75_tdata,
    output s_axis_iarg_75_tready,
    input ap_axis_iarg_75_tready,
    output ap_axis_iarg_75_tlast,
    output ap_axis_iarg_75_tvalid,
    output [S_AXIS_IARG_75_WIDTH/8-1:0] ap_axis_iarg_75_tkeep,
    output [S_AXIS_IARG_75_WIDTH/8-1:0] ap_axis_iarg_75_tstrb,
    output [S_AXIS_IARG_75_WIDTH-1:0] ap_axis_iarg_75_tdata,
    //input AXI-Stream pass-through interface 76
    input s_axis_iarg_76_aclk,
    input s_axis_iarg_76_aresetn,
    input s_axis_iarg_76_tlast,
    input s_axis_iarg_76_tvalid,
    input [S_AXIS_IARG_76_DMWIDTH/8-1:0] s_axis_iarg_76_tkeep,
    input [S_AXIS_IARG_76_DMWIDTH/8-1:0] s_axis_iarg_76_tstrb,
    input [S_AXIS_IARG_76_DMWIDTH-1:0] s_axis_iarg_76_tdata,
    output s_axis_iarg_76_tready,
    input ap_axis_iarg_76_tready,
    output ap_axis_iarg_76_tlast,
    output ap_axis_iarg_76_tvalid,
    output [S_AXIS_IARG_76_WIDTH/8-1:0] ap_axis_iarg_76_tkeep,
    output [S_AXIS_IARG_76_WIDTH/8-1:0] ap_axis_iarg_76_tstrb,
    output [S_AXIS_IARG_76_WIDTH-1:0] ap_axis_iarg_76_tdata,
    //input AXI-Stream pass-through interface 77
    input s_axis_iarg_77_aclk,
    input s_axis_iarg_77_aresetn,
    input s_axis_iarg_77_tlast,
    input s_axis_iarg_77_tvalid,
    input [S_AXIS_IARG_77_DMWIDTH/8-1:0] s_axis_iarg_77_tkeep,
    input [S_AXIS_IARG_77_DMWIDTH/8-1:0] s_axis_iarg_77_tstrb,
    input [S_AXIS_IARG_77_DMWIDTH-1:0] s_axis_iarg_77_tdata,
    output s_axis_iarg_77_tready,
    input ap_axis_iarg_77_tready,
    output ap_axis_iarg_77_tlast,
    output ap_axis_iarg_77_tvalid,
    output [S_AXIS_IARG_77_WIDTH/8-1:0] ap_axis_iarg_77_tkeep,
    output [S_AXIS_IARG_77_WIDTH/8-1:0] ap_axis_iarg_77_tstrb,
    output [S_AXIS_IARG_77_WIDTH-1:0] ap_axis_iarg_77_tdata,
    //input AXI-Stream pass-through interface 78
    input s_axis_iarg_78_aclk,
    input s_axis_iarg_78_aresetn,
    input s_axis_iarg_78_tlast,
    input s_axis_iarg_78_tvalid,
    input [S_AXIS_IARG_78_DMWIDTH/8-1:0] s_axis_iarg_78_tkeep,
    input [S_AXIS_IARG_78_DMWIDTH/8-1:0] s_axis_iarg_78_tstrb,
    input [S_AXIS_IARG_78_DMWIDTH-1:0] s_axis_iarg_78_tdata,
    output s_axis_iarg_78_tready,
    input ap_axis_iarg_78_tready,
    output ap_axis_iarg_78_tlast,
    output ap_axis_iarg_78_tvalid,
    output [S_AXIS_IARG_78_WIDTH/8-1:0] ap_axis_iarg_78_tkeep,
    output [S_AXIS_IARG_78_WIDTH/8-1:0] ap_axis_iarg_78_tstrb,
    output [S_AXIS_IARG_78_WIDTH-1:0] ap_axis_iarg_78_tdata,
    //input AXI-Stream pass-through interface 79
    input s_axis_iarg_79_aclk,
    input s_axis_iarg_79_aresetn,
    input s_axis_iarg_79_tlast,
    input s_axis_iarg_79_tvalid,
    input [S_AXIS_IARG_79_DMWIDTH/8-1:0] s_axis_iarg_79_tkeep,
    input [S_AXIS_IARG_79_DMWIDTH/8-1:0] s_axis_iarg_79_tstrb,
    input [S_AXIS_IARG_79_DMWIDTH-1:0] s_axis_iarg_79_tdata,
    output s_axis_iarg_79_tready,
    input ap_axis_iarg_79_tready,
    output ap_axis_iarg_79_tlast,
    output ap_axis_iarg_79_tvalid,
    output [S_AXIS_IARG_79_WIDTH/8-1:0] ap_axis_iarg_79_tkeep,
    output [S_AXIS_IARG_79_WIDTH/8-1:0] ap_axis_iarg_79_tstrb,
    output [S_AXIS_IARG_79_WIDTH-1:0] ap_axis_iarg_79_tdata,
    //input AXI-Stream pass-through interface 80
    input s_axis_iarg_80_aclk,
    input s_axis_iarg_80_aresetn,
    input s_axis_iarg_80_tlast,
    input s_axis_iarg_80_tvalid,
    input [S_AXIS_IARG_80_DMWIDTH/8-1:0] s_axis_iarg_80_tkeep,
    input [S_AXIS_IARG_80_DMWIDTH/8-1:0] s_axis_iarg_80_tstrb,
    input [S_AXIS_IARG_80_DMWIDTH-1:0] s_axis_iarg_80_tdata,
    output s_axis_iarg_80_tready,
    input ap_axis_iarg_80_tready,
    output ap_axis_iarg_80_tlast,
    output ap_axis_iarg_80_tvalid,
    output [S_AXIS_IARG_80_WIDTH/8-1:0] ap_axis_iarg_80_tkeep,
    output [S_AXIS_IARG_80_WIDTH/8-1:0] ap_axis_iarg_80_tstrb,
    output [S_AXIS_IARG_80_WIDTH-1:0] ap_axis_iarg_80_tdata,
    //input AXI-Stream pass-through interface 81
    input s_axis_iarg_81_aclk,
    input s_axis_iarg_81_aresetn,
    input s_axis_iarg_81_tlast,
    input s_axis_iarg_81_tvalid,
    input [S_AXIS_IARG_81_DMWIDTH/8-1:0] s_axis_iarg_81_tkeep,
    input [S_AXIS_IARG_81_DMWIDTH/8-1:0] s_axis_iarg_81_tstrb,
    input [S_AXIS_IARG_81_DMWIDTH-1:0] s_axis_iarg_81_tdata,
    output s_axis_iarg_81_tready,
    input ap_axis_iarg_81_tready,
    output ap_axis_iarg_81_tlast,
    output ap_axis_iarg_81_tvalid,
    output [S_AXIS_IARG_81_WIDTH/8-1:0] ap_axis_iarg_81_tkeep,
    output [S_AXIS_IARG_81_WIDTH/8-1:0] ap_axis_iarg_81_tstrb,
    output [S_AXIS_IARG_81_WIDTH-1:0] ap_axis_iarg_81_tdata,
    //input AXI-Stream pass-through interface 82
    input s_axis_iarg_82_aclk,
    input s_axis_iarg_82_aresetn,
    input s_axis_iarg_82_tlast,
    input s_axis_iarg_82_tvalid,
    input [S_AXIS_IARG_82_DMWIDTH/8-1:0] s_axis_iarg_82_tkeep,
    input [S_AXIS_IARG_82_DMWIDTH/8-1:0] s_axis_iarg_82_tstrb,
    input [S_AXIS_IARG_82_DMWIDTH-1:0] s_axis_iarg_82_tdata,
    output s_axis_iarg_82_tready,
    input ap_axis_iarg_82_tready,
    output ap_axis_iarg_82_tlast,
    output ap_axis_iarg_82_tvalid,
    output [S_AXIS_IARG_82_WIDTH/8-1:0] ap_axis_iarg_82_tkeep,
    output [S_AXIS_IARG_82_WIDTH/8-1:0] ap_axis_iarg_82_tstrb,
    output [S_AXIS_IARG_82_WIDTH-1:0] ap_axis_iarg_82_tdata,
    //input AXI-Stream pass-through interface 83
    input s_axis_iarg_83_aclk,
    input s_axis_iarg_83_aresetn,
    input s_axis_iarg_83_tlast,
    input s_axis_iarg_83_tvalid,
    input [S_AXIS_IARG_83_DMWIDTH/8-1:0] s_axis_iarg_83_tkeep,
    input [S_AXIS_IARG_83_DMWIDTH/8-1:0] s_axis_iarg_83_tstrb,
    input [S_AXIS_IARG_83_DMWIDTH-1:0] s_axis_iarg_83_tdata,
    output s_axis_iarg_83_tready,
    input ap_axis_iarg_83_tready,
    output ap_axis_iarg_83_tlast,
    output ap_axis_iarg_83_tvalid,
    output [S_AXIS_IARG_83_WIDTH/8-1:0] ap_axis_iarg_83_tkeep,
    output [S_AXIS_IARG_83_WIDTH/8-1:0] ap_axis_iarg_83_tstrb,
    output [S_AXIS_IARG_83_WIDTH-1:0] ap_axis_iarg_83_tdata,
    //input AXI-Stream pass-through interface 84
    input s_axis_iarg_84_aclk,
    input s_axis_iarg_84_aresetn,
    input s_axis_iarg_84_tlast,
    input s_axis_iarg_84_tvalid,
    input [S_AXIS_IARG_84_DMWIDTH/8-1:0] s_axis_iarg_84_tkeep,
    input [S_AXIS_IARG_84_DMWIDTH/8-1:0] s_axis_iarg_84_tstrb,
    input [S_AXIS_IARG_84_DMWIDTH-1:0] s_axis_iarg_84_tdata,
    output s_axis_iarg_84_tready,
    input ap_axis_iarg_84_tready,
    output ap_axis_iarg_84_tlast,
    output ap_axis_iarg_84_tvalid,
    output [S_AXIS_IARG_84_WIDTH/8-1:0] ap_axis_iarg_84_tkeep,
    output [S_AXIS_IARG_84_WIDTH/8-1:0] ap_axis_iarg_84_tstrb,
    output [S_AXIS_IARG_84_WIDTH-1:0] ap_axis_iarg_84_tdata,
    //input AXI-Stream pass-through interface 85
    input s_axis_iarg_85_aclk,
    input s_axis_iarg_85_aresetn,
    input s_axis_iarg_85_tlast,
    input s_axis_iarg_85_tvalid,
    input [S_AXIS_IARG_85_DMWIDTH/8-1:0] s_axis_iarg_85_tkeep,
    input [S_AXIS_IARG_85_DMWIDTH/8-1:0] s_axis_iarg_85_tstrb,
    input [S_AXIS_IARG_85_DMWIDTH-1:0] s_axis_iarg_85_tdata,
    output s_axis_iarg_85_tready,
    input ap_axis_iarg_85_tready,
    output ap_axis_iarg_85_tlast,
    output ap_axis_iarg_85_tvalid,
    output [S_AXIS_IARG_85_WIDTH/8-1:0] ap_axis_iarg_85_tkeep,
    output [S_AXIS_IARG_85_WIDTH/8-1:0] ap_axis_iarg_85_tstrb,
    output [S_AXIS_IARG_85_WIDTH-1:0] ap_axis_iarg_85_tdata,
    //input AXI-Stream pass-through interface 86
    input s_axis_iarg_86_aclk,
    input s_axis_iarg_86_aresetn,
    input s_axis_iarg_86_tlast,
    input s_axis_iarg_86_tvalid,
    input [S_AXIS_IARG_86_DMWIDTH/8-1:0] s_axis_iarg_86_tkeep,
    input [S_AXIS_IARG_86_DMWIDTH/8-1:0] s_axis_iarg_86_tstrb,
    input [S_AXIS_IARG_86_DMWIDTH-1:0] s_axis_iarg_86_tdata,
    output s_axis_iarg_86_tready,
    input ap_axis_iarg_86_tready,
    output ap_axis_iarg_86_tlast,
    output ap_axis_iarg_86_tvalid,
    output [S_AXIS_IARG_86_WIDTH/8-1:0] ap_axis_iarg_86_tkeep,
    output [S_AXIS_IARG_86_WIDTH/8-1:0] ap_axis_iarg_86_tstrb,
    output [S_AXIS_IARG_86_WIDTH-1:0] ap_axis_iarg_86_tdata,
    //input AXI-Stream pass-through interface 87
    input s_axis_iarg_87_aclk,
    input s_axis_iarg_87_aresetn,
    input s_axis_iarg_87_tlast,
    input s_axis_iarg_87_tvalid,
    input [S_AXIS_IARG_87_DMWIDTH/8-1:0] s_axis_iarg_87_tkeep,
    input [S_AXIS_IARG_87_DMWIDTH/8-1:0] s_axis_iarg_87_tstrb,
    input [S_AXIS_IARG_87_DMWIDTH-1:0] s_axis_iarg_87_tdata,
    output s_axis_iarg_87_tready,
    input ap_axis_iarg_87_tready,
    output ap_axis_iarg_87_tlast,
    output ap_axis_iarg_87_tvalid,
    output [S_AXIS_IARG_87_WIDTH/8-1:0] ap_axis_iarg_87_tkeep,
    output [S_AXIS_IARG_87_WIDTH/8-1:0] ap_axis_iarg_87_tstrb,
    output [S_AXIS_IARG_87_WIDTH-1:0] ap_axis_iarg_87_tdata,
    //input AXI-Stream pass-through interface 88
    input s_axis_iarg_88_aclk,
    input s_axis_iarg_88_aresetn,
    input s_axis_iarg_88_tlast,
    input s_axis_iarg_88_tvalid,
    input [S_AXIS_IARG_88_DMWIDTH/8-1:0] s_axis_iarg_88_tkeep,
    input [S_AXIS_IARG_88_DMWIDTH/8-1:0] s_axis_iarg_88_tstrb,
    input [S_AXIS_IARG_88_DMWIDTH-1:0] s_axis_iarg_88_tdata,
    output s_axis_iarg_88_tready,
    input ap_axis_iarg_88_tready,
    output ap_axis_iarg_88_tlast,
    output ap_axis_iarg_88_tvalid,
    output [S_AXIS_IARG_88_WIDTH/8-1:0] ap_axis_iarg_88_tkeep,
    output [S_AXIS_IARG_88_WIDTH/8-1:0] ap_axis_iarg_88_tstrb,
    output [S_AXIS_IARG_88_WIDTH-1:0] ap_axis_iarg_88_tdata,
    //input AXI-Stream pass-through interface 89
    input s_axis_iarg_89_aclk,
    input s_axis_iarg_89_aresetn,
    input s_axis_iarg_89_tlast,
    input s_axis_iarg_89_tvalid,
    input [S_AXIS_IARG_89_DMWIDTH/8-1:0] s_axis_iarg_89_tkeep,
    input [S_AXIS_IARG_89_DMWIDTH/8-1:0] s_axis_iarg_89_tstrb,
    input [S_AXIS_IARG_89_DMWIDTH-1:0] s_axis_iarg_89_tdata,
    output s_axis_iarg_89_tready,
    input ap_axis_iarg_89_tready,
    output ap_axis_iarg_89_tlast,
    output ap_axis_iarg_89_tvalid,
    output [S_AXIS_IARG_89_WIDTH/8-1:0] ap_axis_iarg_89_tkeep,
    output [S_AXIS_IARG_89_WIDTH/8-1:0] ap_axis_iarg_89_tstrb,
    output [S_AXIS_IARG_89_WIDTH-1:0] ap_axis_iarg_89_tdata,
    //input AXI-Stream pass-through interface 90
    input s_axis_iarg_90_aclk,
    input s_axis_iarg_90_aresetn,
    input s_axis_iarg_90_tlast,
    input s_axis_iarg_90_tvalid,
    input [S_AXIS_IARG_90_DMWIDTH/8-1:0] s_axis_iarg_90_tkeep,
    input [S_AXIS_IARG_90_DMWIDTH/8-1:0] s_axis_iarg_90_tstrb,
    input [S_AXIS_IARG_90_DMWIDTH-1:0] s_axis_iarg_90_tdata,
    output s_axis_iarg_90_tready,
    input ap_axis_iarg_90_tready,
    output ap_axis_iarg_90_tlast,
    output ap_axis_iarg_90_tvalid,
    output [S_AXIS_IARG_90_WIDTH/8-1:0] ap_axis_iarg_90_tkeep,
    output [S_AXIS_IARG_90_WIDTH/8-1:0] ap_axis_iarg_90_tstrb,
    output [S_AXIS_IARG_90_WIDTH-1:0] ap_axis_iarg_90_tdata,
    //input AXI-Stream pass-through interface 91
    input s_axis_iarg_91_aclk,
    input s_axis_iarg_91_aresetn,
    input s_axis_iarg_91_tlast,
    input s_axis_iarg_91_tvalid,
    input [S_AXIS_IARG_91_DMWIDTH/8-1:0] s_axis_iarg_91_tkeep,
    input [S_AXIS_IARG_91_DMWIDTH/8-1:0] s_axis_iarg_91_tstrb,
    input [S_AXIS_IARG_91_DMWIDTH-1:0] s_axis_iarg_91_tdata,
    output s_axis_iarg_91_tready,
    input ap_axis_iarg_91_tready,
    output ap_axis_iarg_91_tlast,
    output ap_axis_iarg_91_tvalid,
    output [S_AXIS_IARG_91_WIDTH/8-1:0] ap_axis_iarg_91_tkeep,
    output [S_AXIS_IARG_91_WIDTH/8-1:0] ap_axis_iarg_91_tstrb,
    output [S_AXIS_IARG_91_WIDTH-1:0] ap_axis_iarg_91_tdata,
    //input AXI-Stream pass-through interface 92
    input s_axis_iarg_92_aclk,
    input s_axis_iarg_92_aresetn,
    input s_axis_iarg_92_tlast,
    input s_axis_iarg_92_tvalid,
    input [S_AXIS_IARG_92_DMWIDTH/8-1:0] s_axis_iarg_92_tkeep,
    input [S_AXIS_IARG_92_DMWIDTH/8-1:0] s_axis_iarg_92_tstrb,
    input [S_AXIS_IARG_92_DMWIDTH-1:0] s_axis_iarg_92_tdata,
    output s_axis_iarg_92_tready,
    input ap_axis_iarg_92_tready,
    output ap_axis_iarg_92_tlast,
    output ap_axis_iarg_92_tvalid,
    output [S_AXIS_IARG_92_WIDTH/8-1:0] ap_axis_iarg_92_tkeep,
    output [S_AXIS_IARG_92_WIDTH/8-1:0] ap_axis_iarg_92_tstrb,
    output [S_AXIS_IARG_92_WIDTH-1:0] ap_axis_iarg_92_tdata,
    //input AXI-Stream pass-through interface 93
    input s_axis_iarg_93_aclk,
    input s_axis_iarg_93_aresetn,
    input s_axis_iarg_93_tlast,
    input s_axis_iarg_93_tvalid,
    input [S_AXIS_IARG_93_DMWIDTH/8-1:0] s_axis_iarg_93_tkeep,
    input [S_AXIS_IARG_93_DMWIDTH/8-1:0] s_axis_iarg_93_tstrb,
    input [S_AXIS_IARG_93_DMWIDTH-1:0] s_axis_iarg_93_tdata,
    output s_axis_iarg_93_tready,
    input ap_axis_iarg_93_tready,
    output ap_axis_iarg_93_tlast,
    output ap_axis_iarg_93_tvalid,
    output [S_AXIS_IARG_93_WIDTH/8-1:0] ap_axis_iarg_93_tkeep,
    output [S_AXIS_IARG_93_WIDTH/8-1:0] ap_axis_iarg_93_tstrb,
    output [S_AXIS_IARG_93_WIDTH-1:0] ap_axis_iarg_93_tdata,
    //input AXI-Stream pass-through interface 94
    input s_axis_iarg_94_aclk,
    input s_axis_iarg_94_aresetn,
    input s_axis_iarg_94_tlast,
    input s_axis_iarg_94_tvalid,
    input [S_AXIS_IARG_94_DMWIDTH/8-1:0] s_axis_iarg_94_tkeep,
    input [S_AXIS_IARG_94_DMWIDTH/8-1:0] s_axis_iarg_94_tstrb,
    input [S_AXIS_IARG_94_DMWIDTH-1:0] s_axis_iarg_94_tdata,
    output s_axis_iarg_94_tready,
    input ap_axis_iarg_94_tready,
    output ap_axis_iarg_94_tlast,
    output ap_axis_iarg_94_tvalid,
    output [S_AXIS_IARG_94_WIDTH/8-1:0] ap_axis_iarg_94_tkeep,
    output [S_AXIS_IARG_94_WIDTH/8-1:0] ap_axis_iarg_94_tstrb,
    output [S_AXIS_IARG_94_WIDTH-1:0] ap_axis_iarg_94_tdata,
    //input AXI-Stream pass-through interface 95
    input s_axis_iarg_95_aclk,
    input s_axis_iarg_95_aresetn,
    input s_axis_iarg_95_tlast,
    input s_axis_iarg_95_tvalid,
    input [S_AXIS_IARG_95_DMWIDTH/8-1:0] s_axis_iarg_95_tkeep,
    input [S_AXIS_IARG_95_DMWIDTH/8-1:0] s_axis_iarg_95_tstrb,
    input [S_AXIS_IARG_95_DMWIDTH-1:0] s_axis_iarg_95_tdata,
    output s_axis_iarg_95_tready,
    input ap_axis_iarg_95_tready,
    output ap_axis_iarg_95_tlast,
    output ap_axis_iarg_95_tvalid,
    output [S_AXIS_IARG_95_WIDTH/8-1:0] ap_axis_iarg_95_tkeep,
    output [S_AXIS_IARG_95_WIDTH/8-1:0] ap_axis_iarg_95_tstrb,
    output [S_AXIS_IARG_95_WIDTH-1:0] ap_axis_iarg_95_tdata,
    //input AXI-Stream pass-through interface 96
    input s_axis_iarg_96_aclk,
    input s_axis_iarg_96_aresetn,
    input s_axis_iarg_96_tlast,
    input s_axis_iarg_96_tvalid,
    input [S_AXIS_IARG_96_DMWIDTH/8-1:0] s_axis_iarg_96_tkeep,
    input [S_AXIS_IARG_96_DMWIDTH/8-1:0] s_axis_iarg_96_tstrb,
    input [S_AXIS_IARG_96_DMWIDTH-1:0] s_axis_iarg_96_tdata,
    output s_axis_iarg_96_tready,
    input ap_axis_iarg_96_tready,
    output ap_axis_iarg_96_tlast,
    output ap_axis_iarg_96_tvalid,
    output [S_AXIS_IARG_96_WIDTH/8-1:0] ap_axis_iarg_96_tkeep,
    output [S_AXIS_IARG_96_WIDTH/8-1:0] ap_axis_iarg_96_tstrb,
    output [S_AXIS_IARG_96_WIDTH-1:0] ap_axis_iarg_96_tdata,
    //input AXI-Stream pass-through interface 97
    input s_axis_iarg_97_aclk,
    input s_axis_iarg_97_aresetn,
    input s_axis_iarg_97_tlast,
    input s_axis_iarg_97_tvalid,
    input [S_AXIS_IARG_97_DMWIDTH/8-1:0] s_axis_iarg_97_tkeep,
    input [S_AXIS_IARG_97_DMWIDTH/8-1:0] s_axis_iarg_97_tstrb,
    input [S_AXIS_IARG_97_DMWIDTH-1:0] s_axis_iarg_97_tdata,
    output s_axis_iarg_97_tready,
    input ap_axis_iarg_97_tready,
    output ap_axis_iarg_97_tlast,
    output ap_axis_iarg_97_tvalid,
    output [S_AXIS_IARG_97_WIDTH/8-1:0] ap_axis_iarg_97_tkeep,
    output [S_AXIS_IARG_97_WIDTH/8-1:0] ap_axis_iarg_97_tstrb,
    output [S_AXIS_IARG_97_WIDTH-1:0] ap_axis_iarg_97_tdata,
    //input AXI-Stream pass-through interface 98
    input s_axis_iarg_98_aclk,
    input s_axis_iarg_98_aresetn,
    input s_axis_iarg_98_tlast,
    input s_axis_iarg_98_tvalid,
    input [S_AXIS_IARG_98_DMWIDTH/8-1:0] s_axis_iarg_98_tkeep,
    input [S_AXIS_IARG_98_DMWIDTH/8-1:0] s_axis_iarg_98_tstrb,
    input [S_AXIS_IARG_98_DMWIDTH-1:0] s_axis_iarg_98_tdata,
    output s_axis_iarg_98_tready,
    input ap_axis_iarg_98_tready,
    output ap_axis_iarg_98_tlast,
    output ap_axis_iarg_98_tvalid,
    output [S_AXIS_IARG_98_WIDTH/8-1:0] ap_axis_iarg_98_tkeep,
    output [S_AXIS_IARG_98_WIDTH/8-1:0] ap_axis_iarg_98_tstrb,
    output [S_AXIS_IARG_98_WIDTH-1:0] ap_axis_iarg_98_tdata,
    //input AXI-Stream pass-through interface 99
    input s_axis_iarg_99_aclk,
    input s_axis_iarg_99_aresetn,
    input s_axis_iarg_99_tlast,
    input s_axis_iarg_99_tvalid,
    input [S_AXIS_IARG_99_DMWIDTH/8-1:0] s_axis_iarg_99_tkeep,
    input [S_AXIS_IARG_99_DMWIDTH/8-1:0] s_axis_iarg_99_tstrb,
    input [S_AXIS_IARG_99_DMWIDTH-1:0] s_axis_iarg_99_tdata,
    output s_axis_iarg_99_tready,
    input ap_axis_iarg_99_tready,
    output ap_axis_iarg_99_tlast,
    output ap_axis_iarg_99_tvalid,
    output [S_AXIS_IARG_99_WIDTH/8-1:0] ap_axis_iarg_99_tkeep,
    output [S_AXIS_IARG_99_WIDTH/8-1:0] ap_axis_iarg_99_tstrb,
    output [S_AXIS_IARG_99_WIDTH-1:0] ap_axis_iarg_99_tdata,
    //input AXI-Stream pass-through interface 100
    input s_axis_iarg_100_aclk,
    input s_axis_iarg_100_aresetn,
    input s_axis_iarg_100_tlast,
    input s_axis_iarg_100_tvalid,
    input [S_AXIS_IARG_100_DMWIDTH/8-1:0] s_axis_iarg_100_tkeep,
    input [S_AXIS_IARG_100_DMWIDTH/8-1:0] s_axis_iarg_100_tstrb,
    input [S_AXIS_IARG_100_DMWIDTH-1:0] s_axis_iarg_100_tdata,
    output s_axis_iarg_100_tready,
    input ap_axis_iarg_100_tready,
    output ap_axis_iarg_100_tlast,
    output ap_axis_iarg_100_tvalid,
    output [S_AXIS_IARG_100_WIDTH/8-1:0] ap_axis_iarg_100_tkeep,
    output [S_AXIS_IARG_100_WIDTH/8-1:0] ap_axis_iarg_100_tstrb,
    output [S_AXIS_IARG_100_WIDTH-1:0] ap_axis_iarg_100_tdata,
    //input AXI-Stream pass-through interface 101
    input s_axis_iarg_101_aclk,
    input s_axis_iarg_101_aresetn,
    input s_axis_iarg_101_tlast,
    input s_axis_iarg_101_tvalid,
    input [S_AXIS_IARG_101_DMWIDTH/8-1:0] s_axis_iarg_101_tkeep,
    input [S_AXIS_IARG_101_DMWIDTH/8-1:0] s_axis_iarg_101_tstrb,
    input [S_AXIS_IARG_101_DMWIDTH-1:0] s_axis_iarg_101_tdata,
    output s_axis_iarg_101_tready,
    input ap_axis_iarg_101_tready,
    output ap_axis_iarg_101_tlast,
    output ap_axis_iarg_101_tvalid,
    output [S_AXIS_IARG_101_WIDTH/8-1:0] ap_axis_iarg_101_tkeep,
    output [S_AXIS_IARG_101_WIDTH/8-1:0] ap_axis_iarg_101_tstrb,
    output [S_AXIS_IARG_101_WIDTH-1:0] ap_axis_iarg_101_tdata,
    //input AXI-Stream pass-through interface 102
    input s_axis_iarg_102_aclk,
    input s_axis_iarg_102_aresetn,
    input s_axis_iarg_102_tlast,
    input s_axis_iarg_102_tvalid,
    input [S_AXIS_IARG_102_DMWIDTH/8-1:0] s_axis_iarg_102_tkeep,
    input [S_AXIS_IARG_102_DMWIDTH/8-1:0] s_axis_iarg_102_tstrb,
    input [S_AXIS_IARG_102_DMWIDTH-1:0] s_axis_iarg_102_tdata,
    output s_axis_iarg_102_tready,
    input ap_axis_iarg_102_tready,
    output ap_axis_iarg_102_tlast,
    output ap_axis_iarg_102_tvalid,
    output [S_AXIS_IARG_102_WIDTH/8-1:0] ap_axis_iarg_102_tkeep,
    output [S_AXIS_IARG_102_WIDTH/8-1:0] ap_axis_iarg_102_tstrb,
    output [S_AXIS_IARG_102_WIDTH-1:0] ap_axis_iarg_102_tdata,
    //input AXI-Stream pass-through interface 103
    input s_axis_iarg_103_aclk,
    input s_axis_iarg_103_aresetn,
    input s_axis_iarg_103_tlast,
    input s_axis_iarg_103_tvalid,
    input [S_AXIS_IARG_103_DMWIDTH/8-1:0] s_axis_iarg_103_tkeep,
    input [S_AXIS_IARG_103_DMWIDTH/8-1:0] s_axis_iarg_103_tstrb,
    input [S_AXIS_IARG_103_DMWIDTH-1:0] s_axis_iarg_103_tdata,
    output s_axis_iarg_103_tready,
    input ap_axis_iarg_103_tready,
    output ap_axis_iarg_103_tlast,
    output ap_axis_iarg_103_tvalid,
    output [S_AXIS_IARG_103_WIDTH/8-1:0] ap_axis_iarg_103_tkeep,
    output [S_AXIS_IARG_103_WIDTH/8-1:0] ap_axis_iarg_103_tstrb,
    output [S_AXIS_IARG_103_WIDTH-1:0] ap_axis_iarg_103_tdata,
    //input AXI-Stream pass-through interface 104
    input s_axis_iarg_104_aclk,
    input s_axis_iarg_104_aresetn,
    input s_axis_iarg_104_tlast,
    input s_axis_iarg_104_tvalid,
    input [S_AXIS_IARG_104_DMWIDTH/8-1:0] s_axis_iarg_104_tkeep,
    input [S_AXIS_IARG_104_DMWIDTH/8-1:0] s_axis_iarg_104_tstrb,
    input [S_AXIS_IARG_104_DMWIDTH-1:0] s_axis_iarg_104_tdata,
    output s_axis_iarg_104_tready,
    input ap_axis_iarg_104_tready,
    output ap_axis_iarg_104_tlast,
    output ap_axis_iarg_104_tvalid,
    output [S_AXIS_IARG_104_WIDTH/8-1:0] ap_axis_iarg_104_tkeep,
    output [S_AXIS_IARG_104_WIDTH/8-1:0] ap_axis_iarg_104_tstrb,
    output [S_AXIS_IARG_104_WIDTH-1:0] ap_axis_iarg_104_tdata,
    //input AXI-Stream pass-through interface 105
    input s_axis_iarg_105_aclk,
    input s_axis_iarg_105_aresetn,
    input s_axis_iarg_105_tlast,
    input s_axis_iarg_105_tvalid,
    input [S_AXIS_IARG_105_DMWIDTH/8-1:0] s_axis_iarg_105_tkeep,
    input [S_AXIS_IARG_105_DMWIDTH/8-1:0] s_axis_iarg_105_tstrb,
    input [S_AXIS_IARG_105_DMWIDTH-1:0] s_axis_iarg_105_tdata,
    output s_axis_iarg_105_tready,
    input ap_axis_iarg_105_tready,
    output ap_axis_iarg_105_tlast,
    output ap_axis_iarg_105_tvalid,
    output [S_AXIS_IARG_105_WIDTH/8-1:0] ap_axis_iarg_105_tkeep,
    output [S_AXIS_IARG_105_WIDTH/8-1:0] ap_axis_iarg_105_tstrb,
    output [S_AXIS_IARG_105_WIDTH-1:0] ap_axis_iarg_105_tdata,
    //input AXI-Stream pass-through interface 106
    input s_axis_iarg_106_aclk,
    input s_axis_iarg_106_aresetn,
    input s_axis_iarg_106_tlast,
    input s_axis_iarg_106_tvalid,
    input [S_AXIS_IARG_106_DMWIDTH/8-1:0] s_axis_iarg_106_tkeep,
    input [S_AXIS_IARG_106_DMWIDTH/8-1:0] s_axis_iarg_106_tstrb,
    input [S_AXIS_IARG_106_DMWIDTH-1:0] s_axis_iarg_106_tdata,
    output s_axis_iarg_106_tready,
    input ap_axis_iarg_106_tready,
    output ap_axis_iarg_106_tlast,
    output ap_axis_iarg_106_tvalid,
    output [S_AXIS_IARG_106_WIDTH/8-1:0] ap_axis_iarg_106_tkeep,
    output [S_AXIS_IARG_106_WIDTH/8-1:0] ap_axis_iarg_106_tstrb,
    output [S_AXIS_IARG_106_WIDTH-1:0] ap_axis_iarg_106_tdata,
    //input AXI-Stream pass-through interface 107
    input s_axis_iarg_107_aclk,
    input s_axis_iarg_107_aresetn,
    input s_axis_iarg_107_tlast,
    input s_axis_iarg_107_tvalid,
    input [S_AXIS_IARG_107_DMWIDTH/8-1:0] s_axis_iarg_107_tkeep,
    input [S_AXIS_IARG_107_DMWIDTH/8-1:0] s_axis_iarg_107_tstrb,
    input [S_AXIS_IARG_107_DMWIDTH-1:0] s_axis_iarg_107_tdata,
    output s_axis_iarg_107_tready,
    input ap_axis_iarg_107_tready,
    output ap_axis_iarg_107_tlast,
    output ap_axis_iarg_107_tvalid,
    output [S_AXIS_IARG_107_WIDTH/8-1:0] ap_axis_iarg_107_tkeep,
    output [S_AXIS_IARG_107_WIDTH/8-1:0] ap_axis_iarg_107_tstrb,
    output [S_AXIS_IARG_107_WIDTH-1:0] ap_axis_iarg_107_tdata,
    //input AXI-Stream pass-through interface 108
    input s_axis_iarg_108_aclk,
    input s_axis_iarg_108_aresetn,
    input s_axis_iarg_108_tlast,
    input s_axis_iarg_108_tvalid,
    input [S_AXIS_IARG_108_DMWIDTH/8-1:0] s_axis_iarg_108_tkeep,
    input [S_AXIS_IARG_108_DMWIDTH/8-1:0] s_axis_iarg_108_tstrb,
    input [S_AXIS_IARG_108_DMWIDTH-1:0] s_axis_iarg_108_tdata,
    output s_axis_iarg_108_tready,
    input ap_axis_iarg_108_tready,
    output ap_axis_iarg_108_tlast,
    output ap_axis_iarg_108_tvalid,
    output [S_AXIS_IARG_108_WIDTH/8-1:0] ap_axis_iarg_108_tkeep,
    output [S_AXIS_IARG_108_WIDTH/8-1:0] ap_axis_iarg_108_tstrb,
    output [S_AXIS_IARG_108_WIDTH-1:0] ap_axis_iarg_108_tdata,
    //input AXI-Stream pass-through interface 109
    input s_axis_iarg_109_aclk,
    input s_axis_iarg_109_aresetn,
    input s_axis_iarg_109_tlast,
    input s_axis_iarg_109_tvalid,
    input [S_AXIS_IARG_109_DMWIDTH/8-1:0] s_axis_iarg_109_tkeep,
    input [S_AXIS_IARG_109_DMWIDTH/8-1:0] s_axis_iarg_109_tstrb,
    input [S_AXIS_IARG_109_DMWIDTH-1:0] s_axis_iarg_109_tdata,
    output s_axis_iarg_109_tready,
    input ap_axis_iarg_109_tready,
    output ap_axis_iarg_109_tlast,
    output ap_axis_iarg_109_tvalid,
    output [S_AXIS_IARG_109_WIDTH/8-1:0] ap_axis_iarg_109_tkeep,
    output [S_AXIS_IARG_109_WIDTH/8-1:0] ap_axis_iarg_109_tstrb,
    output [S_AXIS_IARG_109_WIDTH-1:0] ap_axis_iarg_109_tdata,
    //input AXI-Stream pass-through interface 110
    input s_axis_iarg_110_aclk,
    input s_axis_iarg_110_aresetn,
    input s_axis_iarg_110_tlast,
    input s_axis_iarg_110_tvalid,
    input [S_AXIS_IARG_110_DMWIDTH/8-1:0] s_axis_iarg_110_tkeep,
    input [S_AXIS_IARG_110_DMWIDTH/8-1:0] s_axis_iarg_110_tstrb,
    input [S_AXIS_IARG_110_DMWIDTH-1:0] s_axis_iarg_110_tdata,
    output s_axis_iarg_110_tready,
    input ap_axis_iarg_110_tready,
    output ap_axis_iarg_110_tlast,
    output ap_axis_iarg_110_tvalid,
    output [S_AXIS_IARG_110_WIDTH/8-1:0] ap_axis_iarg_110_tkeep,
    output [S_AXIS_IARG_110_WIDTH/8-1:0] ap_axis_iarg_110_tstrb,
    output [S_AXIS_IARG_110_WIDTH-1:0] ap_axis_iarg_110_tdata,
    //input AXI-Stream pass-through interface 111
    input s_axis_iarg_111_aclk,
    input s_axis_iarg_111_aresetn,
    input s_axis_iarg_111_tlast,
    input s_axis_iarg_111_tvalid,
    input [S_AXIS_IARG_111_DMWIDTH/8-1:0] s_axis_iarg_111_tkeep,
    input [S_AXIS_IARG_111_DMWIDTH/8-1:0] s_axis_iarg_111_tstrb,
    input [S_AXIS_IARG_111_DMWIDTH-1:0] s_axis_iarg_111_tdata,
    output s_axis_iarg_111_tready,
    input ap_axis_iarg_111_tready,
    output ap_axis_iarg_111_tlast,
    output ap_axis_iarg_111_tvalid,
    output [S_AXIS_IARG_111_WIDTH/8-1:0] ap_axis_iarg_111_tkeep,
    output [S_AXIS_IARG_111_WIDTH/8-1:0] ap_axis_iarg_111_tstrb,
    output [S_AXIS_IARG_111_WIDTH-1:0] ap_axis_iarg_111_tdata,
    //input AXI-Stream pass-through interface 112
    input s_axis_iarg_112_aclk,
    input s_axis_iarg_112_aresetn,
    input s_axis_iarg_112_tlast,
    input s_axis_iarg_112_tvalid,
    input [S_AXIS_IARG_112_DMWIDTH/8-1:0] s_axis_iarg_112_tkeep,
    input [S_AXIS_IARG_112_DMWIDTH/8-1:0] s_axis_iarg_112_tstrb,
    input [S_AXIS_IARG_112_DMWIDTH-1:0] s_axis_iarg_112_tdata,
    output s_axis_iarg_112_tready,
    input ap_axis_iarg_112_tready,
    output ap_axis_iarg_112_tlast,
    output ap_axis_iarg_112_tvalid,
    output [S_AXIS_IARG_112_WIDTH/8-1:0] ap_axis_iarg_112_tkeep,
    output [S_AXIS_IARG_112_WIDTH/8-1:0] ap_axis_iarg_112_tstrb,
    output [S_AXIS_IARG_112_WIDTH-1:0] ap_axis_iarg_112_tdata,
    //input AXI-Stream pass-through interface 113
    input s_axis_iarg_113_aclk,
    input s_axis_iarg_113_aresetn,
    input s_axis_iarg_113_tlast,
    input s_axis_iarg_113_tvalid,
    input [S_AXIS_IARG_113_DMWIDTH/8-1:0] s_axis_iarg_113_tkeep,
    input [S_AXIS_IARG_113_DMWIDTH/8-1:0] s_axis_iarg_113_tstrb,
    input [S_AXIS_IARG_113_DMWIDTH-1:0] s_axis_iarg_113_tdata,
    output s_axis_iarg_113_tready,
    input ap_axis_iarg_113_tready,
    output ap_axis_iarg_113_tlast,
    output ap_axis_iarg_113_tvalid,
    output [S_AXIS_IARG_113_WIDTH/8-1:0] ap_axis_iarg_113_tkeep,
    output [S_AXIS_IARG_113_WIDTH/8-1:0] ap_axis_iarg_113_tstrb,
    output [S_AXIS_IARG_113_WIDTH-1:0] ap_axis_iarg_113_tdata,
    //input AXI-Stream pass-through interface 114
    input s_axis_iarg_114_aclk,
    input s_axis_iarg_114_aresetn,
    input s_axis_iarg_114_tlast,
    input s_axis_iarg_114_tvalid,
    input [S_AXIS_IARG_114_DMWIDTH/8-1:0] s_axis_iarg_114_tkeep,
    input [S_AXIS_IARG_114_DMWIDTH/8-1:0] s_axis_iarg_114_tstrb,
    input [S_AXIS_IARG_114_DMWIDTH-1:0] s_axis_iarg_114_tdata,
    output s_axis_iarg_114_tready,
    input ap_axis_iarg_114_tready,
    output ap_axis_iarg_114_tlast,
    output ap_axis_iarg_114_tvalid,
    output [S_AXIS_IARG_114_WIDTH/8-1:0] ap_axis_iarg_114_tkeep,
    output [S_AXIS_IARG_114_WIDTH/8-1:0] ap_axis_iarg_114_tstrb,
    output [S_AXIS_IARG_114_WIDTH-1:0] ap_axis_iarg_114_tdata,
    //input AXI-Stream pass-through interface 115
    input s_axis_iarg_115_aclk,
    input s_axis_iarg_115_aresetn,
    input s_axis_iarg_115_tlast,
    input s_axis_iarg_115_tvalid,
    input [S_AXIS_IARG_115_DMWIDTH/8-1:0] s_axis_iarg_115_tkeep,
    input [S_AXIS_IARG_115_DMWIDTH/8-1:0] s_axis_iarg_115_tstrb,
    input [S_AXIS_IARG_115_DMWIDTH-1:0] s_axis_iarg_115_tdata,
    output s_axis_iarg_115_tready,
    input ap_axis_iarg_115_tready,
    output ap_axis_iarg_115_tlast,
    output ap_axis_iarg_115_tvalid,
    output [S_AXIS_IARG_115_WIDTH/8-1:0] ap_axis_iarg_115_tkeep,
    output [S_AXIS_IARG_115_WIDTH/8-1:0] ap_axis_iarg_115_tstrb,
    output [S_AXIS_IARG_115_WIDTH-1:0] ap_axis_iarg_115_tdata,
    //input AXI-Stream pass-through interface 116
    input s_axis_iarg_116_aclk,
    input s_axis_iarg_116_aresetn,
    input s_axis_iarg_116_tlast,
    input s_axis_iarg_116_tvalid,
    input [S_AXIS_IARG_116_DMWIDTH/8-1:0] s_axis_iarg_116_tkeep,
    input [S_AXIS_IARG_116_DMWIDTH/8-1:0] s_axis_iarg_116_tstrb,
    input [S_AXIS_IARG_116_DMWIDTH-1:0] s_axis_iarg_116_tdata,
    output s_axis_iarg_116_tready,
    input ap_axis_iarg_116_tready,
    output ap_axis_iarg_116_tlast,
    output ap_axis_iarg_116_tvalid,
    output [S_AXIS_IARG_116_WIDTH/8-1:0] ap_axis_iarg_116_tkeep,
    output [S_AXIS_IARG_116_WIDTH/8-1:0] ap_axis_iarg_116_tstrb,
    output [S_AXIS_IARG_116_WIDTH-1:0] ap_axis_iarg_116_tdata,
    //input AXI-Stream pass-through interface 117
    input s_axis_iarg_117_aclk,
    input s_axis_iarg_117_aresetn,
    input s_axis_iarg_117_tlast,
    input s_axis_iarg_117_tvalid,
    input [S_AXIS_IARG_117_DMWIDTH/8-1:0] s_axis_iarg_117_tkeep,
    input [S_AXIS_IARG_117_DMWIDTH/8-1:0] s_axis_iarg_117_tstrb,
    input [S_AXIS_IARG_117_DMWIDTH-1:0] s_axis_iarg_117_tdata,
    output s_axis_iarg_117_tready,
    input ap_axis_iarg_117_tready,
    output ap_axis_iarg_117_tlast,
    output ap_axis_iarg_117_tvalid,
    output [S_AXIS_IARG_117_WIDTH/8-1:0] ap_axis_iarg_117_tkeep,
    output [S_AXIS_IARG_117_WIDTH/8-1:0] ap_axis_iarg_117_tstrb,
    output [S_AXIS_IARG_117_WIDTH-1:0] ap_axis_iarg_117_tdata,
    //input AXI-Stream pass-through interface 118
    input s_axis_iarg_118_aclk,
    input s_axis_iarg_118_aresetn,
    input s_axis_iarg_118_tlast,
    input s_axis_iarg_118_tvalid,
    input [S_AXIS_IARG_118_DMWIDTH/8-1:0] s_axis_iarg_118_tkeep,
    input [S_AXIS_IARG_118_DMWIDTH/8-1:0] s_axis_iarg_118_tstrb,
    input [S_AXIS_IARG_118_DMWIDTH-1:0] s_axis_iarg_118_tdata,
    output s_axis_iarg_118_tready,
    input ap_axis_iarg_118_tready,
    output ap_axis_iarg_118_tlast,
    output ap_axis_iarg_118_tvalid,
    output [S_AXIS_IARG_118_WIDTH/8-1:0] ap_axis_iarg_118_tkeep,
    output [S_AXIS_IARG_118_WIDTH/8-1:0] ap_axis_iarg_118_tstrb,
    output [S_AXIS_IARG_118_WIDTH-1:0] ap_axis_iarg_118_tdata,
    //input AXI-Stream pass-through interface 119
    input s_axis_iarg_119_aclk,
    input s_axis_iarg_119_aresetn,
    input s_axis_iarg_119_tlast,
    input s_axis_iarg_119_tvalid,
    input [S_AXIS_IARG_119_DMWIDTH/8-1:0] s_axis_iarg_119_tkeep,
    input [S_AXIS_IARG_119_DMWIDTH/8-1:0] s_axis_iarg_119_tstrb,
    input [S_AXIS_IARG_119_DMWIDTH-1:0] s_axis_iarg_119_tdata,
    output s_axis_iarg_119_tready,
    input ap_axis_iarg_119_tready,
    output ap_axis_iarg_119_tlast,
    output ap_axis_iarg_119_tvalid,
    output [S_AXIS_IARG_119_WIDTH/8-1:0] ap_axis_iarg_119_tkeep,
    output [S_AXIS_IARG_119_WIDTH/8-1:0] ap_axis_iarg_119_tstrb,
    output [S_AXIS_IARG_119_WIDTH-1:0] ap_axis_iarg_119_tdata,
    //input AXI-Stream pass-through interface 120
    input s_axis_iarg_120_aclk,
    input s_axis_iarg_120_aresetn,
    input s_axis_iarg_120_tlast,
    input s_axis_iarg_120_tvalid,
    input [S_AXIS_IARG_120_DMWIDTH/8-1:0] s_axis_iarg_120_tkeep,
    input [S_AXIS_IARG_120_DMWIDTH/8-1:0] s_axis_iarg_120_tstrb,
    input [S_AXIS_IARG_120_DMWIDTH-1:0] s_axis_iarg_120_tdata,
    output s_axis_iarg_120_tready,
    input ap_axis_iarg_120_tready,
    output ap_axis_iarg_120_tlast,
    output ap_axis_iarg_120_tvalid,
    output [S_AXIS_IARG_120_WIDTH/8-1:0] ap_axis_iarg_120_tkeep,
    output [S_AXIS_IARG_120_WIDTH/8-1:0] ap_axis_iarg_120_tstrb,
    output [S_AXIS_IARG_120_WIDTH-1:0] ap_axis_iarg_120_tdata,
    //input AXI-Stream pass-through interface 121
    input s_axis_iarg_121_aclk,
    input s_axis_iarg_121_aresetn,
    input s_axis_iarg_121_tlast,
    input s_axis_iarg_121_tvalid,
    input [S_AXIS_IARG_121_DMWIDTH/8-1:0] s_axis_iarg_121_tkeep,
    input [S_AXIS_IARG_121_DMWIDTH/8-1:0] s_axis_iarg_121_tstrb,
    input [S_AXIS_IARG_121_DMWIDTH-1:0] s_axis_iarg_121_tdata,
    output s_axis_iarg_121_tready,
    input ap_axis_iarg_121_tready,
    output ap_axis_iarg_121_tlast,
    output ap_axis_iarg_121_tvalid,
    output [S_AXIS_IARG_121_WIDTH/8-1:0] ap_axis_iarg_121_tkeep,
    output [S_AXIS_IARG_121_WIDTH/8-1:0] ap_axis_iarg_121_tstrb,
    output [S_AXIS_IARG_121_WIDTH-1:0] ap_axis_iarg_121_tdata,
    //input AXI-Stream pass-through interface 122
    input s_axis_iarg_122_aclk,
    input s_axis_iarg_122_aresetn,
    input s_axis_iarg_122_tlast,
    input s_axis_iarg_122_tvalid,
    input [S_AXIS_IARG_122_DMWIDTH/8-1:0] s_axis_iarg_122_tkeep,
    input [S_AXIS_IARG_122_DMWIDTH/8-1:0] s_axis_iarg_122_tstrb,
    input [S_AXIS_IARG_122_DMWIDTH-1:0] s_axis_iarg_122_tdata,
    output s_axis_iarg_122_tready,
    input ap_axis_iarg_122_tready,
    output ap_axis_iarg_122_tlast,
    output ap_axis_iarg_122_tvalid,
    output [S_AXIS_IARG_122_WIDTH/8-1:0] ap_axis_iarg_122_tkeep,
    output [S_AXIS_IARG_122_WIDTH/8-1:0] ap_axis_iarg_122_tstrb,
    output [S_AXIS_IARG_122_WIDTH-1:0] ap_axis_iarg_122_tdata,
    //input AXI-Stream pass-through interface 123
    input s_axis_iarg_123_aclk,
    input s_axis_iarg_123_aresetn,
    input s_axis_iarg_123_tlast,
    input s_axis_iarg_123_tvalid,
    input [S_AXIS_IARG_123_DMWIDTH/8-1:0] s_axis_iarg_123_tkeep,
    input [S_AXIS_IARG_123_DMWIDTH/8-1:0] s_axis_iarg_123_tstrb,
    input [S_AXIS_IARG_123_DMWIDTH-1:0] s_axis_iarg_123_tdata,
    output s_axis_iarg_123_tready,
    input ap_axis_iarg_123_tready,
    output ap_axis_iarg_123_tlast,
    output ap_axis_iarg_123_tvalid,
    output [S_AXIS_IARG_123_WIDTH/8-1:0] ap_axis_iarg_123_tkeep,
    output [S_AXIS_IARG_123_WIDTH/8-1:0] ap_axis_iarg_123_tstrb,
    output [S_AXIS_IARG_123_WIDTH-1:0] ap_axis_iarg_123_tdata,
    //input AXI-Stream pass-through interface 124
    input s_axis_iarg_124_aclk,
    input s_axis_iarg_124_aresetn,
    input s_axis_iarg_124_tlast,
    input s_axis_iarg_124_tvalid,
    input [S_AXIS_IARG_124_DMWIDTH/8-1:0] s_axis_iarg_124_tkeep,
    input [S_AXIS_IARG_124_DMWIDTH/8-1:0] s_axis_iarg_124_tstrb,
    input [S_AXIS_IARG_124_DMWIDTH-1:0] s_axis_iarg_124_tdata,
    output s_axis_iarg_124_tready,
    input ap_axis_iarg_124_tready,
    output ap_axis_iarg_124_tlast,
    output ap_axis_iarg_124_tvalid,
    output [S_AXIS_IARG_124_WIDTH/8-1:0] ap_axis_iarg_124_tkeep,
    output [S_AXIS_IARG_124_WIDTH/8-1:0] ap_axis_iarg_124_tstrb,
    output [S_AXIS_IARG_124_WIDTH-1:0] ap_axis_iarg_124_tdata,
    //input AXI-Stream pass-through interface 125
    input s_axis_iarg_125_aclk,
    input s_axis_iarg_125_aresetn,
    input s_axis_iarg_125_tlast,
    input s_axis_iarg_125_tvalid,
    input [S_AXIS_IARG_125_DMWIDTH/8-1:0] s_axis_iarg_125_tkeep,
    input [S_AXIS_IARG_125_DMWIDTH/8-1:0] s_axis_iarg_125_tstrb,
    input [S_AXIS_IARG_125_DMWIDTH-1:0] s_axis_iarg_125_tdata,
    output s_axis_iarg_125_tready,
    input ap_axis_iarg_125_tready,
    output ap_axis_iarg_125_tlast,
    output ap_axis_iarg_125_tvalid,
    output [S_AXIS_IARG_125_WIDTH/8-1:0] ap_axis_iarg_125_tkeep,
    output [S_AXIS_IARG_125_WIDTH/8-1:0] ap_axis_iarg_125_tstrb,
    output [S_AXIS_IARG_125_WIDTH-1:0] ap_axis_iarg_125_tdata,
    //input AXI-Stream pass-through interface 126
    input s_axis_iarg_126_aclk,
    input s_axis_iarg_126_aresetn,
    input s_axis_iarg_126_tlast,
    input s_axis_iarg_126_tvalid,
    input [S_AXIS_IARG_126_DMWIDTH/8-1:0] s_axis_iarg_126_tkeep,
    input [S_AXIS_IARG_126_DMWIDTH/8-1:0] s_axis_iarg_126_tstrb,
    input [S_AXIS_IARG_126_DMWIDTH-1:0] s_axis_iarg_126_tdata,
    output s_axis_iarg_126_tready,
    input ap_axis_iarg_126_tready,
    output ap_axis_iarg_126_tlast,
    output ap_axis_iarg_126_tvalid,
    output [S_AXIS_IARG_126_WIDTH/8-1:0] ap_axis_iarg_126_tkeep,
    output [S_AXIS_IARG_126_WIDTH/8-1:0] ap_axis_iarg_126_tstrb,
    output [S_AXIS_IARG_126_WIDTH-1:0] ap_axis_iarg_126_tdata,
    //input AXI-Stream pass-through interface 127
    input s_axis_iarg_127_aclk,
    input s_axis_iarg_127_aresetn,
    input s_axis_iarg_127_tlast,
    input s_axis_iarg_127_tvalid,
    input [S_AXIS_IARG_127_DMWIDTH/8-1:0] s_axis_iarg_127_tkeep,
    input [S_AXIS_IARG_127_DMWIDTH/8-1:0] s_axis_iarg_127_tstrb,
    input [S_AXIS_IARG_127_DMWIDTH-1:0] s_axis_iarg_127_tdata,
    output s_axis_iarg_127_tready,
    input ap_axis_iarg_127_tready,
    output ap_axis_iarg_127_tlast,
    output ap_axis_iarg_127_tvalid,
    output [S_AXIS_IARG_127_WIDTH/8-1:0] ap_axis_iarg_127_tkeep,
    output [S_AXIS_IARG_127_WIDTH/8-1:0] ap_axis_iarg_127_tstrb,
    output [S_AXIS_IARG_127_WIDTH-1:0] ap_axis_iarg_127_tdata,
    //-----------------------------------------------------
    //output AXI-Stream pass-through interface 0
    input m_axis_oarg_0_aclk,
    input m_axis_oarg_0_aresetn,
    output m_axis_oarg_0_tlast,
    output m_axis_oarg_0_tvalid,
    output [M_AXIS_OARG_0_DMWIDTH/8-1:0] m_axis_oarg_0_tkeep,
    output [M_AXIS_OARG_0_DMWIDTH/8-1:0] m_axis_oarg_0_tstrb,
    output [M_AXIS_OARG_0_DMWIDTH-1:0] m_axis_oarg_0_tdata,
    input m_axis_oarg_0_tready,
    input ap_axis_oarg_0_tlast,
    input ap_axis_oarg_0_tvalid,
    input [M_AXIS_OARG_0_WIDTH/8-1:0] ap_axis_oarg_0_tkeep,
    input [M_AXIS_OARG_0_WIDTH/8-1:0] ap_axis_oarg_0_tstrb,
    input [M_AXIS_OARG_0_WIDTH-1:0] ap_axis_oarg_0_tdata,
    output ap_axis_oarg_0_tready,
    //output AXI-Stream pass-through interface 1
    input m_axis_oarg_1_aclk,
    input m_axis_oarg_1_aresetn,
    output m_axis_oarg_1_tlast,
    output m_axis_oarg_1_tvalid,
    output [M_AXIS_OARG_1_DMWIDTH/8-1:0] m_axis_oarg_1_tkeep,
    output [M_AXIS_OARG_1_DMWIDTH/8-1:0] m_axis_oarg_1_tstrb,
    output [M_AXIS_OARG_1_DMWIDTH-1:0] m_axis_oarg_1_tdata,
    input m_axis_oarg_1_tready,
    input ap_axis_oarg_1_tlast,
    input ap_axis_oarg_1_tvalid,
    input [M_AXIS_OARG_1_WIDTH/8-1:0] ap_axis_oarg_1_tkeep,
    input [M_AXIS_OARG_1_WIDTH/8-1:0] ap_axis_oarg_1_tstrb,
    input [M_AXIS_OARG_1_WIDTH-1:0] ap_axis_oarg_1_tdata,
    output ap_axis_oarg_1_tready,
    //output AXI-Stream pass-through interface 2
    input m_axis_oarg_2_aclk,
    input m_axis_oarg_2_aresetn,
    output m_axis_oarg_2_tlast,
    output m_axis_oarg_2_tvalid,
    output [M_AXIS_OARG_2_DMWIDTH/8-1:0] m_axis_oarg_2_tkeep,
    output [M_AXIS_OARG_2_DMWIDTH/8-1:0] m_axis_oarg_2_tstrb,
    output [M_AXIS_OARG_2_DMWIDTH-1:0] m_axis_oarg_2_tdata,
    input m_axis_oarg_2_tready,
    input ap_axis_oarg_2_tlast,
    input ap_axis_oarg_2_tvalid,
    input [M_AXIS_OARG_2_WIDTH/8-1:0] ap_axis_oarg_2_tkeep,
    input [M_AXIS_OARG_2_WIDTH/8-1:0] ap_axis_oarg_2_tstrb,
    input [M_AXIS_OARG_2_WIDTH-1:0] ap_axis_oarg_2_tdata,
    output ap_axis_oarg_2_tready,
    //output AXI-Stream pass-through interface 3
    input m_axis_oarg_3_aclk,
    input m_axis_oarg_3_aresetn,
    output m_axis_oarg_3_tlast,
    output m_axis_oarg_3_tvalid,
    output [M_AXIS_OARG_3_DMWIDTH/8-1:0] m_axis_oarg_3_tkeep,
    output [M_AXIS_OARG_3_DMWIDTH/8-1:0] m_axis_oarg_3_tstrb,
    output [M_AXIS_OARG_3_DMWIDTH-1:0] m_axis_oarg_3_tdata,
    input m_axis_oarg_3_tready,
    input ap_axis_oarg_3_tlast,
    input ap_axis_oarg_3_tvalid,
    input [M_AXIS_OARG_3_WIDTH/8-1:0] ap_axis_oarg_3_tkeep,
    input [M_AXIS_OARG_3_WIDTH/8-1:0] ap_axis_oarg_3_tstrb,
    input [M_AXIS_OARG_3_WIDTH-1:0] ap_axis_oarg_3_tdata,
    output ap_axis_oarg_3_tready,
    //output AXI-Stream pass-through interface 4
    input m_axis_oarg_4_aclk,
    input m_axis_oarg_4_aresetn,
    output m_axis_oarg_4_tlast,
    output m_axis_oarg_4_tvalid,
    output [M_AXIS_OARG_4_DMWIDTH/8-1:0] m_axis_oarg_4_tkeep,
    output [M_AXIS_OARG_4_DMWIDTH/8-1:0] m_axis_oarg_4_tstrb,
    output [M_AXIS_OARG_4_DMWIDTH-1:0] m_axis_oarg_4_tdata,
    input m_axis_oarg_4_tready,
    input ap_axis_oarg_4_tlast,
    input ap_axis_oarg_4_tvalid,
    input [M_AXIS_OARG_4_WIDTH/8-1:0] ap_axis_oarg_4_tkeep,
    input [M_AXIS_OARG_4_WIDTH/8-1:0] ap_axis_oarg_4_tstrb,
    input [M_AXIS_OARG_4_WIDTH-1:0] ap_axis_oarg_4_tdata,
    output ap_axis_oarg_4_tready,
    //output AXI-Stream pass-through interface 5
    input m_axis_oarg_5_aclk,
    input m_axis_oarg_5_aresetn,
    output m_axis_oarg_5_tlast,
    output m_axis_oarg_5_tvalid,
    output [M_AXIS_OARG_5_DMWIDTH/8-1:0] m_axis_oarg_5_tkeep,
    output [M_AXIS_OARG_5_DMWIDTH/8-1:0] m_axis_oarg_5_tstrb,
    output [M_AXIS_OARG_5_DMWIDTH-1:0] m_axis_oarg_5_tdata,
    input m_axis_oarg_5_tready,
    input ap_axis_oarg_5_tlast,
    input ap_axis_oarg_5_tvalid,
    input [M_AXIS_OARG_5_WIDTH/8-1:0] ap_axis_oarg_5_tkeep,
    input [M_AXIS_OARG_5_WIDTH/8-1:0] ap_axis_oarg_5_tstrb,
    input [M_AXIS_OARG_5_WIDTH-1:0] ap_axis_oarg_5_tdata,
    output ap_axis_oarg_5_tready,
    //output AXI-Stream pass-through interface 6
    input m_axis_oarg_6_aclk,
    input m_axis_oarg_6_aresetn,
    output m_axis_oarg_6_tlast,
    output m_axis_oarg_6_tvalid,
    output [M_AXIS_OARG_6_DMWIDTH/8-1:0] m_axis_oarg_6_tkeep,
    output [M_AXIS_OARG_6_DMWIDTH/8-1:0] m_axis_oarg_6_tstrb,
    output [M_AXIS_OARG_6_DMWIDTH-1:0] m_axis_oarg_6_tdata,
    input m_axis_oarg_6_tready,
    input ap_axis_oarg_6_tlast,
    input ap_axis_oarg_6_tvalid,
    input [M_AXIS_OARG_6_WIDTH/8-1:0] ap_axis_oarg_6_tkeep,
    input [M_AXIS_OARG_6_WIDTH/8-1:0] ap_axis_oarg_6_tstrb,
    input [M_AXIS_OARG_6_WIDTH-1:0] ap_axis_oarg_6_tdata,
    output ap_axis_oarg_6_tready,
    //output AXI-Stream pass-through interface 7
    input m_axis_oarg_7_aclk,
    input m_axis_oarg_7_aresetn,
    output m_axis_oarg_7_tlast,
    output m_axis_oarg_7_tvalid,
    output [M_AXIS_OARG_7_DMWIDTH/8-1:0] m_axis_oarg_7_tkeep,
    output [M_AXIS_OARG_7_DMWIDTH/8-1:0] m_axis_oarg_7_tstrb,
    output [M_AXIS_OARG_7_DMWIDTH-1:0] m_axis_oarg_7_tdata,
    input m_axis_oarg_7_tready,
    input ap_axis_oarg_7_tlast,
    input ap_axis_oarg_7_tvalid,
    input [M_AXIS_OARG_7_WIDTH/8-1:0] ap_axis_oarg_7_tkeep,
    input [M_AXIS_OARG_7_WIDTH/8-1:0] ap_axis_oarg_7_tstrb,
    input [M_AXIS_OARG_7_WIDTH-1:0] ap_axis_oarg_7_tdata,
    output ap_axis_oarg_7_tready,
    //output AXI-Stream pass-through interface 8
    input m_axis_oarg_8_aclk,
    input m_axis_oarg_8_aresetn,
    output m_axis_oarg_8_tlast,
    output m_axis_oarg_8_tvalid,
    output [M_AXIS_OARG_8_DMWIDTH/8-1:0] m_axis_oarg_8_tkeep,
    output [M_AXIS_OARG_8_DMWIDTH/8-1:0] m_axis_oarg_8_tstrb,
    output [M_AXIS_OARG_8_DMWIDTH-1:0] m_axis_oarg_8_tdata,
    input m_axis_oarg_8_tready,
    input ap_axis_oarg_8_tlast,
    input ap_axis_oarg_8_tvalid,
    input [M_AXIS_OARG_8_WIDTH/8-1:0] ap_axis_oarg_8_tkeep,
    input [M_AXIS_OARG_8_WIDTH/8-1:0] ap_axis_oarg_8_tstrb,
    input [M_AXIS_OARG_8_WIDTH-1:0] ap_axis_oarg_8_tdata,
    output ap_axis_oarg_8_tready,
    //output AXI-Stream pass-through interface 9
    input m_axis_oarg_9_aclk,
    input m_axis_oarg_9_aresetn,
    output m_axis_oarg_9_tlast,
    output m_axis_oarg_9_tvalid,
    output [M_AXIS_OARG_9_DMWIDTH/8-1:0] m_axis_oarg_9_tkeep,
    output [M_AXIS_OARG_9_DMWIDTH/8-1:0] m_axis_oarg_9_tstrb,
    output [M_AXIS_OARG_9_DMWIDTH-1:0] m_axis_oarg_9_tdata,
    input m_axis_oarg_9_tready,
    input ap_axis_oarg_9_tlast,
    input ap_axis_oarg_9_tvalid,
    input [M_AXIS_OARG_9_WIDTH/8-1:0] ap_axis_oarg_9_tkeep,
    input [M_AXIS_OARG_9_WIDTH/8-1:0] ap_axis_oarg_9_tstrb,
    input [M_AXIS_OARG_9_WIDTH-1:0] ap_axis_oarg_9_tdata,
    output ap_axis_oarg_9_tready,
    //output AXI-Stream pass-through interface 10
    input m_axis_oarg_10_aclk,
    input m_axis_oarg_10_aresetn,
    output m_axis_oarg_10_tlast,
    output m_axis_oarg_10_tvalid,
    output [M_AXIS_OARG_10_DMWIDTH/8-1:0] m_axis_oarg_10_tkeep,
    output [M_AXIS_OARG_10_DMWIDTH/8-1:0] m_axis_oarg_10_tstrb,
    output [M_AXIS_OARG_10_DMWIDTH-1:0] m_axis_oarg_10_tdata,
    input m_axis_oarg_10_tready,
    input ap_axis_oarg_10_tlast,
    input ap_axis_oarg_10_tvalid,
    input [M_AXIS_OARG_10_WIDTH/8-1:0] ap_axis_oarg_10_tkeep,
    input [M_AXIS_OARG_10_WIDTH/8-1:0] ap_axis_oarg_10_tstrb,
    input [M_AXIS_OARG_10_WIDTH-1:0] ap_axis_oarg_10_tdata,
    output ap_axis_oarg_10_tready,
    //output AXI-Stream pass-through interface 11
    input m_axis_oarg_11_aclk,
    input m_axis_oarg_11_aresetn,
    output m_axis_oarg_11_tlast,
    output m_axis_oarg_11_tvalid,
    output [M_AXIS_OARG_11_DMWIDTH/8-1:0] m_axis_oarg_11_tkeep,
    output [M_AXIS_OARG_11_DMWIDTH/8-1:0] m_axis_oarg_11_tstrb,
    output [M_AXIS_OARG_11_DMWIDTH-1:0] m_axis_oarg_11_tdata,
    input m_axis_oarg_11_tready,
    input ap_axis_oarg_11_tlast,
    input ap_axis_oarg_11_tvalid,
    input [M_AXIS_OARG_11_WIDTH/8-1:0] ap_axis_oarg_11_tkeep,
    input [M_AXIS_OARG_11_WIDTH/8-1:0] ap_axis_oarg_11_tstrb,
    input [M_AXIS_OARG_11_WIDTH-1:0] ap_axis_oarg_11_tdata,
    output ap_axis_oarg_11_tready,
    //output AXI-Stream pass-through interface 12
    input m_axis_oarg_12_aclk,
    input m_axis_oarg_12_aresetn,
    output m_axis_oarg_12_tlast,
    output m_axis_oarg_12_tvalid,
    output [M_AXIS_OARG_12_DMWIDTH/8-1:0] m_axis_oarg_12_tkeep,
    output [M_AXIS_OARG_12_DMWIDTH/8-1:0] m_axis_oarg_12_tstrb,
    output [M_AXIS_OARG_12_DMWIDTH-1:0] m_axis_oarg_12_tdata,
    input m_axis_oarg_12_tready,
    input ap_axis_oarg_12_tlast,
    input ap_axis_oarg_12_tvalid,
    input [M_AXIS_OARG_12_WIDTH/8-1:0] ap_axis_oarg_12_tkeep,
    input [M_AXIS_OARG_12_WIDTH/8-1:0] ap_axis_oarg_12_tstrb,
    input [M_AXIS_OARG_12_WIDTH-1:0] ap_axis_oarg_12_tdata,
    output ap_axis_oarg_12_tready,
    //output AXI-Stream pass-through interface 13
    input m_axis_oarg_13_aclk,
    input m_axis_oarg_13_aresetn,
    output m_axis_oarg_13_tlast,
    output m_axis_oarg_13_tvalid,
    output [M_AXIS_OARG_13_DMWIDTH/8-1:0] m_axis_oarg_13_tkeep,
    output [M_AXIS_OARG_13_DMWIDTH/8-1:0] m_axis_oarg_13_tstrb,
    output [M_AXIS_OARG_13_DMWIDTH-1:0] m_axis_oarg_13_tdata,
    input m_axis_oarg_13_tready,
    input ap_axis_oarg_13_tlast,
    input ap_axis_oarg_13_tvalid,
    input [M_AXIS_OARG_13_WIDTH/8-1:0] ap_axis_oarg_13_tkeep,
    input [M_AXIS_OARG_13_WIDTH/8-1:0] ap_axis_oarg_13_tstrb,
    input [M_AXIS_OARG_13_WIDTH-1:0] ap_axis_oarg_13_tdata,
    output ap_axis_oarg_13_tready,
    //output AXI-Stream pass-through interface 14
    input m_axis_oarg_14_aclk,
    input m_axis_oarg_14_aresetn,
    output m_axis_oarg_14_tlast,
    output m_axis_oarg_14_tvalid,
    output [M_AXIS_OARG_14_DMWIDTH/8-1:0] m_axis_oarg_14_tkeep,
    output [M_AXIS_OARG_14_DMWIDTH/8-1:0] m_axis_oarg_14_tstrb,
    output [M_AXIS_OARG_14_DMWIDTH-1:0] m_axis_oarg_14_tdata,
    input m_axis_oarg_14_tready,
    input ap_axis_oarg_14_tlast,
    input ap_axis_oarg_14_tvalid,
    input [M_AXIS_OARG_14_WIDTH/8-1:0] ap_axis_oarg_14_tkeep,
    input [M_AXIS_OARG_14_WIDTH/8-1:0] ap_axis_oarg_14_tstrb,
    input [M_AXIS_OARG_14_WIDTH-1:0] ap_axis_oarg_14_tdata,
    output ap_axis_oarg_14_tready,
    //output AXI-Stream pass-through interface 15
    input m_axis_oarg_15_aclk,
    input m_axis_oarg_15_aresetn,
    output m_axis_oarg_15_tlast,
    output m_axis_oarg_15_tvalid,
    output [M_AXIS_OARG_15_DMWIDTH/8-1:0] m_axis_oarg_15_tkeep,
    output [M_AXIS_OARG_15_DMWIDTH/8-1:0] m_axis_oarg_15_tstrb,
    output [M_AXIS_OARG_15_DMWIDTH-1:0] m_axis_oarg_15_tdata,
    input m_axis_oarg_15_tready,
    input ap_axis_oarg_15_tlast,
    input ap_axis_oarg_15_tvalid,
    input [M_AXIS_OARG_15_WIDTH/8-1:0] ap_axis_oarg_15_tkeep,
    input [M_AXIS_OARG_15_WIDTH/8-1:0] ap_axis_oarg_15_tstrb,
    input [M_AXIS_OARG_15_WIDTH-1:0] ap_axis_oarg_15_tdata,
    output ap_axis_oarg_15_tready,
    //output AXI-Stream pass-through interface 16
    input m_axis_oarg_16_aclk,
    input m_axis_oarg_16_aresetn,
    output m_axis_oarg_16_tlast,
    output m_axis_oarg_16_tvalid,
    output [M_AXIS_OARG_16_DMWIDTH/8-1:0] m_axis_oarg_16_tkeep,
    output [M_AXIS_OARG_16_DMWIDTH/8-1:0] m_axis_oarg_16_tstrb,
    output [M_AXIS_OARG_16_DMWIDTH-1:0] m_axis_oarg_16_tdata,
    input m_axis_oarg_16_tready,
    input ap_axis_oarg_16_tlast,
    input ap_axis_oarg_16_tvalid,
    input [M_AXIS_OARG_16_WIDTH/8-1:0] ap_axis_oarg_16_tkeep,
    input [M_AXIS_OARG_16_WIDTH/8-1:0] ap_axis_oarg_16_tstrb,
    input [M_AXIS_OARG_16_WIDTH-1:0] ap_axis_oarg_16_tdata,
    output ap_axis_oarg_16_tready,
    //output AXI-Stream pass-through interface 17
    input m_axis_oarg_17_aclk,
    input m_axis_oarg_17_aresetn,
    output m_axis_oarg_17_tlast,
    output m_axis_oarg_17_tvalid,
    output [M_AXIS_OARG_17_DMWIDTH/8-1:0] m_axis_oarg_17_tkeep,
    output [M_AXIS_OARG_17_DMWIDTH/8-1:0] m_axis_oarg_17_tstrb,
    output [M_AXIS_OARG_17_DMWIDTH-1:0] m_axis_oarg_17_tdata,
    input m_axis_oarg_17_tready,
    input ap_axis_oarg_17_tlast,
    input ap_axis_oarg_17_tvalid,
    input [M_AXIS_OARG_17_WIDTH/8-1:0] ap_axis_oarg_17_tkeep,
    input [M_AXIS_OARG_17_WIDTH/8-1:0] ap_axis_oarg_17_tstrb,
    input [M_AXIS_OARG_17_WIDTH-1:0] ap_axis_oarg_17_tdata,
    output ap_axis_oarg_17_tready,
    //output AXI-Stream pass-through interface 18
    input m_axis_oarg_18_aclk,
    input m_axis_oarg_18_aresetn,
    output m_axis_oarg_18_tlast,
    output m_axis_oarg_18_tvalid,
    output [M_AXIS_OARG_18_DMWIDTH/8-1:0] m_axis_oarg_18_tkeep,
    output [M_AXIS_OARG_18_DMWIDTH/8-1:0] m_axis_oarg_18_tstrb,
    output [M_AXIS_OARG_18_DMWIDTH-1:0] m_axis_oarg_18_tdata,
    input m_axis_oarg_18_tready,
    input ap_axis_oarg_18_tlast,
    input ap_axis_oarg_18_tvalid,
    input [M_AXIS_OARG_18_WIDTH/8-1:0] ap_axis_oarg_18_tkeep,
    input [M_AXIS_OARG_18_WIDTH/8-1:0] ap_axis_oarg_18_tstrb,
    input [M_AXIS_OARG_18_WIDTH-1:0] ap_axis_oarg_18_tdata,
    output ap_axis_oarg_18_tready,
    //output AXI-Stream pass-through interface 19
    input m_axis_oarg_19_aclk,
    input m_axis_oarg_19_aresetn,
    output m_axis_oarg_19_tlast,
    output m_axis_oarg_19_tvalid,
    output [M_AXIS_OARG_19_DMWIDTH/8-1:0] m_axis_oarg_19_tkeep,
    output [M_AXIS_OARG_19_DMWIDTH/8-1:0] m_axis_oarg_19_tstrb,
    output [M_AXIS_OARG_19_DMWIDTH-1:0] m_axis_oarg_19_tdata,
    input m_axis_oarg_19_tready,
    input ap_axis_oarg_19_tlast,
    input ap_axis_oarg_19_tvalid,
    input [M_AXIS_OARG_19_WIDTH/8-1:0] ap_axis_oarg_19_tkeep,
    input [M_AXIS_OARG_19_WIDTH/8-1:0] ap_axis_oarg_19_tstrb,
    input [M_AXIS_OARG_19_WIDTH-1:0] ap_axis_oarg_19_tdata,
    output ap_axis_oarg_19_tready,
    //output AXI-Stream pass-through interface 20
    input m_axis_oarg_20_aclk,
    input m_axis_oarg_20_aresetn,
    output m_axis_oarg_20_tlast,
    output m_axis_oarg_20_tvalid,
    output [M_AXIS_OARG_20_DMWIDTH/8-1:0] m_axis_oarg_20_tkeep,
    output [M_AXIS_OARG_20_DMWIDTH/8-1:0] m_axis_oarg_20_tstrb,
    output [M_AXIS_OARG_20_DMWIDTH-1:0] m_axis_oarg_20_tdata,
    input m_axis_oarg_20_tready,
    input ap_axis_oarg_20_tlast,
    input ap_axis_oarg_20_tvalid,
    input [M_AXIS_OARG_20_WIDTH/8-1:0] ap_axis_oarg_20_tkeep,
    input [M_AXIS_OARG_20_WIDTH/8-1:0] ap_axis_oarg_20_tstrb,
    input [M_AXIS_OARG_20_WIDTH-1:0] ap_axis_oarg_20_tdata,
    output ap_axis_oarg_20_tready,
    //output AXI-Stream pass-through interface 21
    input m_axis_oarg_21_aclk,
    input m_axis_oarg_21_aresetn,
    output m_axis_oarg_21_tlast,
    output m_axis_oarg_21_tvalid,
    output [M_AXIS_OARG_21_DMWIDTH/8-1:0] m_axis_oarg_21_tkeep,
    output [M_AXIS_OARG_21_DMWIDTH/8-1:0] m_axis_oarg_21_tstrb,
    output [M_AXIS_OARG_21_DMWIDTH-1:0] m_axis_oarg_21_tdata,
    input m_axis_oarg_21_tready,
    input ap_axis_oarg_21_tlast,
    input ap_axis_oarg_21_tvalid,
    input [M_AXIS_OARG_21_WIDTH/8-1:0] ap_axis_oarg_21_tkeep,
    input [M_AXIS_OARG_21_WIDTH/8-1:0] ap_axis_oarg_21_tstrb,
    input [M_AXIS_OARG_21_WIDTH-1:0] ap_axis_oarg_21_tdata,
    output ap_axis_oarg_21_tready,
    //output AXI-Stream pass-through interface 22
    input m_axis_oarg_22_aclk,
    input m_axis_oarg_22_aresetn,
    output m_axis_oarg_22_tlast,
    output m_axis_oarg_22_tvalid,
    output [M_AXIS_OARG_22_DMWIDTH/8-1:0] m_axis_oarg_22_tkeep,
    output [M_AXIS_OARG_22_DMWIDTH/8-1:0] m_axis_oarg_22_tstrb,
    output [M_AXIS_OARG_22_DMWIDTH-1:0] m_axis_oarg_22_tdata,
    input m_axis_oarg_22_tready,
    input ap_axis_oarg_22_tlast,
    input ap_axis_oarg_22_tvalid,
    input [M_AXIS_OARG_22_WIDTH/8-1:0] ap_axis_oarg_22_tkeep,
    input [M_AXIS_OARG_22_WIDTH/8-1:0] ap_axis_oarg_22_tstrb,
    input [M_AXIS_OARG_22_WIDTH-1:0] ap_axis_oarg_22_tdata,
    output ap_axis_oarg_22_tready,
    //output AXI-Stream pass-through interface 23
    input m_axis_oarg_23_aclk,
    input m_axis_oarg_23_aresetn,
    output m_axis_oarg_23_tlast,
    output m_axis_oarg_23_tvalid,
    output [M_AXIS_OARG_23_DMWIDTH/8-1:0] m_axis_oarg_23_tkeep,
    output [M_AXIS_OARG_23_DMWIDTH/8-1:0] m_axis_oarg_23_tstrb,
    output [M_AXIS_OARG_23_DMWIDTH-1:0] m_axis_oarg_23_tdata,
    input m_axis_oarg_23_tready,
    input ap_axis_oarg_23_tlast,
    input ap_axis_oarg_23_tvalid,
    input [M_AXIS_OARG_23_WIDTH/8-1:0] ap_axis_oarg_23_tkeep,
    input [M_AXIS_OARG_23_WIDTH/8-1:0] ap_axis_oarg_23_tstrb,
    input [M_AXIS_OARG_23_WIDTH-1:0] ap_axis_oarg_23_tdata,
    output ap_axis_oarg_23_tready,
    //output AXI-Stream pass-through interface 24
    input m_axis_oarg_24_aclk,
    input m_axis_oarg_24_aresetn,
    output m_axis_oarg_24_tlast,
    output m_axis_oarg_24_tvalid,
    output [M_AXIS_OARG_24_DMWIDTH/8-1:0] m_axis_oarg_24_tkeep,
    output [M_AXIS_OARG_24_DMWIDTH/8-1:0] m_axis_oarg_24_tstrb,
    output [M_AXIS_OARG_24_DMWIDTH-1:0] m_axis_oarg_24_tdata,
    input m_axis_oarg_24_tready,
    input ap_axis_oarg_24_tlast,
    input ap_axis_oarg_24_tvalid,
    input [M_AXIS_OARG_24_WIDTH/8-1:0] ap_axis_oarg_24_tkeep,
    input [M_AXIS_OARG_24_WIDTH/8-1:0] ap_axis_oarg_24_tstrb,
    input [M_AXIS_OARG_24_WIDTH-1:0] ap_axis_oarg_24_tdata,
    output ap_axis_oarg_24_tready,
    //output AXI-Stream pass-through interface 25
    input m_axis_oarg_25_aclk,
    input m_axis_oarg_25_aresetn,
    output m_axis_oarg_25_tlast,
    output m_axis_oarg_25_tvalid,
    output [M_AXIS_OARG_25_DMWIDTH/8-1:0] m_axis_oarg_25_tkeep,
    output [M_AXIS_OARG_25_DMWIDTH/8-1:0] m_axis_oarg_25_tstrb,
    output [M_AXIS_OARG_25_DMWIDTH-1:0] m_axis_oarg_25_tdata,
    input m_axis_oarg_25_tready,
    input ap_axis_oarg_25_tlast,
    input ap_axis_oarg_25_tvalid,
    input [M_AXIS_OARG_25_WIDTH/8-1:0] ap_axis_oarg_25_tkeep,
    input [M_AXIS_OARG_25_WIDTH/8-1:0] ap_axis_oarg_25_tstrb,
    input [M_AXIS_OARG_25_WIDTH-1:0] ap_axis_oarg_25_tdata,
    output ap_axis_oarg_25_tready,
    //output AXI-Stream pass-through interface 26
    input m_axis_oarg_26_aclk,
    input m_axis_oarg_26_aresetn,
    output m_axis_oarg_26_tlast,
    output m_axis_oarg_26_tvalid,
    output [M_AXIS_OARG_26_DMWIDTH/8-1:0] m_axis_oarg_26_tkeep,
    output [M_AXIS_OARG_26_DMWIDTH/8-1:0] m_axis_oarg_26_tstrb,
    output [M_AXIS_OARG_26_DMWIDTH-1:0] m_axis_oarg_26_tdata,
    input m_axis_oarg_26_tready,
    input ap_axis_oarg_26_tlast,
    input ap_axis_oarg_26_tvalid,
    input [M_AXIS_OARG_26_WIDTH/8-1:0] ap_axis_oarg_26_tkeep,
    input [M_AXIS_OARG_26_WIDTH/8-1:0] ap_axis_oarg_26_tstrb,
    input [M_AXIS_OARG_26_WIDTH-1:0] ap_axis_oarg_26_tdata,
    output ap_axis_oarg_26_tready,
    //output AXI-Stream pass-through interface 27
    input m_axis_oarg_27_aclk,
    input m_axis_oarg_27_aresetn,
    output m_axis_oarg_27_tlast,
    output m_axis_oarg_27_tvalid,
    output [M_AXIS_OARG_27_DMWIDTH/8-1:0] m_axis_oarg_27_tkeep,
    output [M_AXIS_OARG_27_DMWIDTH/8-1:0] m_axis_oarg_27_tstrb,
    output [M_AXIS_OARG_27_DMWIDTH-1:0] m_axis_oarg_27_tdata,
    input m_axis_oarg_27_tready,
    input ap_axis_oarg_27_tlast,
    input ap_axis_oarg_27_tvalid,
    input [M_AXIS_OARG_27_WIDTH/8-1:0] ap_axis_oarg_27_tkeep,
    input [M_AXIS_OARG_27_WIDTH/8-1:0] ap_axis_oarg_27_tstrb,
    input [M_AXIS_OARG_27_WIDTH-1:0] ap_axis_oarg_27_tdata,
    output ap_axis_oarg_27_tready,
    //output AXI-Stream pass-through interface 28
    input m_axis_oarg_28_aclk,
    input m_axis_oarg_28_aresetn,
    output m_axis_oarg_28_tlast,
    output m_axis_oarg_28_tvalid,
    output [M_AXIS_OARG_28_DMWIDTH/8-1:0] m_axis_oarg_28_tkeep,
    output [M_AXIS_OARG_28_DMWIDTH/8-1:0] m_axis_oarg_28_tstrb,
    output [M_AXIS_OARG_28_DMWIDTH-1:0] m_axis_oarg_28_tdata,
    input m_axis_oarg_28_tready,
    input ap_axis_oarg_28_tlast,
    input ap_axis_oarg_28_tvalid,
    input [M_AXIS_OARG_28_WIDTH/8-1:0] ap_axis_oarg_28_tkeep,
    input [M_AXIS_OARG_28_WIDTH/8-1:0] ap_axis_oarg_28_tstrb,
    input [M_AXIS_OARG_28_WIDTH-1:0] ap_axis_oarg_28_tdata,
    output ap_axis_oarg_28_tready,
    //output AXI-Stream pass-through interface 29
    input m_axis_oarg_29_aclk,
    input m_axis_oarg_29_aresetn,
    output m_axis_oarg_29_tlast,
    output m_axis_oarg_29_tvalid,
    output [M_AXIS_OARG_29_DMWIDTH/8-1:0] m_axis_oarg_29_tkeep,
    output [M_AXIS_OARG_29_DMWIDTH/8-1:0] m_axis_oarg_29_tstrb,
    output [M_AXIS_OARG_29_DMWIDTH-1:0] m_axis_oarg_29_tdata,
    input m_axis_oarg_29_tready,
    input ap_axis_oarg_29_tlast,
    input ap_axis_oarg_29_tvalid,
    input [M_AXIS_OARG_29_WIDTH/8-1:0] ap_axis_oarg_29_tkeep,
    input [M_AXIS_OARG_29_WIDTH/8-1:0] ap_axis_oarg_29_tstrb,
    input [M_AXIS_OARG_29_WIDTH-1:0] ap_axis_oarg_29_tdata,
    output ap_axis_oarg_29_tready,
    //output AXI-Stream pass-through interface 30
    input m_axis_oarg_30_aclk,
    input m_axis_oarg_30_aresetn,
    output m_axis_oarg_30_tlast,
    output m_axis_oarg_30_tvalid,
    output [M_AXIS_OARG_30_DMWIDTH/8-1:0] m_axis_oarg_30_tkeep,
    output [M_AXIS_OARG_30_DMWIDTH/8-1:0] m_axis_oarg_30_tstrb,
    output [M_AXIS_OARG_30_DMWIDTH-1:0] m_axis_oarg_30_tdata,
    input m_axis_oarg_30_tready,
    input ap_axis_oarg_30_tlast,
    input ap_axis_oarg_30_tvalid,
    input [M_AXIS_OARG_30_WIDTH/8-1:0] ap_axis_oarg_30_tkeep,
    input [M_AXIS_OARG_30_WIDTH/8-1:0] ap_axis_oarg_30_tstrb,
    input [M_AXIS_OARG_30_WIDTH-1:0] ap_axis_oarg_30_tdata,
    output ap_axis_oarg_30_tready,
    //output AXI-Stream pass-through interface 31
    input m_axis_oarg_31_aclk,
    input m_axis_oarg_31_aresetn,
    output m_axis_oarg_31_tlast,
    output m_axis_oarg_31_tvalid,
    output [M_AXIS_OARG_31_DMWIDTH/8-1:0] m_axis_oarg_31_tkeep,
    output [M_AXIS_OARG_31_DMWIDTH/8-1:0] m_axis_oarg_31_tstrb,
    output [M_AXIS_OARG_31_DMWIDTH-1:0] m_axis_oarg_31_tdata,
    input m_axis_oarg_31_tready,
    input ap_axis_oarg_31_tlast,
    input ap_axis_oarg_31_tvalid,
    input [M_AXIS_OARG_31_WIDTH/8-1:0] ap_axis_oarg_31_tkeep,
    input [M_AXIS_OARG_31_WIDTH/8-1:0] ap_axis_oarg_31_tstrb,
    input [M_AXIS_OARG_31_WIDTH-1:0] ap_axis_oarg_31_tdata,
    output ap_axis_oarg_31_tready,
    //output AXI-Stream pass-through interface 32
    input m_axis_oarg_32_aclk,
    input m_axis_oarg_32_aresetn,
    output m_axis_oarg_32_tlast,
    output m_axis_oarg_32_tvalid,
    output [M_AXIS_OARG_32_DMWIDTH/8-1:0] m_axis_oarg_32_tkeep,
    output [M_AXIS_OARG_32_DMWIDTH/8-1:0] m_axis_oarg_32_tstrb,
    output [M_AXIS_OARG_32_DMWIDTH-1:0] m_axis_oarg_32_tdata,
    input m_axis_oarg_32_tready,
    input ap_axis_oarg_32_tlast,
    input ap_axis_oarg_32_tvalid,
    input [M_AXIS_OARG_32_WIDTH/8-1:0] ap_axis_oarg_32_tkeep,
    input [M_AXIS_OARG_32_WIDTH/8-1:0] ap_axis_oarg_32_tstrb,
    input [M_AXIS_OARG_32_WIDTH-1:0] ap_axis_oarg_32_tdata,
    output ap_axis_oarg_32_tready,
    //output AXI-Stream pass-through interface 33
    input m_axis_oarg_33_aclk,
    input m_axis_oarg_33_aresetn,
    output m_axis_oarg_33_tlast,
    output m_axis_oarg_33_tvalid,
    output [M_AXIS_OARG_33_DMWIDTH/8-1:0] m_axis_oarg_33_tkeep,
    output [M_AXIS_OARG_33_DMWIDTH/8-1:0] m_axis_oarg_33_tstrb,
    output [M_AXIS_OARG_33_DMWIDTH-1:0] m_axis_oarg_33_tdata,
    input m_axis_oarg_33_tready,
    input ap_axis_oarg_33_tlast,
    input ap_axis_oarg_33_tvalid,
    input [M_AXIS_OARG_33_WIDTH/8-1:0] ap_axis_oarg_33_tkeep,
    input [M_AXIS_OARG_33_WIDTH/8-1:0] ap_axis_oarg_33_tstrb,
    input [M_AXIS_OARG_33_WIDTH-1:0] ap_axis_oarg_33_tdata,
    output ap_axis_oarg_33_tready,
    //output AXI-Stream pass-through interface 34
    input m_axis_oarg_34_aclk,
    input m_axis_oarg_34_aresetn,
    output m_axis_oarg_34_tlast,
    output m_axis_oarg_34_tvalid,
    output [M_AXIS_OARG_34_DMWIDTH/8-1:0] m_axis_oarg_34_tkeep,
    output [M_AXIS_OARG_34_DMWIDTH/8-1:0] m_axis_oarg_34_tstrb,
    output [M_AXIS_OARG_34_DMWIDTH-1:0] m_axis_oarg_34_tdata,
    input m_axis_oarg_34_tready,
    input ap_axis_oarg_34_tlast,
    input ap_axis_oarg_34_tvalid,
    input [M_AXIS_OARG_34_WIDTH/8-1:0] ap_axis_oarg_34_tkeep,
    input [M_AXIS_OARG_34_WIDTH/8-1:0] ap_axis_oarg_34_tstrb,
    input [M_AXIS_OARG_34_WIDTH-1:0] ap_axis_oarg_34_tdata,
    output ap_axis_oarg_34_tready,
    //output AXI-Stream pass-through interface 35
    input m_axis_oarg_35_aclk,
    input m_axis_oarg_35_aresetn,
    output m_axis_oarg_35_tlast,
    output m_axis_oarg_35_tvalid,
    output [M_AXIS_OARG_35_DMWIDTH/8-1:0] m_axis_oarg_35_tkeep,
    output [M_AXIS_OARG_35_DMWIDTH/8-1:0] m_axis_oarg_35_tstrb,
    output [M_AXIS_OARG_35_DMWIDTH-1:0] m_axis_oarg_35_tdata,
    input m_axis_oarg_35_tready,
    input ap_axis_oarg_35_tlast,
    input ap_axis_oarg_35_tvalid,
    input [M_AXIS_OARG_35_WIDTH/8-1:0] ap_axis_oarg_35_tkeep,
    input [M_AXIS_OARG_35_WIDTH/8-1:0] ap_axis_oarg_35_tstrb,
    input [M_AXIS_OARG_35_WIDTH-1:0] ap_axis_oarg_35_tdata,
    output ap_axis_oarg_35_tready,
    //output AXI-Stream pass-through interface 36
    input m_axis_oarg_36_aclk,
    input m_axis_oarg_36_aresetn,
    output m_axis_oarg_36_tlast,
    output m_axis_oarg_36_tvalid,
    output [M_AXIS_OARG_36_DMWIDTH/8-1:0] m_axis_oarg_36_tkeep,
    output [M_AXIS_OARG_36_DMWIDTH/8-1:0] m_axis_oarg_36_tstrb,
    output [M_AXIS_OARG_36_DMWIDTH-1:0] m_axis_oarg_36_tdata,
    input m_axis_oarg_36_tready,
    input ap_axis_oarg_36_tlast,
    input ap_axis_oarg_36_tvalid,
    input [M_AXIS_OARG_36_WIDTH/8-1:0] ap_axis_oarg_36_tkeep,
    input [M_AXIS_OARG_36_WIDTH/8-1:0] ap_axis_oarg_36_tstrb,
    input [M_AXIS_OARG_36_WIDTH-1:0] ap_axis_oarg_36_tdata,
    output ap_axis_oarg_36_tready,
    //output AXI-Stream pass-through interface 37
    input m_axis_oarg_37_aclk,
    input m_axis_oarg_37_aresetn,
    output m_axis_oarg_37_tlast,
    output m_axis_oarg_37_tvalid,
    output [M_AXIS_OARG_37_DMWIDTH/8-1:0] m_axis_oarg_37_tkeep,
    output [M_AXIS_OARG_37_DMWIDTH/8-1:0] m_axis_oarg_37_tstrb,
    output [M_AXIS_OARG_37_DMWIDTH-1:0] m_axis_oarg_37_tdata,
    input m_axis_oarg_37_tready,
    input ap_axis_oarg_37_tlast,
    input ap_axis_oarg_37_tvalid,
    input [M_AXIS_OARG_37_WIDTH/8-1:0] ap_axis_oarg_37_tkeep,
    input [M_AXIS_OARG_37_WIDTH/8-1:0] ap_axis_oarg_37_tstrb,
    input [M_AXIS_OARG_37_WIDTH-1:0] ap_axis_oarg_37_tdata,
    output ap_axis_oarg_37_tready,
    //output AXI-Stream pass-through interface 38
    input m_axis_oarg_38_aclk,
    input m_axis_oarg_38_aresetn,
    output m_axis_oarg_38_tlast,
    output m_axis_oarg_38_tvalid,
    output [M_AXIS_OARG_38_DMWIDTH/8-1:0] m_axis_oarg_38_tkeep,
    output [M_AXIS_OARG_38_DMWIDTH/8-1:0] m_axis_oarg_38_tstrb,
    output [M_AXIS_OARG_38_DMWIDTH-1:0] m_axis_oarg_38_tdata,
    input m_axis_oarg_38_tready,
    input ap_axis_oarg_38_tlast,
    input ap_axis_oarg_38_tvalid,
    input [M_AXIS_OARG_38_WIDTH/8-1:0] ap_axis_oarg_38_tkeep,
    input [M_AXIS_OARG_38_WIDTH/8-1:0] ap_axis_oarg_38_tstrb,
    input [M_AXIS_OARG_38_WIDTH-1:0] ap_axis_oarg_38_tdata,
    output ap_axis_oarg_38_tready,
    //output AXI-Stream pass-through interface 39
    input m_axis_oarg_39_aclk,
    input m_axis_oarg_39_aresetn,
    output m_axis_oarg_39_tlast,
    output m_axis_oarg_39_tvalid,
    output [M_AXIS_OARG_39_DMWIDTH/8-1:0] m_axis_oarg_39_tkeep,
    output [M_AXIS_OARG_39_DMWIDTH/8-1:0] m_axis_oarg_39_tstrb,
    output [M_AXIS_OARG_39_DMWIDTH-1:0] m_axis_oarg_39_tdata,
    input m_axis_oarg_39_tready,
    input ap_axis_oarg_39_tlast,
    input ap_axis_oarg_39_tvalid,
    input [M_AXIS_OARG_39_WIDTH/8-1:0] ap_axis_oarg_39_tkeep,
    input [M_AXIS_OARG_39_WIDTH/8-1:0] ap_axis_oarg_39_tstrb,
    input [M_AXIS_OARG_39_WIDTH-1:0] ap_axis_oarg_39_tdata,
    output ap_axis_oarg_39_tready,
    //output AXI-Stream pass-through interface 40
    input m_axis_oarg_40_aclk,
    input m_axis_oarg_40_aresetn,
    output m_axis_oarg_40_tlast,
    output m_axis_oarg_40_tvalid,
    output [M_AXIS_OARG_40_DMWIDTH/8-1:0] m_axis_oarg_40_tkeep,
    output [M_AXIS_OARG_40_DMWIDTH/8-1:0] m_axis_oarg_40_tstrb,
    output [M_AXIS_OARG_40_DMWIDTH-1:0] m_axis_oarg_40_tdata,
    input m_axis_oarg_40_tready,
    input ap_axis_oarg_40_tlast,
    input ap_axis_oarg_40_tvalid,
    input [M_AXIS_OARG_40_WIDTH/8-1:0] ap_axis_oarg_40_tkeep,
    input [M_AXIS_OARG_40_WIDTH/8-1:0] ap_axis_oarg_40_tstrb,
    input [M_AXIS_OARG_40_WIDTH-1:0] ap_axis_oarg_40_tdata,
    output ap_axis_oarg_40_tready,
    //output AXI-Stream pass-through interface 41
    input m_axis_oarg_41_aclk,
    input m_axis_oarg_41_aresetn,
    output m_axis_oarg_41_tlast,
    output m_axis_oarg_41_tvalid,
    output [M_AXIS_OARG_41_DMWIDTH/8-1:0] m_axis_oarg_41_tkeep,
    output [M_AXIS_OARG_41_DMWIDTH/8-1:0] m_axis_oarg_41_tstrb,
    output [M_AXIS_OARG_41_DMWIDTH-1:0] m_axis_oarg_41_tdata,
    input m_axis_oarg_41_tready,
    input ap_axis_oarg_41_tlast,
    input ap_axis_oarg_41_tvalid,
    input [M_AXIS_OARG_41_WIDTH/8-1:0] ap_axis_oarg_41_tkeep,
    input [M_AXIS_OARG_41_WIDTH/8-1:0] ap_axis_oarg_41_tstrb,
    input [M_AXIS_OARG_41_WIDTH-1:0] ap_axis_oarg_41_tdata,
    output ap_axis_oarg_41_tready,
    //output AXI-Stream pass-through interface 42
    input m_axis_oarg_42_aclk,
    input m_axis_oarg_42_aresetn,
    output m_axis_oarg_42_tlast,
    output m_axis_oarg_42_tvalid,
    output [M_AXIS_OARG_42_DMWIDTH/8-1:0] m_axis_oarg_42_tkeep,
    output [M_AXIS_OARG_42_DMWIDTH/8-1:0] m_axis_oarg_42_tstrb,
    output [M_AXIS_OARG_42_DMWIDTH-1:0] m_axis_oarg_42_tdata,
    input m_axis_oarg_42_tready,
    input ap_axis_oarg_42_tlast,
    input ap_axis_oarg_42_tvalid,
    input [M_AXIS_OARG_42_WIDTH/8-1:0] ap_axis_oarg_42_tkeep,
    input [M_AXIS_OARG_42_WIDTH/8-1:0] ap_axis_oarg_42_tstrb,
    input [M_AXIS_OARG_42_WIDTH-1:0] ap_axis_oarg_42_tdata,
    output ap_axis_oarg_42_tready,
    //output AXI-Stream pass-through interface 43
    input m_axis_oarg_43_aclk,
    input m_axis_oarg_43_aresetn,
    output m_axis_oarg_43_tlast,
    output m_axis_oarg_43_tvalid,
    output [M_AXIS_OARG_43_DMWIDTH/8-1:0] m_axis_oarg_43_tkeep,
    output [M_AXIS_OARG_43_DMWIDTH/8-1:0] m_axis_oarg_43_tstrb,
    output [M_AXIS_OARG_43_DMWIDTH-1:0] m_axis_oarg_43_tdata,
    input m_axis_oarg_43_tready,
    input ap_axis_oarg_43_tlast,
    input ap_axis_oarg_43_tvalid,
    input [M_AXIS_OARG_43_WIDTH/8-1:0] ap_axis_oarg_43_tkeep,
    input [M_AXIS_OARG_43_WIDTH/8-1:0] ap_axis_oarg_43_tstrb,
    input [M_AXIS_OARG_43_WIDTH-1:0] ap_axis_oarg_43_tdata,
    output ap_axis_oarg_43_tready,
    //output AXI-Stream pass-through interface 44
    input m_axis_oarg_44_aclk,
    input m_axis_oarg_44_aresetn,
    output m_axis_oarg_44_tlast,
    output m_axis_oarg_44_tvalid,
    output [M_AXIS_OARG_44_DMWIDTH/8-1:0] m_axis_oarg_44_tkeep,
    output [M_AXIS_OARG_44_DMWIDTH/8-1:0] m_axis_oarg_44_tstrb,
    output [M_AXIS_OARG_44_DMWIDTH-1:0] m_axis_oarg_44_tdata,
    input m_axis_oarg_44_tready,
    input ap_axis_oarg_44_tlast,
    input ap_axis_oarg_44_tvalid,
    input [M_AXIS_OARG_44_WIDTH/8-1:0] ap_axis_oarg_44_tkeep,
    input [M_AXIS_OARG_44_WIDTH/8-1:0] ap_axis_oarg_44_tstrb,
    input [M_AXIS_OARG_44_WIDTH-1:0] ap_axis_oarg_44_tdata,
    output ap_axis_oarg_44_tready,
    //output AXI-Stream pass-through interface 45
    input m_axis_oarg_45_aclk,
    input m_axis_oarg_45_aresetn,
    output m_axis_oarg_45_tlast,
    output m_axis_oarg_45_tvalid,
    output [M_AXIS_OARG_45_DMWIDTH/8-1:0] m_axis_oarg_45_tkeep,
    output [M_AXIS_OARG_45_DMWIDTH/8-1:0] m_axis_oarg_45_tstrb,
    output [M_AXIS_OARG_45_DMWIDTH-1:0] m_axis_oarg_45_tdata,
    input m_axis_oarg_45_tready,
    input ap_axis_oarg_45_tlast,
    input ap_axis_oarg_45_tvalid,
    input [M_AXIS_OARG_45_WIDTH/8-1:0] ap_axis_oarg_45_tkeep,
    input [M_AXIS_OARG_45_WIDTH/8-1:0] ap_axis_oarg_45_tstrb,
    input [M_AXIS_OARG_45_WIDTH-1:0] ap_axis_oarg_45_tdata,
    output ap_axis_oarg_45_tready,
    //output AXI-Stream pass-through interface 46
    input m_axis_oarg_46_aclk,
    input m_axis_oarg_46_aresetn,
    output m_axis_oarg_46_tlast,
    output m_axis_oarg_46_tvalid,
    output [M_AXIS_OARG_46_DMWIDTH/8-1:0] m_axis_oarg_46_tkeep,
    output [M_AXIS_OARG_46_DMWIDTH/8-1:0] m_axis_oarg_46_tstrb,
    output [M_AXIS_OARG_46_DMWIDTH-1:0] m_axis_oarg_46_tdata,
    input m_axis_oarg_46_tready,
    input ap_axis_oarg_46_tlast,
    input ap_axis_oarg_46_tvalid,
    input [M_AXIS_OARG_46_WIDTH/8-1:0] ap_axis_oarg_46_tkeep,
    input [M_AXIS_OARG_46_WIDTH/8-1:0] ap_axis_oarg_46_tstrb,
    input [M_AXIS_OARG_46_WIDTH-1:0] ap_axis_oarg_46_tdata,
    output ap_axis_oarg_46_tready,
    //output AXI-Stream pass-through interface 47
    input m_axis_oarg_47_aclk,
    input m_axis_oarg_47_aresetn,
    output m_axis_oarg_47_tlast,
    output m_axis_oarg_47_tvalid,
    output [M_AXIS_OARG_47_DMWIDTH/8-1:0] m_axis_oarg_47_tkeep,
    output [M_AXIS_OARG_47_DMWIDTH/8-1:0] m_axis_oarg_47_tstrb,
    output [M_AXIS_OARG_47_DMWIDTH-1:0] m_axis_oarg_47_tdata,
    input m_axis_oarg_47_tready,
    input ap_axis_oarg_47_tlast,
    input ap_axis_oarg_47_tvalid,
    input [M_AXIS_OARG_47_WIDTH/8-1:0] ap_axis_oarg_47_tkeep,
    input [M_AXIS_OARG_47_WIDTH/8-1:0] ap_axis_oarg_47_tstrb,
    input [M_AXIS_OARG_47_WIDTH-1:0] ap_axis_oarg_47_tdata,
    output ap_axis_oarg_47_tready,
    //output AXI-Stream pass-through interface 48
    input m_axis_oarg_48_aclk,
    input m_axis_oarg_48_aresetn,
    output m_axis_oarg_48_tlast,
    output m_axis_oarg_48_tvalid,
    output [M_AXIS_OARG_48_DMWIDTH/8-1:0] m_axis_oarg_48_tkeep,
    output [M_AXIS_OARG_48_DMWIDTH/8-1:0] m_axis_oarg_48_tstrb,
    output [M_AXIS_OARG_48_DMWIDTH-1:0] m_axis_oarg_48_tdata,
    input m_axis_oarg_48_tready,
    input ap_axis_oarg_48_tlast,
    input ap_axis_oarg_48_tvalid,
    input [M_AXIS_OARG_48_WIDTH/8-1:0] ap_axis_oarg_48_tkeep,
    input [M_AXIS_OARG_48_WIDTH/8-1:0] ap_axis_oarg_48_tstrb,
    input [M_AXIS_OARG_48_WIDTH-1:0] ap_axis_oarg_48_tdata,
    output ap_axis_oarg_48_tready,
    //output AXI-Stream pass-through interface 49
    input m_axis_oarg_49_aclk,
    input m_axis_oarg_49_aresetn,
    output m_axis_oarg_49_tlast,
    output m_axis_oarg_49_tvalid,
    output [M_AXIS_OARG_49_DMWIDTH/8-1:0] m_axis_oarg_49_tkeep,
    output [M_AXIS_OARG_49_DMWIDTH/8-1:0] m_axis_oarg_49_tstrb,
    output [M_AXIS_OARG_49_DMWIDTH-1:0] m_axis_oarg_49_tdata,
    input m_axis_oarg_49_tready,
    input ap_axis_oarg_49_tlast,
    input ap_axis_oarg_49_tvalid,
    input [M_AXIS_OARG_49_WIDTH/8-1:0] ap_axis_oarg_49_tkeep,
    input [M_AXIS_OARG_49_WIDTH/8-1:0] ap_axis_oarg_49_tstrb,
    input [M_AXIS_OARG_49_WIDTH-1:0] ap_axis_oarg_49_tdata,
    output ap_axis_oarg_49_tready,
    //output AXI-Stream pass-through interface 50
    input m_axis_oarg_50_aclk,
    input m_axis_oarg_50_aresetn,
    output m_axis_oarg_50_tlast,
    output m_axis_oarg_50_tvalid,
    output [M_AXIS_OARG_50_DMWIDTH/8-1:0] m_axis_oarg_50_tkeep,
    output [M_AXIS_OARG_50_DMWIDTH/8-1:0] m_axis_oarg_50_tstrb,
    output [M_AXIS_OARG_50_DMWIDTH-1:0] m_axis_oarg_50_tdata,
    input m_axis_oarg_50_tready,
    input ap_axis_oarg_50_tlast,
    input ap_axis_oarg_50_tvalid,
    input [M_AXIS_OARG_50_WIDTH/8-1:0] ap_axis_oarg_50_tkeep,
    input [M_AXIS_OARG_50_WIDTH/8-1:0] ap_axis_oarg_50_tstrb,
    input [M_AXIS_OARG_50_WIDTH-1:0] ap_axis_oarg_50_tdata,
    output ap_axis_oarg_50_tready,
    //output AXI-Stream pass-through interface 51
    input m_axis_oarg_51_aclk,
    input m_axis_oarg_51_aresetn,
    output m_axis_oarg_51_tlast,
    output m_axis_oarg_51_tvalid,
    output [M_AXIS_OARG_51_DMWIDTH/8-1:0] m_axis_oarg_51_tkeep,
    output [M_AXIS_OARG_51_DMWIDTH/8-1:0] m_axis_oarg_51_tstrb,
    output [M_AXIS_OARG_51_DMWIDTH-1:0] m_axis_oarg_51_tdata,
    input m_axis_oarg_51_tready,
    input ap_axis_oarg_51_tlast,
    input ap_axis_oarg_51_tvalid,
    input [M_AXIS_OARG_51_WIDTH/8-1:0] ap_axis_oarg_51_tkeep,
    input [M_AXIS_OARG_51_WIDTH/8-1:0] ap_axis_oarg_51_tstrb,
    input [M_AXIS_OARG_51_WIDTH-1:0] ap_axis_oarg_51_tdata,
    output ap_axis_oarg_51_tready,
    //output AXI-Stream pass-through interface 52
    input m_axis_oarg_52_aclk,
    input m_axis_oarg_52_aresetn,
    output m_axis_oarg_52_tlast,
    output m_axis_oarg_52_tvalid,
    output [M_AXIS_OARG_52_DMWIDTH/8-1:0] m_axis_oarg_52_tkeep,
    output [M_AXIS_OARG_52_DMWIDTH/8-1:0] m_axis_oarg_52_tstrb,
    output [M_AXIS_OARG_52_DMWIDTH-1:0] m_axis_oarg_52_tdata,
    input m_axis_oarg_52_tready,
    input ap_axis_oarg_52_tlast,
    input ap_axis_oarg_52_tvalid,
    input [M_AXIS_OARG_52_WIDTH/8-1:0] ap_axis_oarg_52_tkeep,
    input [M_AXIS_OARG_52_WIDTH/8-1:0] ap_axis_oarg_52_tstrb,
    input [M_AXIS_OARG_52_WIDTH-1:0] ap_axis_oarg_52_tdata,
    output ap_axis_oarg_52_tready,
    //output AXI-Stream pass-through interface 53
    input m_axis_oarg_53_aclk,
    input m_axis_oarg_53_aresetn,
    output m_axis_oarg_53_tlast,
    output m_axis_oarg_53_tvalid,
    output [M_AXIS_OARG_53_DMWIDTH/8-1:0] m_axis_oarg_53_tkeep,
    output [M_AXIS_OARG_53_DMWIDTH/8-1:0] m_axis_oarg_53_tstrb,
    output [M_AXIS_OARG_53_DMWIDTH-1:0] m_axis_oarg_53_tdata,
    input m_axis_oarg_53_tready,
    input ap_axis_oarg_53_tlast,
    input ap_axis_oarg_53_tvalid,
    input [M_AXIS_OARG_53_WIDTH/8-1:0] ap_axis_oarg_53_tkeep,
    input [M_AXIS_OARG_53_WIDTH/8-1:0] ap_axis_oarg_53_tstrb,
    input [M_AXIS_OARG_53_WIDTH-1:0] ap_axis_oarg_53_tdata,
    output ap_axis_oarg_53_tready,
    //output AXI-Stream pass-through interface 54
    input m_axis_oarg_54_aclk,
    input m_axis_oarg_54_aresetn,
    output m_axis_oarg_54_tlast,
    output m_axis_oarg_54_tvalid,
    output [M_AXIS_OARG_54_DMWIDTH/8-1:0] m_axis_oarg_54_tkeep,
    output [M_AXIS_OARG_54_DMWIDTH/8-1:0] m_axis_oarg_54_tstrb,
    output [M_AXIS_OARG_54_DMWIDTH-1:0] m_axis_oarg_54_tdata,
    input m_axis_oarg_54_tready,
    input ap_axis_oarg_54_tlast,
    input ap_axis_oarg_54_tvalid,
    input [M_AXIS_OARG_54_WIDTH/8-1:0] ap_axis_oarg_54_tkeep,
    input [M_AXIS_OARG_54_WIDTH/8-1:0] ap_axis_oarg_54_tstrb,
    input [M_AXIS_OARG_54_WIDTH-1:0] ap_axis_oarg_54_tdata,
    output ap_axis_oarg_54_tready,
    //output AXI-Stream pass-through interface 55
    input m_axis_oarg_55_aclk,
    input m_axis_oarg_55_aresetn,
    output m_axis_oarg_55_tlast,
    output m_axis_oarg_55_tvalid,
    output [M_AXIS_OARG_55_DMWIDTH/8-1:0] m_axis_oarg_55_tkeep,
    output [M_AXIS_OARG_55_DMWIDTH/8-1:0] m_axis_oarg_55_tstrb,
    output [M_AXIS_OARG_55_DMWIDTH-1:0] m_axis_oarg_55_tdata,
    input m_axis_oarg_55_tready,
    input ap_axis_oarg_55_tlast,
    input ap_axis_oarg_55_tvalid,
    input [M_AXIS_OARG_55_WIDTH/8-1:0] ap_axis_oarg_55_tkeep,
    input [M_AXIS_OARG_55_WIDTH/8-1:0] ap_axis_oarg_55_tstrb,
    input [M_AXIS_OARG_55_WIDTH-1:0] ap_axis_oarg_55_tdata,
    output ap_axis_oarg_55_tready,
    //output AXI-Stream pass-through interface 56
    input m_axis_oarg_56_aclk,
    input m_axis_oarg_56_aresetn,
    output m_axis_oarg_56_tlast,
    output m_axis_oarg_56_tvalid,
    output [M_AXIS_OARG_56_DMWIDTH/8-1:0] m_axis_oarg_56_tkeep,
    output [M_AXIS_OARG_56_DMWIDTH/8-1:0] m_axis_oarg_56_tstrb,
    output [M_AXIS_OARG_56_DMWIDTH-1:0] m_axis_oarg_56_tdata,
    input m_axis_oarg_56_tready,
    input ap_axis_oarg_56_tlast,
    input ap_axis_oarg_56_tvalid,
    input [M_AXIS_OARG_56_WIDTH/8-1:0] ap_axis_oarg_56_tkeep,
    input [M_AXIS_OARG_56_WIDTH/8-1:0] ap_axis_oarg_56_tstrb,
    input [M_AXIS_OARG_56_WIDTH-1:0] ap_axis_oarg_56_tdata,
    output ap_axis_oarg_56_tready,
    //output AXI-Stream pass-through interface 57
    input m_axis_oarg_57_aclk,
    input m_axis_oarg_57_aresetn,
    output m_axis_oarg_57_tlast,
    output m_axis_oarg_57_tvalid,
    output [M_AXIS_OARG_57_DMWIDTH/8-1:0] m_axis_oarg_57_tkeep,
    output [M_AXIS_OARG_57_DMWIDTH/8-1:0] m_axis_oarg_57_tstrb,
    output [M_AXIS_OARG_57_DMWIDTH-1:0] m_axis_oarg_57_tdata,
    input m_axis_oarg_57_tready,
    input ap_axis_oarg_57_tlast,
    input ap_axis_oarg_57_tvalid,
    input [M_AXIS_OARG_57_WIDTH/8-1:0] ap_axis_oarg_57_tkeep,
    input [M_AXIS_OARG_57_WIDTH/8-1:0] ap_axis_oarg_57_tstrb,
    input [M_AXIS_OARG_57_WIDTH-1:0] ap_axis_oarg_57_tdata,
    output ap_axis_oarg_57_tready,
    //output AXI-Stream pass-through interface 58
    input m_axis_oarg_58_aclk,
    input m_axis_oarg_58_aresetn,
    output m_axis_oarg_58_tlast,
    output m_axis_oarg_58_tvalid,
    output [M_AXIS_OARG_58_DMWIDTH/8-1:0] m_axis_oarg_58_tkeep,
    output [M_AXIS_OARG_58_DMWIDTH/8-1:0] m_axis_oarg_58_tstrb,
    output [M_AXIS_OARG_58_DMWIDTH-1:0] m_axis_oarg_58_tdata,
    input m_axis_oarg_58_tready,
    input ap_axis_oarg_58_tlast,
    input ap_axis_oarg_58_tvalid,
    input [M_AXIS_OARG_58_WIDTH/8-1:0] ap_axis_oarg_58_tkeep,
    input [M_AXIS_OARG_58_WIDTH/8-1:0] ap_axis_oarg_58_tstrb,
    input [M_AXIS_OARG_58_WIDTH-1:0] ap_axis_oarg_58_tdata,
    output ap_axis_oarg_58_tready,
    //output AXI-Stream pass-through interface 59
    input m_axis_oarg_59_aclk,
    input m_axis_oarg_59_aresetn,
    output m_axis_oarg_59_tlast,
    output m_axis_oarg_59_tvalid,
    output [M_AXIS_OARG_59_DMWIDTH/8-1:0] m_axis_oarg_59_tkeep,
    output [M_AXIS_OARG_59_DMWIDTH/8-1:0] m_axis_oarg_59_tstrb,
    output [M_AXIS_OARG_59_DMWIDTH-1:0] m_axis_oarg_59_tdata,
    input m_axis_oarg_59_tready,
    input ap_axis_oarg_59_tlast,
    input ap_axis_oarg_59_tvalid,
    input [M_AXIS_OARG_59_WIDTH/8-1:0] ap_axis_oarg_59_tkeep,
    input [M_AXIS_OARG_59_WIDTH/8-1:0] ap_axis_oarg_59_tstrb,
    input [M_AXIS_OARG_59_WIDTH-1:0] ap_axis_oarg_59_tdata,
    output ap_axis_oarg_59_tready,
    //output AXI-Stream pass-through interface 60
    input m_axis_oarg_60_aclk,
    input m_axis_oarg_60_aresetn,
    output m_axis_oarg_60_tlast,
    output m_axis_oarg_60_tvalid,
    output [M_AXIS_OARG_60_DMWIDTH/8-1:0] m_axis_oarg_60_tkeep,
    output [M_AXIS_OARG_60_DMWIDTH/8-1:0] m_axis_oarg_60_tstrb,
    output [M_AXIS_OARG_60_DMWIDTH-1:0] m_axis_oarg_60_tdata,
    input m_axis_oarg_60_tready,
    input ap_axis_oarg_60_tlast,
    input ap_axis_oarg_60_tvalid,
    input [M_AXIS_OARG_60_WIDTH/8-1:0] ap_axis_oarg_60_tkeep,
    input [M_AXIS_OARG_60_WIDTH/8-1:0] ap_axis_oarg_60_tstrb,
    input [M_AXIS_OARG_60_WIDTH-1:0] ap_axis_oarg_60_tdata,
    output ap_axis_oarg_60_tready,
    //output AXI-Stream pass-through interface 61
    input m_axis_oarg_61_aclk,
    input m_axis_oarg_61_aresetn,
    output m_axis_oarg_61_tlast,
    output m_axis_oarg_61_tvalid,
    output [M_AXIS_OARG_61_DMWIDTH/8-1:0] m_axis_oarg_61_tkeep,
    output [M_AXIS_OARG_61_DMWIDTH/8-1:0] m_axis_oarg_61_tstrb,
    output [M_AXIS_OARG_61_DMWIDTH-1:0] m_axis_oarg_61_tdata,
    input m_axis_oarg_61_tready,
    input ap_axis_oarg_61_tlast,
    input ap_axis_oarg_61_tvalid,
    input [M_AXIS_OARG_61_WIDTH/8-1:0] ap_axis_oarg_61_tkeep,
    input [M_AXIS_OARG_61_WIDTH/8-1:0] ap_axis_oarg_61_tstrb,
    input [M_AXIS_OARG_61_WIDTH-1:0] ap_axis_oarg_61_tdata,
    output ap_axis_oarg_61_tready,
    //output AXI-Stream pass-through interface 62
    input m_axis_oarg_62_aclk,
    input m_axis_oarg_62_aresetn,
    output m_axis_oarg_62_tlast,
    output m_axis_oarg_62_tvalid,
    output [M_AXIS_OARG_62_DMWIDTH/8-1:0] m_axis_oarg_62_tkeep,
    output [M_AXIS_OARG_62_DMWIDTH/8-1:0] m_axis_oarg_62_tstrb,
    output [M_AXIS_OARG_62_DMWIDTH-1:0] m_axis_oarg_62_tdata,
    input m_axis_oarg_62_tready,
    input ap_axis_oarg_62_tlast,
    input ap_axis_oarg_62_tvalid,
    input [M_AXIS_OARG_62_WIDTH/8-1:0] ap_axis_oarg_62_tkeep,
    input [M_AXIS_OARG_62_WIDTH/8-1:0] ap_axis_oarg_62_tstrb,
    input [M_AXIS_OARG_62_WIDTH-1:0] ap_axis_oarg_62_tdata,
    output ap_axis_oarg_62_tready,
    //output AXI-Stream pass-through interface 63
    input m_axis_oarg_63_aclk,
    input m_axis_oarg_63_aresetn,
    output m_axis_oarg_63_tlast,
    output m_axis_oarg_63_tvalid,
    output [M_AXIS_OARG_63_DMWIDTH/8-1:0] m_axis_oarg_63_tkeep,
    output [M_AXIS_OARG_63_DMWIDTH/8-1:0] m_axis_oarg_63_tstrb,
    output [M_AXIS_OARG_63_DMWIDTH-1:0] m_axis_oarg_63_tdata,
    input m_axis_oarg_63_tready,
    input ap_axis_oarg_63_tlast,
    input ap_axis_oarg_63_tvalid,
    input [M_AXIS_OARG_63_WIDTH/8-1:0] ap_axis_oarg_63_tkeep,
    input [M_AXIS_OARG_63_WIDTH/8-1:0] ap_axis_oarg_63_tstrb,
    input [M_AXIS_OARG_63_WIDTH-1:0] ap_axis_oarg_63_tdata,
    output ap_axis_oarg_63_tready,
    //output AXI-Stream pass-through interface 64
    input m_axis_oarg_64_aclk,
    input m_axis_oarg_64_aresetn,
    output m_axis_oarg_64_tlast,
    output m_axis_oarg_64_tvalid,
    output [M_AXIS_OARG_64_DMWIDTH/8-1:0] m_axis_oarg_64_tkeep,
    output [M_AXIS_OARG_64_DMWIDTH/8-1:0] m_axis_oarg_64_tstrb,
    output [M_AXIS_OARG_64_DMWIDTH-1:0] m_axis_oarg_64_tdata,
    input m_axis_oarg_64_tready,
    input ap_axis_oarg_64_tlast,
    input ap_axis_oarg_64_tvalid,
    input [M_AXIS_OARG_64_WIDTH/8-1:0] ap_axis_oarg_64_tkeep,
    input [M_AXIS_OARG_64_WIDTH/8-1:0] ap_axis_oarg_64_tstrb,
    input [M_AXIS_OARG_64_WIDTH-1:0] ap_axis_oarg_64_tdata,
    output ap_axis_oarg_64_tready,
    //output AXI-Stream pass-through interface 65
    input m_axis_oarg_65_aclk,
    input m_axis_oarg_65_aresetn,
    output m_axis_oarg_65_tlast,
    output m_axis_oarg_65_tvalid,
    output [M_AXIS_OARG_65_DMWIDTH/8-1:0] m_axis_oarg_65_tkeep,
    output [M_AXIS_OARG_65_DMWIDTH/8-1:0] m_axis_oarg_65_tstrb,
    output [M_AXIS_OARG_65_DMWIDTH-1:0] m_axis_oarg_65_tdata,
    input m_axis_oarg_65_tready,
    input ap_axis_oarg_65_tlast,
    input ap_axis_oarg_65_tvalid,
    input [M_AXIS_OARG_65_WIDTH/8-1:0] ap_axis_oarg_65_tkeep,
    input [M_AXIS_OARG_65_WIDTH/8-1:0] ap_axis_oarg_65_tstrb,
    input [M_AXIS_OARG_65_WIDTH-1:0] ap_axis_oarg_65_tdata,
    output ap_axis_oarg_65_tready,
    //output AXI-Stream pass-through interface 66
    input m_axis_oarg_66_aclk,
    input m_axis_oarg_66_aresetn,
    output m_axis_oarg_66_tlast,
    output m_axis_oarg_66_tvalid,
    output [M_AXIS_OARG_66_DMWIDTH/8-1:0] m_axis_oarg_66_tkeep,
    output [M_AXIS_OARG_66_DMWIDTH/8-1:0] m_axis_oarg_66_tstrb,
    output [M_AXIS_OARG_66_DMWIDTH-1:0] m_axis_oarg_66_tdata,
    input m_axis_oarg_66_tready,
    input ap_axis_oarg_66_tlast,
    input ap_axis_oarg_66_tvalid,
    input [M_AXIS_OARG_66_WIDTH/8-1:0] ap_axis_oarg_66_tkeep,
    input [M_AXIS_OARG_66_WIDTH/8-1:0] ap_axis_oarg_66_tstrb,
    input [M_AXIS_OARG_66_WIDTH-1:0] ap_axis_oarg_66_tdata,
    output ap_axis_oarg_66_tready,
    //output AXI-Stream pass-through interface 67
    input m_axis_oarg_67_aclk,
    input m_axis_oarg_67_aresetn,
    output m_axis_oarg_67_tlast,
    output m_axis_oarg_67_tvalid,
    output [M_AXIS_OARG_67_DMWIDTH/8-1:0] m_axis_oarg_67_tkeep,
    output [M_AXIS_OARG_67_DMWIDTH/8-1:0] m_axis_oarg_67_tstrb,
    output [M_AXIS_OARG_67_DMWIDTH-1:0] m_axis_oarg_67_tdata,
    input m_axis_oarg_67_tready,
    input ap_axis_oarg_67_tlast,
    input ap_axis_oarg_67_tvalid,
    input [M_AXIS_OARG_67_WIDTH/8-1:0] ap_axis_oarg_67_tkeep,
    input [M_AXIS_OARG_67_WIDTH/8-1:0] ap_axis_oarg_67_tstrb,
    input [M_AXIS_OARG_67_WIDTH-1:0] ap_axis_oarg_67_tdata,
    output ap_axis_oarg_67_tready,
    //output AXI-Stream pass-through interface 68
    input m_axis_oarg_68_aclk,
    input m_axis_oarg_68_aresetn,
    output m_axis_oarg_68_tlast,
    output m_axis_oarg_68_tvalid,
    output [M_AXIS_OARG_68_DMWIDTH/8-1:0] m_axis_oarg_68_tkeep,
    output [M_AXIS_OARG_68_DMWIDTH/8-1:0] m_axis_oarg_68_tstrb,
    output [M_AXIS_OARG_68_DMWIDTH-1:0] m_axis_oarg_68_tdata,
    input m_axis_oarg_68_tready,
    input ap_axis_oarg_68_tlast,
    input ap_axis_oarg_68_tvalid,
    input [M_AXIS_OARG_68_WIDTH/8-1:0] ap_axis_oarg_68_tkeep,
    input [M_AXIS_OARG_68_WIDTH/8-1:0] ap_axis_oarg_68_tstrb,
    input [M_AXIS_OARG_68_WIDTH-1:0] ap_axis_oarg_68_tdata,
    output ap_axis_oarg_68_tready,
    //output AXI-Stream pass-through interface 69
    input m_axis_oarg_69_aclk,
    input m_axis_oarg_69_aresetn,
    output m_axis_oarg_69_tlast,
    output m_axis_oarg_69_tvalid,
    output [M_AXIS_OARG_69_DMWIDTH/8-1:0] m_axis_oarg_69_tkeep,
    output [M_AXIS_OARG_69_DMWIDTH/8-1:0] m_axis_oarg_69_tstrb,
    output [M_AXIS_OARG_69_DMWIDTH-1:0] m_axis_oarg_69_tdata,
    input m_axis_oarg_69_tready,
    input ap_axis_oarg_69_tlast,
    input ap_axis_oarg_69_tvalid,
    input [M_AXIS_OARG_69_WIDTH/8-1:0] ap_axis_oarg_69_tkeep,
    input [M_AXIS_OARG_69_WIDTH/8-1:0] ap_axis_oarg_69_tstrb,
    input [M_AXIS_OARG_69_WIDTH-1:0] ap_axis_oarg_69_tdata,
    output ap_axis_oarg_69_tready,
    //output AXI-Stream pass-through interface 70
    input m_axis_oarg_70_aclk,
    input m_axis_oarg_70_aresetn,
    output m_axis_oarg_70_tlast,
    output m_axis_oarg_70_tvalid,
    output [M_AXIS_OARG_70_DMWIDTH/8-1:0] m_axis_oarg_70_tkeep,
    output [M_AXIS_OARG_70_DMWIDTH/8-1:0] m_axis_oarg_70_tstrb,
    output [M_AXIS_OARG_70_DMWIDTH-1:0] m_axis_oarg_70_tdata,
    input m_axis_oarg_70_tready,
    input ap_axis_oarg_70_tlast,
    input ap_axis_oarg_70_tvalid,
    input [M_AXIS_OARG_70_WIDTH/8-1:0] ap_axis_oarg_70_tkeep,
    input [M_AXIS_OARG_70_WIDTH/8-1:0] ap_axis_oarg_70_tstrb,
    input [M_AXIS_OARG_70_WIDTH-1:0] ap_axis_oarg_70_tdata,
    output ap_axis_oarg_70_tready,
    //output AXI-Stream pass-through interface 71
    input m_axis_oarg_71_aclk,
    input m_axis_oarg_71_aresetn,
    output m_axis_oarg_71_tlast,
    output m_axis_oarg_71_tvalid,
    output [M_AXIS_OARG_71_DMWIDTH/8-1:0] m_axis_oarg_71_tkeep,
    output [M_AXIS_OARG_71_DMWIDTH/8-1:0] m_axis_oarg_71_tstrb,
    output [M_AXIS_OARG_71_DMWIDTH-1:0] m_axis_oarg_71_tdata,
    input m_axis_oarg_71_tready,
    input ap_axis_oarg_71_tlast,
    input ap_axis_oarg_71_tvalid,
    input [M_AXIS_OARG_71_WIDTH/8-1:0] ap_axis_oarg_71_tkeep,
    input [M_AXIS_OARG_71_WIDTH/8-1:0] ap_axis_oarg_71_tstrb,
    input [M_AXIS_OARG_71_WIDTH-1:0] ap_axis_oarg_71_tdata,
    output ap_axis_oarg_71_tready,
    //output AXI-Stream pass-through interface 72
    input m_axis_oarg_72_aclk,
    input m_axis_oarg_72_aresetn,
    output m_axis_oarg_72_tlast,
    output m_axis_oarg_72_tvalid,
    output [M_AXIS_OARG_72_DMWIDTH/8-1:0] m_axis_oarg_72_tkeep,
    output [M_AXIS_OARG_72_DMWIDTH/8-1:0] m_axis_oarg_72_tstrb,
    output [M_AXIS_OARG_72_DMWIDTH-1:0] m_axis_oarg_72_tdata,
    input m_axis_oarg_72_tready,
    input ap_axis_oarg_72_tlast,
    input ap_axis_oarg_72_tvalid,
    input [M_AXIS_OARG_72_WIDTH/8-1:0] ap_axis_oarg_72_tkeep,
    input [M_AXIS_OARG_72_WIDTH/8-1:0] ap_axis_oarg_72_tstrb,
    input [M_AXIS_OARG_72_WIDTH-1:0] ap_axis_oarg_72_tdata,
    output ap_axis_oarg_72_tready,
    //output AXI-Stream pass-through interface 73
    input m_axis_oarg_73_aclk,
    input m_axis_oarg_73_aresetn,
    output m_axis_oarg_73_tlast,
    output m_axis_oarg_73_tvalid,
    output [M_AXIS_OARG_73_DMWIDTH/8-1:0] m_axis_oarg_73_tkeep,
    output [M_AXIS_OARG_73_DMWIDTH/8-1:0] m_axis_oarg_73_tstrb,
    output [M_AXIS_OARG_73_DMWIDTH-1:0] m_axis_oarg_73_tdata,
    input m_axis_oarg_73_tready,
    input ap_axis_oarg_73_tlast,
    input ap_axis_oarg_73_tvalid,
    input [M_AXIS_OARG_73_WIDTH/8-1:0] ap_axis_oarg_73_tkeep,
    input [M_AXIS_OARG_73_WIDTH/8-1:0] ap_axis_oarg_73_tstrb,
    input [M_AXIS_OARG_73_WIDTH-1:0] ap_axis_oarg_73_tdata,
    output ap_axis_oarg_73_tready,
    //output AXI-Stream pass-through interface 74
    input m_axis_oarg_74_aclk,
    input m_axis_oarg_74_aresetn,
    output m_axis_oarg_74_tlast,
    output m_axis_oarg_74_tvalid,
    output [M_AXIS_OARG_74_DMWIDTH/8-1:0] m_axis_oarg_74_tkeep,
    output [M_AXIS_OARG_74_DMWIDTH/8-1:0] m_axis_oarg_74_tstrb,
    output [M_AXIS_OARG_74_DMWIDTH-1:0] m_axis_oarg_74_tdata,
    input m_axis_oarg_74_tready,
    input ap_axis_oarg_74_tlast,
    input ap_axis_oarg_74_tvalid,
    input [M_AXIS_OARG_74_WIDTH/8-1:0] ap_axis_oarg_74_tkeep,
    input [M_AXIS_OARG_74_WIDTH/8-1:0] ap_axis_oarg_74_tstrb,
    input [M_AXIS_OARG_74_WIDTH-1:0] ap_axis_oarg_74_tdata,
    output ap_axis_oarg_74_tready,
    //output AXI-Stream pass-through interface 75
    input m_axis_oarg_75_aclk,
    input m_axis_oarg_75_aresetn,
    output m_axis_oarg_75_tlast,
    output m_axis_oarg_75_tvalid,
    output [M_AXIS_OARG_75_DMWIDTH/8-1:0] m_axis_oarg_75_tkeep,
    output [M_AXIS_OARG_75_DMWIDTH/8-1:0] m_axis_oarg_75_tstrb,
    output [M_AXIS_OARG_75_DMWIDTH-1:0] m_axis_oarg_75_tdata,
    input m_axis_oarg_75_tready,
    input ap_axis_oarg_75_tlast,
    input ap_axis_oarg_75_tvalid,
    input [M_AXIS_OARG_75_WIDTH/8-1:0] ap_axis_oarg_75_tkeep,
    input [M_AXIS_OARG_75_WIDTH/8-1:0] ap_axis_oarg_75_tstrb,
    input [M_AXIS_OARG_75_WIDTH-1:0] ap_axis_oarg_75_tdata,
    output ap_axis_oarg_75_tready,
    //output AXI-Stream pass-through interface 76
    input m_axis_oarg_76_aclk,
    input m_axis_oarg_76_aresetn,
    output m_axis_oarg_76_tlast,
    output m_axis_oarg_76_tvalid,
    output [M_AXIS_OARG_76_DMWIDTH/8-1:0] m_axis_oarg_76_tkeep,
    output [M_AXIS_OARG_76_DMWIDTH/8-1:0] m_axis_oarg_76_tstrb,
    output [M_AXIS_OARG_76_DMWIDTH-1:0] m_axis_oarg_76_tdata,
    input m_axis_oarg_76_tready,
    input ap_axis_oarg_76_tlast,
    input ap_axis_oarg_76_tvalid,
    input [M_AXIS_OARG_76_WIDTH/8-1:0] ap_axis_oarg_76_tkeep,
    input [M_AXIS_OARG_76_WIDTH/8-1:0] ap_axis_oarg_76_tstrb,
    input [M_AXIS_OARG_76_WIDTH-1:0] ap_axis_oarg_76_tdata,
    output ap_axis_oarg_76_tready,
    //output AXI-Stream pass-through interface 77
    input m_axis_oarg_77_aclk,
    input m_axis_oarg_77_aresetn,
    output m_axis_oarg_77_tlast,
    output m_axis_oarg_77_tvalid,
    output [M_AXIS_OARG_77_DMWIDTH/8-1:0] m_axis_oarg_77_tkeep,
    output [M_AXIS_OARG_77_DMWIDTH/8-1:0] m_axis_oarg_77_tstrb,
    output [M_AXIS_OARG_77_DMWIDTH-1:0] m_axis_oarg_77_tdata,
    input m_axis_oarg_77_tready,
    input ap_axis_oarg_77_tlast,
    input ap_axis_oarg_77_tvalid,
    input [M_AXIS_OARG_77_WIDTH/8-1:0] ap_axis_oarg_77_tkeep,
    input [M_AXIS_OARG_77_WIDTH/8-1:0] ap_axis_oarg_77_tstrb,
    input [M_AXIS_OARG_77_WIDTH-1:0] ap_axis_oarg_77_tdata,
    output ap_axis_oarg_77_tready,
    //output AXI-Stream pass-through interface 78
    input m_axis_oarg_78_aclk,
    input m_axis_oarg_78_aresetn,
    output m_axis_oarg_78_tlast,
    output m_axis_oarg_78_tvalid,
    output [M_AXIS_OARG_78_DMWIDTH/8-1:0] m_axis_oarg_78_tkeep,
    output [M_AXIS_OARG_78_DMWIDTH/8-1:0] m_axis_oarg_78_tstrb,
    output [M_AXIS_OARG_78_DMWIDTH-1:0] m_axis_oarg_78_tdata,
    input m_axis_oarg_78_tready,
    input ap_axis_oarg_78_tlast,
    input ap_axis_oarg_78_tvalid,
    input [M_AXIS_OARG_78_WIDTH/8-1:0] ap_axis_oarg_78_tkeep,
    input [M_AXIS_OARG_78_WIDTH/8-1:0] ap_axis_oarg_78_tstrb,
    input [M_AXIS_OARG_78_WIDTH-1:0] ap_axis_oarg_78_tdata,
    output ap_axis_oarg_78_tready,
    //output AXI-Stream pass-through interface 79
    input m_axis_oarg_79_aclk,
    input m_axis_oarg_79_aresetn,
    output m_axis_oarg_79_tlast,
    output m_axis_oarg_79_tvalid,
    output [M_AXIS_OARG_79_DMWIDTH/8-1:0] m_axis_oarg_79_tkeep,
    output [M_AXIS_OARG_79_DMWIDTH/8-1:0] m_axis_oarg_79_tstrb,
    output [M_AXIS_OARG_79_DMWIDTH-1:0] m_axis_oarg_79_tdata,
    input m_axis_oarg_79_tready,
    input ap_axis_oarg_79_tlast,
    input ap_axis_oarg_79_tvalid,
    input [M_AXIS_OARG_79_WIDTH/8-1:0] ap_axis_oarg_79_tkeep,
    input [M_AXIS_OARG_79_WIDTH/8-1:0] ap_axis_oarg_79_tstrb,
    input [M_AXIS_OARG_79_WIDTH-1:0] ap_axis_oarg_79_tdata,
    output ap_axis_oarg_79_tready,
    //output AXI-Stream pass-through interface 80
    input m_axis_oarg_80_aclk,
    input m_axis_oarg_80_aresetn,
    output m_axis_oarg_80_tlast,
    output m_axis_oarg_80_tvalid,
    output [M_AXIS_OARG_80_DMWIDTH/8-1:0] m_axis_oarg_80_tkeep,
    output [M_AXIS_OARG_80_DMWIDTH/8-1:0] m_axis_oarg_80_tstrb,
    output [M_AXIS_OARG_80_DMWIDTH-1:0] m_axis_oarg_80_tdata,
    input m_axis_oarg_80_tready,
    input ap_axis_oarg_80_tlast,
    input ap_axis_oarg_80_tvalid,
    input [M_AXIS_OARG_80_WIDTH/8-1:0] ap_axis_oarg_80_tkeep,
    input [M_AXIS_OARG_80_WIDTH/8-1:0] ap_axis_oarg_80_tstrb,
    input [M_AXIS_OARG_80_WIDTH-1:0] ap_axis_oarg_80_tdata,
    output ap_axis_oarg_80_tready,
    //output AXI-Stream pass-through interface 81
    input m_axis_oarg_81_aclk,
    input m_axis_oarg_81_aresetn,
    output m_axis_oarg_81_tlast,
    output m_axis_oarg_81_tvalid,
    output [M_AXIS_OARG_81_DMWIDTH/8-1:0] m_axis_oarg_81_tkeep,
    output [M_AXIS_OARG_81_DMWIDTH/8-1:0] m_axis_oarg_81_tstrb,
    output [M_AXIS_OARG_81_DMWIDTH-1:0] m_axis_oarg_81_tdata,
    input m_axis_oarg_81_tready,
    input ap_axis_oarg_81_tlast,
    input ap_axis_oarg_81_tvalid,
    input [M_AXIS_OARG_81_WIDTH/8-1:0] ap_axis_oarg_81_tkeep,
    input [M_AXIS_OARG_81_WIDTH/8-1:0] ap_axis_oarg_81_tstrb,
    input [M_AXIS_OARG_81_WIDTH-1:0] ap_axis_oarg_81_tdata,
    output ap_axis_oarg_81_tready,
    //output AXI-Stream pass-through interface 82
    input m_axis_oarg_82_aclk,
    input m_axis_oarg_82_aresetn,
    output m_axis_oarg_82_tlast,
    output m_axis_oarg_82_tvalid,
    output [M_AXIS_OARG_82_DMWIDTH/8-1:0] m_axis_oarg_82_tkeep,
    output [M_AXIS_OARG_82_DMWIDTH/8-1:0] m_axis_oarg_82_tstrb,
    output [M_AXIS_OARG_82_DMWIDTH-1:0] m_axis_oarg_82_tdata,
    input m_axis_oarg_82_tready,
    input ap_axis_oarg_82_tlast,
    input ap_axis_oarg_82_tvalid,
    input [M_AXIS_OARG_82_WIDTH/8-1:0] ap_axis_oarg_82_tkeep,
    input [M_AXIS_OARG_82_WIDTH/8-1:0] ap_axis_oarg_82_tstrb,
    input [M_AXIS_OARG_82_WIDTH-1:0] ap_axis_oarg_82_tdata,
    output ap_axis_oarg_82_tready,
    //output AXI-Stream pass-through interface 83
    input m_axis_oarg_83_aclk,
    input m_axis_oarg_83_aresetn,
    output m_axis_oarg_83_tlast,
    output m_axis_oarg_83_tvalid,
    output [M_AXIS_OARG_83_DMWIDTH/8-1:0] m_axis_oarg_83_tkeep,
    output [M_AXIS_OARG_83_DMWIDTH/8-1:0] m_axis_oarg_83_tstrb,
    output [M_AXIS_OARG_83_DMWIDTH-1:0] m_axis_oarg_83_tdata,
    input m_axis_oarg_83_tready,
    input ap_axis_oarg_83_tlast,
    input ap_axis_oarg_83_tvalid,
    input [M_AXIS_OARG_83_WIDTH/8-1:0] ap_axis_oarg_83_tkeep,
    input [M_AXIS_OARG_83_WIDTH/8-1:0] ap_axis_oarg_83_tstrb,
    input [M_AXIS_OARG_83_WIDTH-1:0] ap_axis_oarg_83_tdata,
    output ap_axis_oarg_83_tready,
    //output AXI-Stream pass-through interface 84
    input m_axis_oarg_84_aclk,
    input m_axis_oarg_84_aresetn,
    output m_axis_oarg_84_tlast,
    output m_axis_oarg_84_tvalid,
    output [M_AXIS_OARG_84_DMWIDTH/8-1:0] m_axis_oarg_84_tkeep,
    output [M_AXIS_OARG_84_DMWIDTH/8-1:0] m_axis_oarg_84_tstrb,
    output [M_AXIS_OARG_84_DMWIDTH-1:0] m_axis_oarg_84_tdata,
    input m_axis_oarg_84_tready,
    input ap_axis_oarg_84_tlast,
    input ap_axis_oarg_84_tvalid,
    input [M_AXIS_OARG_84_WIDTH/8-1:0] ap_axis_oarg_84_tkeep,
    input [M_AXIS_OARG_84_WIDTH/8-1:0] ap_axis_oarg_84_tstrb,
    input [M_AXIS_OARG_84_WIDTH-1:0] ap_axis_oarg_84_tdata,
    output ap_axis_oarg_84_tready,
    //output AXI-Stream pass-through interface 85
    input m_axis_oarg_85_aclk,
    input m_axis_oarg_85_aresetn,
    output m_axis_oarg_85_tlast,
    output m_axis_oarg_85_tvalid,
    output [M_AXIS_OARG_85_DMWIDTH/8-1:0] m_axis_oarg_85_tkeep,
    output [M_AXIS_OARG_85_DMWIDTH/8-1:0] m_axis_oarg_85_tstrb,
    output [M_AXIS_OARG_85_DMWIDTH-1:0] m_axis_oarg_85_tdata,
    input m_axis_oarg_85_tready,
    input ap_axis_oarg_85_tlast,
    input ap_axis_oarg_85_tvalid,
    input [M_AXIS_OARG_85_WIDTH/8-1:0] ap_axis_oarg_85_tkeep,
    input [M_AXIS_OARG_85_WIDTH/8-1:0] ap_axis_oarg_85_tstrb,
    input [M_AXIS_OARG_85_WIDTH-1:0] ap_axis_oarg_85_tdata,
    output ap_axis_oarg_85_tready,
    //output AXI-Stream pass-through interface 86
    input m_axis_oarg_86_aclk,
    input m_axis_oarg_86_aresetn,
    output m_axis_oarg_86_tlast,
    output m_axis_oarg_86_tvalid,
    output [M_AXIS_OARG_86_DMWIDTH/8-1:0] m_axis_oarg_86_tkeep,
    output [M_AXIS_OARG_86_DMWIDTH/8-1:0] m_axis_oarg_86_tstrb,
    output [M_AXIS_OARG_86_DMWIDTH-1:0] m_axis_oarg_86_tdata,
    input m_axis_oarg_86_tready,
    input ap_axis_oarg_86_tlast,
    input ap_axis_oarg_86_tvalid,
    input [M_AXIS_OARG_86_WIDTH/8-1:0] ap_axis_oarg_86_tkeep,
    input [M_AXIS_OARG_86_WIDTH/8-1:0] ap_axis_oarg_86_tstrb,
    input [M_AXIS_OARG_86_WIDTH-1:0] ap_axis_oarg_86_tdata,
    output ap_axis_oarg_86_tready,
    //output AXI-Stream pass-through interface 87
    input m_axis_oarg_87_aclk,
    input m_axis_oarg_87_aresetn,
    output m_axis_oarg_87_tlast,
    output m_axis_oarg_87_tvalid,
    output [M_AXIS_OARG_87_DMWIDTH/8-1:0] m_axis_oarg_87_tkeep,
    output [M_AXIS_OARG_87_DMWIDTH/8-1:0] m_axis_oarg_87_tstrb,
    output [M_AXIS_OARG_87_DMWIDTH-1:0] m_axis_oarg_87_tdata,
    input m_axis_oarg_87_tready,
    input ap_axis_oarg_87_tlast,
    input ap_axis_oarg_87_tvalid,
    input [M_AXIS_OARG_87_WIDTH/8-1:0] ap_axis_oarg_87_tkeep,
    input [M_AXIS_OARG_87_WIDTH/8-1:0] ap_axis_oarg_87_tstrb,
    input [M_AXIS_OARG_87_WIDTH-1:0] ap_axis_oarg_87_tdata,
    output ap_axis_oarg_87_tready,
    //output AXI-Stream pass-through interface 88
    input m_axis_oarg_88_aclk,
    input m_axis_oarg_88_aresetn,
    output m_axis_oarg_88_tlast,
    output m_axis_oarg_88_tvalid,
    output [M_AXIS_OARG_88_DMWIDTH/8-1:0] m_axis_oarg_88_tkeep,
    output [M_AXIS_OARG_88_DMWIDTH/8-1:0] m_axis_oarg_88_tstrb,
    output [M_AXIS_OARG_88_DMWIDTH-1:0] m_axis_oarg_88_tdata,
    input m_axis_oarg_88_tready,
    input ap_axis_oarg_88_tlast,
    input ap_axis_oarg_88_tvalid,
    input [M_AXIS_OARG_88_WIDTH/8-1:0] ap_axis_oarg_88_tkeep,
    input [M_AXIS_OARG_88_WIDTH/8-1:0] ap_axis_oarg_88_tstrb,
    input [M_AXIS_OARG_88_WIDTH-1:0] ap_axis_oarg_88_tdata,
    output ap_axis_oarg_88_tready,
    //output AXI-Stream pass-through interface 89
    input m_axis_oarg_89_aclk,
    input m_axis_oarg_89_aresetn,
    output m_axis_oarg_89_tlast,
    output m_axis_oarg_89_tvalid,
    output [M_AXIS_OARG_89_DMWIDTH/8-1:0] m_axis_oarg_89_tkeep,
    output [M_AXIS_OARG_89_DMWIDTH/8-1:0] m_axis_oarg_89_tstrb,
    output [M_AXIS_OARG_89_DMWIDTH-1:0] m_axis_oarg_89_tdata,
    input m_axis_oarg_89_tready,
    input ap_axis_oarg_89_tlast,
    input ap_axis_oarg_89_tvalid,
    input [M_AXIS_OARG_89_WIDTH/8-1:0] ap_axis_oarg_89_tkeep,
    input [M_AXIS_OARG_89_WIDTH/8-1:0] ap_axis_oarg_89_tstrb,
    input [M_AXIS_OARG_89_WIDTH-1:0] ap_axis_oarg_89_tdata,
    output ap_axis_oarg_89_tready,
    //output AXI-Stream pass-through interface 90
    input m_axis_oarg_90_aclk,
    input m_axis_oarg_90_aresetn,
    output m_axis_oarg_90_tlast,
    output m_axis_oarg_90_tvalid,
    output [M_AXIS_OARG_90_DMWIDTH/8-1:0] m_axis_oarg_90_tkeep,
    output [M_AXIS_OARG_90_DMWIDTH/8-1:0] m_axis_oarg_90_tstrb,
    output [M_AXIS_OARG_90_DMWIDTH-1:0] m_axis_oarg_90_tdata,
    input m_axis_oarg_90_tready,
    input ap_axis_oarg_90_tlast,
    input ap_axis_oarg_90_tvalid,
    input [M_AXIS_OARG_90_WIDTH/8-1:0] ap_axis_oarg_90_tkeep,
    input [M_AXIS_OARG_90_WIDTH/8-1:0] ap_axis_oarg_90_tstrb,
    input [M_AXIS_OARG_90_WIDTH-1:0] ap_axis_oarg_90_tdata,
    output ap_axis_oarg_90_tready,
    //output AXI-Stream pass-through interface 91
    input m_axis_oarg_91_aclk,
    input m_axis_oarg_91_aresetn,
    output m_axis_oarg_91_tlast,
    output m_axis_oarg_91_tvalid,
    output [M_AXIS_OARG_91_DMWIDTH/8-1:0] m_axis_oarg_91_tkeep,
    output [M_AXIS_OARG_91_DMWIDTH/8-1:0] m_axis_oarg_91_tstrb,
    output [M_AXIS_OARG_91_DMWIDTH-1:0] m_axis_oarg_91_tdata,
    input m_axis_oarg_91_tready,
    input ap_axis_oarg_91_tlast,
    input ap_axis_oarg_91_tvalid,
    input [M_AXIS_OARG_91_WIDTH/8-1:0] ap_axis_oarg_91_tkeep,
    input [M_AXIS_OARG_91_WIDTH/8-1:0] ap_axis_oarg_91_tstrb,
    input [M_AXIS_OARG_91_WIDTH-1:0] ap_axis_oarg_91_tdata,
    output ap_axis_oarg_91_tready,
    //output AXI-Stream pass-through interface 92
    input m_axis_oarg_92_aclk,
    input m_axis_oarg_92_aresetn,
    output m_axis_oarg_92_tlast,
    output m_axis_oarg_92_tvalid,
    output [M_AXIS_OARG_92_DMWIDTH/8-1:0] m_axis_oarg_92_tkeep,
    output [M_AXIS_OARG_92_DMWIDTH/8-1:0] m_axis_oarg_92_tstrb,
    output [M_AXIS_OARG_92_DMWIDTH-1:0] m_axis_oarg_92_tdata,
    input m_axis_oarg_92_tready,
    input ap_axis_oarg_92_tlast,
    input ap_axis_oarg_92_tvalid,
    input [M_AXIS_OARG_92_WIDTH/8-1:0] ap_axis_oarg_92_tkeep,
    input [M_AXIS_OARG_92_WIDTH/8-1:0] ap_axis_oarg_92_tstrb,
    input [M_AXIS_OARG_92_WIDTH-1:0] ap_axis_oarg_92_tdata,
    output ap_axis_oarg_92_tready,
    //output AXI-Stream pass-through interface 93
    input m_axis_oarg_93_aclk,
    input m_axis_oarg_93_aresetn,
    output m_axis_oarg_93_tlast,
    output m_axis_oarg_93_tvalid,
    output [M_AXIS_OARG_93_DMWIDTH/8-1:0] m_axis_oarg_93_tkeep,
    output [M_AXIS_OARG_93_DMWIDTH/8-1:0] m_axis_oarg_93_tstrb,
    output [M_AXIS_OARG_93_DMWIDTH-1:0] m_axis_oarg_93_tdata,
    input m_axis_oarg_93_tready,
    input ap_axis_oarg_93_tlast,
    input ap_axis_oarg_93_tvalid,
    input [M_AXIS_OARG_93_WIDTH/8-1:0] ap_axis_oarg_93_tkeep,
    input [M_AXIS_OARG_93_WIDTH/8-1:0] ap_axis_oarg_93_tstrb,
    input [M_AXIS_OARG_93_WIDTH-1:0] ap_axis_oarg_93_tdata,
    output ap_axis_oarg_93_tready,
    //output AXI-Stream pass-through interface 94
    input m_axis_oarg_94_aclk,
    input m_axis_oarg_94_aresetn,
    output m_axis_oarg_94_tlast,
    output m_axis_oarg_94_tvalid,
    output [M_AXIS_OARG_94_DMWIDTH/8-1:0] m_axis_oarg_94_tkeep,
    output [M_AXIS_OARG_94_DMWIDTH/8-1:0] m_axis_oarg_94_tstrb,
    output [M_AXIS_OARG_94_DMWIDTH-1:0] m_axis_oarg_94_tdata,
    input m_axis_oarg_94_tready,
    input ap_axis_oarg_94_tlast,
    input ap_axis_oarg_94_tvalid,
    input [M_AXIS_OARG_94_WIDTH/8-1:0] ap_axis_oarg_94_tkeep,
    input [M_AXIS_OARG_94_WIDTH/8-1:0] ap_axis_oarg_94_tstrb,
    input [M_AXIS_OARG_94_WIDTH-1:0] ap_axis_oarg_94_tdata,
    output ap_axis_oarg_94_tready,
    //output AXI-Stream pass-through interface 95
    input m_axis_oarg_95_aclk,
    input m_axis_oarg_95_aresetn,
    output m_axis_oarg_95_tlast,
    output m_axis_oarg_95_tvalid,
    output [M_AXIS_OARG_95_DMWIDTH/8-1:0] m_axis_oarg_95_tkeep,
    output [M_AXIS_OARG_95_DMWIDTH/8-1:0] m_axis_oarg_95_tstrb,
    output [M_AXIS_OARG_95_DMWIDTH-1:0] m_axis_oarg_95_tdata,
    input m_axis_oarg_95_tready,
    input ap_axis_oarg_95_tlast,
    input ap_axis_oarg_95_tvalid,
    input [M_AXIS_OARG_95_WIDTH/8-1:0] ap_axis_oarg_95_tkeep,
    input [M_AXIS_OARG_95_WIDTH/8-1:0] ap_axis_oarg_95_tstrb,
    input [M_AXIS_OARG_95_WIDTH-1:0] ap_axis_oarg_95_tdata,
    output ap_axis_oarg_95_tready,
    //output AXI-Stream pass-through interface 96
    input m_axis_oarg_96_aclk,
    input m_axis_oarg_96_aresetn,
    output m_axis_oarg_96_tlast,
    output m_axis_oarg_96_tvalid,
    output [M_AXIS_OARG_96_DMWIDTH/8-1:0] m_axis_oarg_96_tkeep,
    output [M_AXIS_OARG_96_DMWIDTH/8-1:0] m_axis_oarg_96_tstrb,
    output [M_AXIS_OARG_96_DMWIDTH-1:0] m_axis_oarg_96_tdata,
    input m_axis_oarg_96_tready,
    input ap_axis_oarg_96_tlast,
    input ap_axis_oarg_96_tvalid,
    input [M_AXIS_OARG_96_WIDTH/8-1:0] ap_axis_oarg_96_tkeep,
    input [M_AXIS_OARG_96_WIDTH/8-1:0] ap_axis_oarg_96_tstrb,
    input [M_AXIS_OARG_96_WIDTH-1:0] ap_axis_oarg_96_tdata,
    output ap_axis_oarg_96_tready,
    //output AXI-Stream pass-through interface 97
    input m_axis_oarg_97_aclk,
    input m_axis_oarg_97_aresetn,
    output m_axis_oarg_97_tlast,
    output m_axis_oarg_97_tvalid,
    output [M_AXIS_OARG_97_DMWIDTH/8-1:0] m_axis_oarg_97_tkeep,
    output [M_AXIS_OARG_97_DMWIDTH/8-1:0] m_axis_oarg_97_tstrb,
    output [M_AXIS_OARG_97_DMWIDTH-1:0] m_axis_oarg_97_tdata,
    input m_axis_oarg_97_tready,
    input ap_axis_oarg_97_tlast,
    input ap_axis_oarg_97_tvalid,
    input [M_AXIS_OARG_97_WIDTH/8-1:0] ap_axis_oarg_97_tkeep,
    input [M_AXIS_OARG_97_WIDTH/8-1:0] ap_axis_oarg_97_tstrb,
    input [M_AXIS_OARG_97_WIDTH-1:0] ap_axis_oarg_97_tdata,
    output ap_axis_oarg_97_tready,
    //output AXI-Stream pass-through interface 98
    input m_axis_oarg_98_aclk,
    input m_axis_oarg_98_aresetn,
    output m_axis_oarg_98_tlast,
    output m_axis_oarg_98_tvalid,
    output [M_AXIS_OARG_98_DMWIDTH/8-1:0] m_axis_oarg_98_tkeep,
    output [M_AXIS_OARG_98_DMWIDTH/8-1:0] m_axis_oarg_98_tstrb,
    output [M_AXIS_OARG_98_DMWIDTH-1:0] m_axis_oarg_98_tdata,
    input m_axis_oarg_98_tready,
    input ap_axis_oarg_98_tlast,
    input ap_axis_oarg_98_tvalid,
    input [M_AXIS_OARG_98_WIDTH/8-1:0] ap_axis_oarg_98_tkeep,
    input [M_AXIS_OARG_98_WIDTH/8-1:0] ap_axis_oarg_98_tstrb,
    input [M_AXIS_OARG_98_WIDTH-1:0] ap_axis_oarg_98_tdata,
    output ap_axis_oarg_98_tready,
    //output AXI-Stream pass-through interface 99
    input m_axis_oarg_99_aclk,
    input m_axis_oarg_99_aresetn,
    output m_axis_oarg_99_tlast,
    output m_axis_oarg_99_tvalid,
    output [M_AXIS_OARG_99_DMWIDTH/8-1:0] m_axis_oarg_99_tkeep,
    output [M_AXIS_OARG_99_DMWIDTH/8-1:0] m_axis_oarg_99_tstrb,
    output [M_AXIS_OARG_99_DMWIDTH-1:0] m_axis_oarg_99_tdata,
    input m_axis_oarg_99_tready,
    input ap_axis_oarg_99_tlast,
    input ap_axis_oarg_99_tvalid,
    input [M_AXIS_OARG_99_WIDTH/8-1:0] ap_axis_oarg_99_tkeep,
    input [M_AXIS_OARG_99_WIDTH/8-1:0] ap_axis_oarg_99_tstrb,
    input [M_AXIS_OARG_99_WIDTH-1:0] ap_axis_oarg_99_tdata,
    output ap_axis_oarg_99_tready,
    //output AXI-Stream pass-through interface 100
    input m_axis_oarg_100_aclk,
    input m_axis_oarg_100_aresetn,
    output m_axis_oarg_100_tlast,
    output m_axis_oarg_100_tvalid,
    output [M_AXIS_OARG_100_DMWIDTH/8-1:0] m_axis_oarg_100_tkeep,
    output [M_AXIS_OARG_100_DMWIDTH/8-1:0] m_axis_oarg_100_tstrb,
    output [M_AXIS_OARG_100_DMWIDTH-1:0] m_axis_oarg_100_tdata,
    input m_axis_oarg_100_tready,
    input ap_axis_oarg_100_tlast,
    input ap_axis_oarg_100_tvalid,
    input [M_AXIS_OARG_100_WIDTH/8-1:0] ap_axis_oarg_100_tkeep,
    input [M_AXIS_OARG_100_WIDTH/8-1:0] ap_axis_oarg_100_tstrb,
    input [M_AXIS_OARG_100_WIDTH-1:0] ap_axis_oarg_100_tdata,
    output ap_axis_oarg_100_tready,
    //output AXI-Stream pass-through interface 101
    input m_axis_oarg_101_aclk,
    input m_axis_oarg_101_aresetn,
    output m_axis_oarg_101_tlast,
    output m_axis_oarg_101_tvalid,
    output [M_AXIS_OARG_101_DMWIDTH/8-1:0] m_axis_oarg_101_tkeep,
    output [M_AXIS_OARG_101_DMWIDTH/8-1:0] m_axis_oarg_101_tstrb,
    output [M_AXIS_OARG_101_DMWIDTH-1:0] m_axis_oarg_101_tdata,
    input m_axis_oarg_101_tready,
    input ap_axis_oarg_101_tlast,
    input ap_axis_oarg_101_tvalid,
    input [M_AXIS_OARG_101_WIDTH/8-1:0] ap_axis_oarg_101_tkeep,
    input [M_AXIS_OARG_101_WIDTH/8-1:0] ap_axis_oarg_101_tstrb,
    input [M_AXIS_OARG_101_WIDTH-1:0] ap_axis_oarg_101_tdata,
    output ap_axis_oarg_101_tready,
    //output AXI-Stream pass-through interface 102
    input m_axis_oarg_102_aclk,
    input m_axis_oarg_102_aresetn,
    output m_axis_oarg_102_tlast,
    output m_axis_oarg_102_tvalid,
    output [M_AXIS_OARG_102_DMWIDTH/8-1:0] m_axis_oarg_102_tkeep,
    output [M_AXIS_OARG_102_DMWIDTH/8-1:0] m_axis_oarg_102_tstrb,
    output [M_AXIS_OARG_102_DMWIDTH-1:0] m_axis_oarg_102_tdata,
    input m_axis_oarg_102_tready,
    input ap_axis_oarg_102_tlast,
    input ap_axis_oarg_102_tvalid,
    input [M_AXIS_OARG_102_WIDTH/8-1:0] ap_axis_oarg_102_tkeep,
    input [M_AXIS_OARG_102_WIDTH/8-1:0] ap_axis_oarg_102_tstrb,
    input [M_AXIS_OARG_102_WIDTH-1:0] ap_axis_oarg_102_tdata,
    output ap_axis_oarg_102_tready,
    //output AXI-Stream pass-through interface 103
    input m_axis_oarg_103_aclk,
    input m_axis_oarg_103_aresetn,
    output m_axis_oarg_103_tlast,
    output m_axis_oarg_103_tvalid,
    output [M_AXIS_OARG_103_DMWIDTH/8-1:0] m_axis_oarg_103_tkeep,
    output [M_AXIS_OARG_103_DMWIDTH/8-1:0] m_axis_oarg_103_tstrb,
    output [M_AXIS_OARG_103_DMWIDTH-1:0] m_axis_oarg_103_tdata,
    input m_axis_oarg_103_tready,
    input ap_axis_oarg_103_tlast,
    input ap_axis_oarg_103_tvalid,
    input [M_AXIS_OARG_103_WIDTH/8-1:0] ap_axis_oarg_103_tkeep,
    input [M_AXIS_OARG_103_WIDTH/8-1:0] ap_axis_oarg_103_tstrb,
    input [M_AXIS_OARG_103_WIDTH-1:0] ap_axis_oarg_103_tdata,
    output ap_axis_oarg_103_tready,
    //output AXI-Stream pass-through interface 104
    input m_axis_oarg_104_aclk,
    input m_axis_oarg_104_aresetn,
    output m_axis_oarg_104_tlast,
    output m_axis_oarg_104_tvalid,
    output [M_AXIS_OARG_104_DMWIDTH/8-1:0] m_axis_oarg_104_tkeep,
    output [M_AXIS_OARG_104_DMWIDTH/8-1:0] m_axis_oarg_104_tstrb,
    output [M_AXIS_OARG_104_DMWIDTH-1:0] m_axis_oarg_104_tdata,
    input m_axis_oarg_104_tready,
    input ap_axis_oarg_104_tlast,
    input ap_axis_oarg_104_tvalid,
    input [M_AXIS_OARG_104_WIDTH/8-1:0] ap_axis_oarg_104_tkeep,
    input [M_AXIS_OARG_104_WIDTH/8-1:0] ap_axis_oarg_104_tstrb,
    input [M_AXIS_OARG_104_WIDTH-1:0] ap_axis_oarg_104_tdata,
    output ap_axis_oarg_104_tready,
    //output AXI-Stream pass-through interface 105
    input m_axis_oarg_105_aclk,
    input m_axis_oarg_105_aresetn,
    output m_axis_oarg_105_tlast,
    output m_axis_oarg_105_tvalid,
    output [M_AXIS_OARG_105_DMWIDTH/8-1:0] m_axis_oarg_105_tkeep,
    output [M_AXIS_OARG_105_DMWIDTH/8-1:0] m_axis_oarg_105_tstrb,
    output [M_AXIS_OARG_105_DMWIDTH-1:0] m_axis_oarg_105_tdata,
    input m_axis_oarg_105_tready,
    input ap_axis_oarg_105_tlast,
    input ap_axis_oarg_105_tvalid,
    input [M_AXIS_OARG_105_WIDTH/8-1:0] ap_axis_oarg_105_tkeep,
    input [M_AXIS_OARG_105_WIDTH/8-1:0] ap_axis_oarg_105_tstrb,
    input [M_AXIS_OARG_105_WIDTH-1:0] ap_axis_oarg_105_tdata,
    output ap_axis_oarg_105_tready,
    //output AXI-Stream pass-through interface 106
    input m_axis_oarg_106_aclk,
    input m_axis_oarg_106_aresetn,
    output m_axis_oarg_106_tlast,
    output m_axis_oarg_106_tvalid,
    output [M_AXIS_OARG_106_DMWIDTH/8-1:0] m_axis_oarg_106_tkeep,
    output [M_AXIS_OARG_106_DMWIDTH/8-1:0] m_axis_oarg_106_tstrb,
    output [M_AXIS_OARG_106_DMWIDTH-1:0] m_axis_oarg_106_tdata,
    input m_axis_oarg_106_tready,
    input ap_axis_oarg_106_tlast,
    input ap_axis_oarg_106_tvalid,
    input [M_AXIS_OARG_106_WIDTH/8-1:0] ap_axis_oarg_106_tkeep,
    input [M_AXIS_OARG_106_WIDTH/8-1:0] ap_axis_oarg_106_tstrb,
    input [M_AXIS_OARG_106_WIDTH-1:0] ap_axis_oarg_106_tdata,
    output ap_axis_oarg_106_tready,
    //output AXI-Stream pass-through interface 107
    input m_axis_oarg_107_aclk,
    input m_axis_oarg_107_aresetn,
    output m_axis_oarg_107_tlast,
    output m_axis_oarg_107_tvalid,
    output [M_AXIS_OARG_107_DMWIDTH/8-1:0] m_axis_oarg_107_tkeep,
    output [M_AXIS_OARG_107_DMWIDTH/8-1:0] m_axis_oarg_107_tstrb,
    output [M_AXIS_OARG_107_DMWIDTH-1:0] m_axis_oarg_107_tdata,
    input m_axis_oarg_107_tready,
    input ap_axis_oarg_107_tlast,
    input ap_axis_oarg_107_tvalid,
    input [M_AXIS_OARG_107_WIDTH/8-1:0] ap_axis_oarg_107_tkeep,
    input [M_AXIS_OARG_107_WIDTH/8-1:0] ap_axis_oarg_107_tstrb,
    input [M_AXIS_OARG_107_WIDTH-1:0] ap_axis_oarg_107_tdata,
    output ap_axis_oarg_107_tready,
    //output AXI-Stream pass-through interface 108
    input m_axis_oarg_108_aclk,
    input m_axis_oarg_108_aresetn,
    output m_axis_oarg_108_tlast,
    output m_axis_oarg_108_tvalid,
    output [M_AXIS_OARG_108_DMWIDTH/8-1:0] m_axis_oarg_108_tkeep,
    output [M_AXIS_OARG_108_DMWIDTH/8-1:0] m_axis_oarg_108_tstrb,
    output [M_AXIS_OARG_108_DMWIDTH-1:0] m_axis_oarg_108_tdata,
    input m_axis_oarg_108_tready,
    input ap_axis_oarg_108_tlast,
    input ap_axis_oarg_108_tvalid,
    input [M_AXIS_OARG_108_WIDTH/8-1:0] ap_axis_oarg_108_tkeep,
    input [M_AXIS_OARG_108_WIDTH/8-1:0] ap_axis_oarg_108_tstrb,
    input [M_AXIS_OARG_108_WIDTH-1:0] ap_axis_oarg_108_tdata,
    output ap_axis_oarg_108_tready,
    //output AXI-Stream pass-through interface 109
    input m_axis_oarg_109_aclk,
    input m_axis_oarg_109_aresetn,
    output m_axis_oarg_109_tlast,
    output m_axis_oarg_109_tvalid,
    output [M_AXIS_OARG_109_DMWIDTH/8-1:0] m_axis_oarg_109_tkeep,
    output [M_AXIS_OARG_109_DMWIDTH/8-1:0] m_axis_oarg_109_tstrb,
    output [M_AXIS_OARG_109_DMWIDTH-1:0] m_axis_oarg_109_tdata,
    input m_axis_oarg_109_tready,
    input ap_axis_oarg_109_tlast,
    input ap_axis_oarg_109_tvalid,
    input [M_AXIS_OARG_109_WIDTH/8-1:0] ap_axis_oarg_109_tkeep,
    input [M_AXIS_OARG_109_WIDTH/8-1:0] ap_axis_oarg_109_tstrb,
    input [M_AXIS_OARG_109_WIDTH-1:0] ap_axis_oarg_109_tdata,
    output ap_axis_oarg_109_tready,
    //output AXI-Stream pass-through interface 110
    input m_axis_oarg_110_aclk,
    input m_axis_oarg_110_aresetn,
    output m_axis_oarg_110_tlast,
    output m_axis_oarg_110_tvalid,
    output [M_AXIS_OARG_110_DMWIDTH/8-1:0] m_axis_oarg_110_tkeep,
    output [M_AXIS_OARG_110_DMWIDTH/8-1:0] m_axis_oarg_110_tstrb,
    output [M_AXIS_OARG_110_DMWIDTH-1:0] m_axis_oarg_110_tdata,
    input m_axis_oarg_110_tready,
    input ap_axis_oarg_110_tlast,
    input ap_axis_oarg_110_tvalid,
    input [M_AXIS_OARG_110_WIDTH/8-1:0] ap_axis_oarg_110_tkeep,
    input [M_AXIS_OARG_110_WIDTH/8-1:0] ap_axis_oarg_110_tstrb,
    input [M_AXIS_OARG_110_WIDTH-1:0] ap_axis_oarg_110_tdata,
    output ap_axis_oarg_110_tready,
    //output AXI-Stream pass-through interface 111
    input m_axis_oarg_111_aclk,
    input m_axis_oarg_111_aresetn,
    output m_axis_oarg_111_tlast,
    output m_axis_oarg_111_tvalid,
    output [M_AXIS_OARG_111_DMWIDTH/8-1:0] m_axis_oarg_111_tkeep,
    output [M_AXIS_OARG_111_DMWIDTH/8-1:0] m_axis_oarg_111_tstrb,
    output [M_AXIS_OARG_111_DMWIDTH-1:0] m_axis_oarg_111_tdata,
    input m_axis_oarg_111_tready,
    input ap_axis_oarg_111_tlast,
    input ap_axis_oarg_111_tvalid,
    input [M_AXIS_OARG_111_WIDTH/8-1:0] ap_axis_oarg_111_tkeep,
    input [M_AXIS_OARG_111_WIDTH/8-1:0] ap_axis_oarg_111_tstrb,
    input [M_AXIS_OARG_111_WIDTH-1:0] ap_axis_oarg_111_tdata,
    output ap_axis_oarg_111_tready,
    //output AXI-Stream pass-through interface 112
    input m_axis_oarg_112_aclk,
    input m_axis_oarg_112_aresetn,
    output m_axis_oarg_112_tlast,
    output m_axis_oarg_112_tvalid,
    output [M_AXIS_OARG_112_DMWIDTH/8-1:0] m_axis_oarg_112_tkeep,
    output [M_AXIS_OARG_112_DMWIDTH/8-1:0] m_axis_oarg_112_tstrb,
    output [M_AXIS_OARG_112_DMWIDTH-1:0] m_axis_oarg_112_tdata,
    input m_axis_oarg_112_tready,
    input ap_axis_oarg_112_tlast,
    input ap_axis_oarg_112_tvalid,
    input [M_AXIS_OARG_112_WIDTH/8-1:0] ap_axis_oarg_112_tkeep,
    input [M_AXIS_OARG_112_WIDTH/8-1:0] ap_axis_oarg_112_tstrb,
    input [M_AXIS_OARG_112_WIDTH-1:0] ap_axis_oarg_112_tdata,
    output ap_axis_oarg_112_tready,
    //output AXI-Stream pass-through interface 113
    input m_axis_oarg_113_aclk,
    input m_axis_oarg_113_aresetn,
    output m_axis_oarg_113_tlast,
    output m_axis_oarg_113_tvalid,
    output [M_AXIS_OARG_113_DMWIDTH/8-1:0] m_axis_oarg_113_tkeep,
    output [M_AXIS_OARG_113_DMWIDTH/8-1:0] m_axis_oarg_113_tstrb,
    output [M_AXIS_OARG_113_DMWIDTH-1:0] m_axis_oarg_113_tdata,
    input m_axis_oarg_113_tready,
    input ap_axis_oarg_113_tlast,
    input ap_axis_oarg_113_tvalid,
    input [M_AXIS_OARG_113_WIDTH/8-1:0] ap_axis_oarg_113_tkeep,
    input [M_AXIS_OARG_113_WIDTH/8-1:0] ap_axis_oarg_113_tstrb,
    input [M_AXIS_OARG_113_WIDTH-1:0] ap_axis_oarg_113_tdata,
    output ap_axis_oarg_113_tready,
    //output AXI-Stream pass-through interface 114
    input m_axis_oarg_114_aclk,
    input m_axis_oarg_114_aresetn,
    output m_axis_oarg_114_tlast,
    output m_axis_oarg_114_tvalid,
    output [M_AXIS_OARG_114_DMWIDTH/8-1:0] m_axis_oarg_114_tkeep,
    output [M_AXIS_OARG_114_DMWIDTH/8-1:0] m_axis_oarg_114_tstrb,
    output [M_AXIS_OARG_114_DMWIDTH-1:0] m_axis_oarg_114_tdata,
    input m_axis_oarg_114_tready,
    input ap_axis_oarg_114_tlast,
    input ap_axis_oarg_114_tvalid,
    input [M_AXIS_OARG_114_WIDTH/8-1:0] ap_axis_oarg_114_tkeep,
    input [M_AXIS_OARG_114_WIDTH/8-1:0] ap_axis_oarg_114_tstrb,
    input [M_AXIS_OARG_114_WIDTH-1:0] ap_axis_oarg_114_tdata,
    output ap_axis_oarg_114_tready,
    //output AXI-Stream pass-through interface 115
    input m_axis_oarg_115_aclk,
    input m_axis_oarg_115_aresetn,
    output m_axis_oarg_115_tlast,
    output m_axis_oarg_115_tvalid,
    output [M_AXIS_OARG_115_DMWIDTH/8-1:0] m_axis_oarg_115_tkeep,
    output [M_AXIS_OARG_115_DMWIDTH/8-1:0] m_axis_oarg_115_tstrb,
    output [M_AXIS_OARG_115_DMWIDTH-1:0] m_axis_oarg_115_tdata,
    input m_axis_oarg_115_tready,
    input ap_axis_oarg_115_tlast,
    input ap_axis_oarg_115_tvalid,
    input [M_AXIS_OARG_115_WIDTH/8-1:0] ap_axis_oarg_115_tkeep,
    input [M_AXIS_OARG_115_WIDTH/8-1:0] ap_axis_oarg_115_tstrb,
    input [M_AXIS_OARG_115_WIDTH-1:0] ap_axis_oarg_115_tdata,
    output ap_axis_oarg_115_tready,
    //output AXI-Stream pass-through interface 116
    input m_axis_oarg_116_aclk,
    input m_axis_oarg_116_aresetn,
    output m_axis_oarg_116_tlast,
    output m_axis_oarg_116_tvalid,
    output [M_AXIS_OARG_116_DMWIDTH/8-1:0] m_axis_oarg_116_tkeep,
    output [M_AXIS_OARG_116_DMWIDTH/8-1:0] m_axis_oarg_116_tstrb,
    output [M_AXIS_OARG_116_DMWIDTH-1:0] m_axis_oarg_116_tdata,
    input m_axis_oarg_116_tready,
    input ap_axis_oarg_116_tlast,
    input ap_axis_oarg_116_tvalid,
    input [M_AXIS_OARG_116_WIDTH/8-1:0] ap_axis_oarg_116_tkeep,
    input [M_AXIS_OARG_116_WIDTH/8-1:0] ap_axis_oarg_116_tstrb,
    input [M_AXIS_OARG_116_WIDTH-1:0] ap_axis_oarg_116_tdata,
    output ap_axis_oarg_116_tready,
    //output AXI-Stream pass-through interface 117
    input m_axis_oarg_117_aclk,
    input m_axis_oarg_117_aresetn,
    output m_axis_oarg_117_tlast,
    output m_axis_oarg_117_tvalid,
    output [M_AXIS_OARG_117_DMWIDTH/8-1:0] m_axis_oarg_117_tkeep,
    output [M_AXIS_OARG_117_DMWIDTH/8-1:0] m_axis_oarg_117_tstrb,
    output [M_AXIS_OARG_117_DMWIDTH-1:0] m_axis_oarg_117_tdata,
    input m_axis_oarg_117_tready,
    input ap_axis_oarg_117_tlast,
    input ap_axis_oarg_117_tvalid,
    input [M_AXIS_OARG_117_WIDTH/8-1:0] ap_axis_oarg_117_tkeep,
    input [M_AXIS_OARG_117_WIDTH/8-1:0] ap_axis_oarg_117_tstrb,
    input [M_AXIS_OARG_117_WIDTH-1:0] ap_axis_oarg_117_tdata,
    output ap_axis_oarg_117_tready,
    //output AXI-Stream pass-through interface 118
    input m_axis_oarg_118_aclk,
    input m_axis_oarg_118_aresetn,
    output m_axis_oarg_118_tlast,
    output m_axis_oarg_118_tvalid,
    output [M_AXIS_OARG_118_DMWIDTH/8-1:0] m_axis_oarg_118_tkeep,
    output [M_AXIS_OARG_118_DMWIDTH/8-1:0] m_axis_oarg_118_tstrb,
    output [M_AXIS_OARG_118_DMWIDTH-1:0] m_axis_oarg_118_tdata,
    input m_axis_oarg_118_tready,
    input ap_axis_oarg_118_tlast,
    input ap_axis_oarg_118_tvalid,
    input [M_AXIS_OARG_118_WIDTH/8-1:0] ap_axis_oarg_118_tkeep,
    input [M_AXIS_OARG_118_WIDTH/8-1:0] ap_axis_oarg_118_tstrb,
    input [M_AXIS_OARG_118_WIDTH-1:0] ap_axis_oarg_118_tdata,
    output ap_axis_oarg_118_tready,
    //output AXI-Stream pass-through interface 119
    input m_axis_oarg_119_aclk,
    input m_axis_oarg_119_aresetn,
    output m_axis_oarg_119_tlast,
    output m_axis_oarg_119_tvalid,
    output [M_AXIS_OARG_119_DMWIDTH/8-1:0] m_axis_oarg_119_tkeep,
    output [M_AXIS_OARG_119_DMWIDTH/8-1:0] m_axis_oarg_119_tstrb,
    output [M_AXIS_OARG_119_DMWIDTH-1:0] m_axis_oarg_119_tdata,
    input m_axis_oarg_119_tready,
    input ap_axis_oarg_119_tlast,
    input ap_axis_oarg_119_tvalid,
    input [M_AXIS_OARG_119_WIDTH/8-1:0] ap_axis_oarg_119_tkeep,
    input [M_AXIS_OARG_119_WIDTH/8-1:0] ap_axis_oarg_119_tstrb,
    input [M_AXIS_OARG_119_WIDTH-1:0] ap_axis_oarg_119_tdata,
    output ap_axis_oarg_119_tready,
    //output AXI-Stream pass-through interface 120
    input m_axis_oarg_120_aclk,
    input m_axis_oarg_120_aresetn,
    output m_axis_oarg_120_tlast,
    output m_axis_oarg_120_tvalid,
    output [M_AXIS_OARG_120_DMWIDTH/8-1:0] m_axis_oarg_120_tkeep,
    output [M_AXIS_OARG_120_DMWIDTH/8-1:0] m_axis_oarg_120_tstrb,
    output [M_AXIS_OARG_120_DMWIDTH-1:0] m_axis_oarg_120_tdata,
    input m_axis_oarg_120_tready,
    input ap_axis_oarg_120_tlast,
    input ap_axis_oarg_120_tvalid,
    input [M_AXIS_OARG_120_WIDTH/8-1:0] ap_axis_oarg_120_tkeep,
    input [M_AXIS_OARG_120_WIDTH/8-1:0] ap_axis_oarg_120_tstrb,
    input [M_AXIS_OARG_120_WIDTH-1:0] ap_axis_oarg_120_tdata,
    output ap_axis_oarg_120_tready,
    //output AXI-Stream pass-through interface 121
    input m_axis_oarg_121_aclk,
    input m_axis_oarg_121_aresetn,
    output m_axis_oarg_121_tlast,
    output m_axis_oarg_121_tvalid,
    output [M_AXIS_OARG_121_DMWIDTH/8-1:0] m_axis_oarg_121_tkeep,
    output [M_AXIS_OARG_121_DMWIDTH/8-1:0] m_axis_oarg_121_tstrb,
    output [M_AXIS_OARG_121_DMWIDTH-1:0] m_axis_oarg_121_tdata,
    input m_axis_oarg_121_tready,
    input ap_axis_oarg_121_tlast,
    input ap_axis_oarg_121_tvalid,
    input [M_AXIS_OARG_121_WIDTH/8-1:0] ap_axis_oarg_121_tkeep,
    input [M_AXIS_OARG_121_WIDTH/8-1:0] ap_axis_oarg_121_tstrb,
    input [M_AXIS_OARG_121_WIDTH-1:0] ap_axis_oarg_121_tdata,
    output ap_axis_oarg_121_tready,
    //output AXI-Stream pass-through interface 122
    input m_axis_oarg_122_aclk,
    input m_axis_oarg_122_aresetn,
    output m_axis_oarg_122_tlast,
    output m_axis_oarg_122_tvalid,
    output [M_AXIS_OARG_122_DMWIDTH/8-1:0] m_axis_oarg_122_tkeep,
    output [M_AXIS_OARG_122_DMWIDTH/8-1:0] m_axis_oarg_122_tstrb,
    output [M_AXIS_OARG_122_DMWIDTH-1:0] m_axis_oarg_122_tdata,
    input m_axis_oarg_122_tready,
    input ap_axis_oarg_122_tlast,
    input ap_axis_oarg_122_tvalid,
    input [M_AXIS_OARG_122_WIDTH/8-1:0] ap_axis_oarg_122_tkeep,
    input [M_AXIS_OARG_122_WIDTH/8-1:0] ap_axis_oarg_122_tstrb,
    input [M_AXIS_OARG_122_WIDTH-1:0] ap_axis_oarg_122_tdata,
    output ap_axis_oarg_122_tready,
    //output AXI-Stream pass-through interface 123
    input m_axis_oarg_123_aclk,
    input m_axis_oarg_123_aresetn,
    output m_axis_oarg_123_tlast,
    output m_axis_oarg_123_tvalid,
    output [M_AXIS_OARG_123_DMWIDTH/8-1:0] m_axis_oarg_123_tkeep,
    output [M_AXIS_OARG_123_DMWIDTH/8-1:0] m_axis_oarg_123_tstrb,
    output [M_AXIS_OARG_123_DMWIDTH-1:0] m_axis_oarg_123_tdata,
    input m_axis_oarg_123_tready,
    input ap_axis_oarg_123_tlast,
    input ap_axis_oarg_123_tvalid,
    input [M_AXIS_OARG_123_WIDTH/8-1:0] ap_axis_oarg_123_tkeep,
    input [M_AXIS_OARG_123_WIDTH/8-1:0] ap_axis_oarg_123_tstrb,
    input [M_AXIS_OARG_123_WIDTH-1:0] ap_axis_oarg_123_tdata,
    output ap_axis_oarg_123_tready,
    //output AXI-Stream pass-through interface 124
    input m_axis_oarg_124_aclk,
    input m_axis_oarg_124_aresetn,
    output m_axis_oarg_124_tlast,
    output m_axis_oarg_124_tvalid,
    output [M_AXIS_OARG_124_DMWIDTH/8-1:0] m_axis_oarg_124_tkeep,
    output [M_AXIS_OARG_124_DMWIDTH/8-1:0] m_axis_oarg_124_tstrb,
    output [M_AXIS_OARG_124_DMWIDTH-1:0] m_axis_oarg_124_tdata,
    input m_axis_oarg_124_tready,
    input ap_axis_oarg_124_tlast,
    input ap_axis_oarg_124_tvalid,
    input [M_AXIS_OARG_124_WIDTH/8-1:0] ap_axis_oarg_124_tkeep,
    input [M_AXIS_OARG_124_WIDTH/8-1:0] ap_axis_oarg_124_tstrb,
    input [M_AXIS_OARG_124_WIDTH-1:0] ap_axis_oarg_124_tdata,
    output ap_axis_oarg_124_tready,
    //output AXI-Stream pass-through interface 125
    input m_axis_oarg_125_aclk,
    input m_axis_oarg_125_aresetn,
    output m_axis_oarg_125_tlast,
    output m_axis_oarg_125_tvalid,
    output [M_AXIS_OARG_125_DMWIDTH/8-1:0] m_axis_oarg_125_tkeep,
    output [M_AXIS_OARG_125_DMWIDTH/8-1:0] m_axis_oarg_125_tstrb,
    output [M_AXIS_OARG_125_DMWIDTH-1:0] m_axis_oarg_125_tdata,
    input m_axis_oarg_125_tready,
    input ap_axis_oarg_125_tlast,
    input ap_axis_oarg_125_tvalid,
    input [M_AXIS_OARG_125_WIDTH/8-1:0] ap_axis_oarg_125_tkeep,
    input [M_AXIS_OARG_125_WIDTH/8-1:0] ap_axis_oarg_125_tstrb,
    input [M_AXIS_OARG_125_WIDTH-1:0] ap_axis_oarg_125_tdata,
    output ap_axis_oarg_125_tready,
    //output AXI-Stream pass-through interface 126
    input m_axis_oarg_126_aclk,
    input m_axis_oarg_126_aresetn,
    output m_axis_oarg_126_tlast,
    output m_axis_oarg_126_tvalid,
    output [M_AXIS_OARG_126_DMWIDTH/8-1:0] m_axis_oarg_126_tkeep,
    output [M_AXIS_OARG_126_DMWIDTH/8-1:0] m_axis_oarg_126_tstrb,
    output [M_AXIS_OARG_126_DMWIDTH-1:0] m_axis_oarg_126_tdata,
    input m_axis_oarg_126_tready,
    input ap_axis_oarg_126_tlast,
    input ap_axis_oarg_126_tvalid,
    input [M_AXIS_OARG_126_WIDTH/8-1:0] ap_axis_oarg_126_tkeep,
    input [M_AXIS_OARG_126_WIDTH/8-1:0] ap_axis_oarg_126_tstrb,
    input [M_AXIS_OARG_126_WIDTH-1:0] ap_axis_oarg_126_tdata,
    output ap_axis_oarg_126_tready,
    //output AXI-Stream pass-through interface 127
    input m_axis_oarg_127_aclk,
    input m_axis_oarg_127_aresetn,
    output m_axis_oarg_127_tlast,
    output m_axis_oarg_127_tvalid,
    output [M_AXIS_OARG_127_DMWIDTH/8-1:0] m_axis_oarg_127_tkeep,
    output [M_AXIS_OARG_127_DMWIDTH/8-1:0] m_axis_oarg_127_tstrb,
    output [M_AXIS_OARG_127_DMWIDTH-1:0] m_axis_oarg_127_tdata,
    input m_axis_oarg_127_tready,
    input ap_axis_oarg_127_tlast,
    input ap_axis_oarg_127_tvalid,
    input [M_AXIS_OARG_127_WIDTH/8-1:0] ap_axis_oarg_127_tkeep,
    input [M_AXIS_OARG_127_WIDTH/8-1:0] ap_axis_oarg_127_tstrb,
    input [M_AXIS_OARG_127_WIDTH-1:0] ap_axis_oarg_127_tdata,
    output ap_axis_oarg_127_tready,
    //-----------------------------------------------------
    //AXI-MM pass-through interface 0
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_0_AWADDR,
    input wire [7:0]                      AP_AXIMM_0_AWLEN,
    input wire [2:0]                      AP_AXIMM_0_AWSIZE,
    input wire [1:0]                      AP_AXIMM_0_AWBURST,
    input wire [1:0]                      AP_AXIMM_0_AWLOCK,
    input wire [3:0]                      AP_AXIMM_0_AWCACHE,
    input wire [2:0]                      AP_AXIMM_0_AWPROT,
    input wire [3:0]                      AP_AXIMM_0_AWREGION,
    input wire [3:0]                      AP_AXIMM_0_AWQOS,
    input wire                            AP_AXIMM_0_AWVALID,
    output  wire                            AP_AXIMM_0_AWREADY,
    input wire [M_AXIMM_0_DATA_WIDTH-1:0]   AP_AXIMM_0_WDATA,
    input wire [M_AXIMM_0_DATA_WIDTH/8-1:0] AP_AXIMM_0_WSTRB,
    input wire                            AP_AXIMM_0_WLAST,
    input wire                            AP_AXIMM_0_WVALID,
    output  wire                            AP_AXIMM_0_WREADY,
    output  wire [1:0]                      AP_AXIMM_0_BRESP,
    output  wire                            AP_AXIMM_0_BVALID,
    input wire                            AP_AXIMM_0_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_0_ARADDR,
    input wire [7:0]                      AP_AXIMM_0_ARLEN,
    input wire [2:0]                      AP_AXIMM_0_ARSIZE,
    input wire [1:0]                      AP_AXIMM_0_ARBURST,
    input wire [1:0]                      AP_AXIMM_0_ARLOCK,
    input wire [3:0]                      AP_AXIMM_0_ARCACHE,
    input wire [2:0]                      AP_AXIMM_0_ARPROT,
    input wire [3:0]                      AP_AXIMM_0_ARREGION,
    input wire [3:0]                      AP_AXIMM_0_ARQOS,
    input wire                            AP_AXIMM_0_ARVALID,
    output  wire                            AP_AXIMM_0_ARREADY,
    output  wire [M_AXIMM_0_DATA_WIDTH-1:0]   AP_AXIMM_0_RDATA,
    output  wire [1:0]                      AP_AXIMM_0_RRESP,
    output  wire                            AP_AXIMM_0_RLAST,
    output  wire                            AP_AXIMM_0_RVALID,
    input  wire                            AP_AXIMM_0_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_0_AWADDR,
    output wire [7:0]                      M_AXIMM_0_AWLEN,
    output wire [2:0]                      M_AXIMM_0_AWSIZE,
    output wire [1:0]                      M_AXIMM_0_AWBURST,
    output wire [1:0]                      M_AXIMM_0_AWLOCK,
    output wire [3:0]                      M_AXIMM_0_AWCACHE,
    output wire [2:0]                      M_AXIMM_0_AWPROT,
    output wire [3:0]                      M_AXIMM_0_AWREGION,
    output wire [3:0]                      M_AXIMM_0_AWQOS,
    output wire                            M_AXIMM_0_AWVALID,
    input  wire                            M_AXIMM_0_AWREADY,
    output wire [M_AXIMM_0_DATA_WIDTH-1:0]   M_AXIMM_0_WDATA,
    output wire [M_AXIMM_0_DATA_WIDTH/8-1:0] M_AXIMM_0_WSTRB,
    output wire                            M_AXIMM_0_WLAST,
    output wire                            M_AXIMM_0_WVALID,
    input  wire                            M_AXIMM_0_WREADY,
    input  wire [1:0]                      M_AXIMM_0_BRESP,
    input  wire                            M_AXIMM_0_BVALID,
    output wire                            M_AXIMM_0_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_0_ARADDR,
    output wire [7:0]                      M_AXIMM_0_ARLEN,
    output wire [2:0]                      M_AXIMM_0_ARSIZE,
    output wire [1:0]                      M_AXIMM_0_ARBURST,
    output wire [1:0]                      M_AXIMM_0_ARLOCK,
    output wire [3:0]                      M_AXIMM_0_ARCACHE,
    output wire [2:0]                      M_AXIMM_0_ARPROT,
    output wire [3:0]                      M_AXIMM_0_ARREGION,
    output wire [3:0]                      M_AXIMM_0_ARQOS,
    output wire                            M_AXIMM_0_ARVALID,
    input  wire                            M_AXIMM_0_ARREADY,
    input  wire [M_AXIMM_0_DATA_WIDTH-1:0]   M_AXIMM_0_RDATA,
    input  wire [1:0]                      M_AXIMM_0_RRESP,
    input  wire                            M_AXIMM_0_RLAST,
    input  wire                            M_AXIMM_0_RVALID,
    output wire                            M_AXIMM_0_RREADY,
    //AXI-MM pass-through interface 1
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_1_AWADDR,
    input wire [7:0]                      AP_AXIMM_1_AWLEN,
    input wire [2:0]                      AP_AXIMM_1_AWSIZE,
    input wire [1:0]                      AP_AXIMM_1_AWBURST,
    input wire [1:0]                      AP_AXIMM_1_AWLOCK,
    input wire [3:0]                      AP_AXIMM_1_AWCACHE,
    input wire [2:0]                      AP_AXIMM_1_AWPROT,
    input wire [3:0]                      AP_AXIMM_1_AWREGION,
    input wire [3:0]                      AP_AXIMM_1_AWQOS,
    input wire                            AP_AXIMM_1_AWVALID,
    output  wire                            AP_AXIMM_1_AWREADY,
    input wire [M_AXIMM_1_DATA_WIDTH-1:0]   AP_AXIMM_1_WDATA,
    input wire [M_AXIMM_1_DATA_WIDTH/8-1:0] AP_AXIMM_1_WSTRB,
    input wire                            AP_AXIMM_1_WLAST,
    input wire                            AP_AXIMM_1_WVALID,
    output  wire                            AP_AXIMM_1_WREADY,
    output  wire [1:0]                      AP_AXIMM_1_BRESP,
    output  wire                            AP_AXIMM_1_BVALID,
    input wire                            AP_AXIMM_1_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_1_ARADDR,
    input wire [7:0]                      AP_AXIMM_1_ARLEN,
    input wire [2:0]                      AP_AXIMM_1_ARSIZE,
    input wire [1:0]                      AP_AXIMM_1_ARBURST,
    input wire [1:0]                      AP_AXIMM_1_ARLOCK,
    input wire [3:0]                      AP_AXIMM_1_ARCACHE,
    input wire [2:0]                      AP_AXIMM_1_ARPROT,
    input wire [3:0]                      AP_AXIMM_1_ARREGION,
    input wire [3:0]                      AP_AXIMM_1_ARQOS,
    input wire                            AP_AXIMM_1_ARVALID,
    output  wire                            AP_AXIMM_1_ARREADY,
    output  wire [M_AXIMM_1_DATA_WIDTH-1:0]   AP_AXIMM_1_RDATA,
    output  wire [1:0]                      AP_AXIMM_1_RRESP,
    output  wire                            AP_AXIMM_1_RLAST,
    output  wire                            AP_AXIMM_1_RVALID,
    input  wire                            AP_AXIMM_1_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_1_AWADDR,
    output wire [7:0]                      M_AXIMM_1_AWLEN,
    output wire [2:0]                      M_AXIMM_1_AWSIZE,
    output wire [1:0]                      M_AXIMM_1_AWBURST,
    output wire [1:0]                      M_AXIMM_1_AWLOCK,
    output wire [3:0]                      M_AXIMM_1_AWCACHE,
    output wire [2:0]                      M_AXIMM_1_AWPROT,
    output wire [3:0]                      M_AXIMM_1_AWREGION,
    output wire [3:0]                      M_AXIMM_1_AWQOS,
    output wire                            M_AXIMM_1_AWVALID,
    input  wire                            M_AXIMM_1_AWREADY,
    output wire [M_AXIMM_1_DATA_WIDTH-1:0]   M_AXIMM_1_WDATA,
    output wire [M_AXIMM_1_DATA_WIDTH/8-1:0] M_AXIMM_1_WSTRB,
    output wire                            M_AXIMM_1_WLAST,
    output wire                            M_AXIMM_1_WVALID,
    input  wire                            M_AXIMM_1_WREADY,
    input  wire [1:0]                      M_AXIMM_1_BRESP,
    input  wire                            M_AXIMM_1_BVALID,
    output wire                            M_AXIMM_1_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_1_ARADDR,
    output wire [7:0]                      M_AXIMM_1_ARLEN,
    output wire [2:0]                      M_AXIMM_1_ARSIZE,
    output wire [1:0]                      M_AXIMM_1_ARBURST,
    output wire [1:0]                      M_AXIMM_1_ARLOCK,
    output wire [3:0]                      M_AXIMM_1_ARCACHE,
    output wire [2:0]                      M_AXIMM_1_ARPROT,
    output wire [3:0]                      M_AXIMM_1_ARREGION,
    output wire [3:0]                      M_AXIMM_1_ARQOS,
    output wire                            M_AXIMM_1_ARVALID,
    input  wire                            M_AXIMM_1_ARREADY,
    input  wire [M_AXIMM_1_DATA_WIDTH-1:0]   M_AXIMM_1_RDATA,
    input  wire [1:0]                      M_AXIMM_1_RRESP,
    input  wire                            M_AXIMM_1_RLAST,
    input  wire                            M_AXIMM_1_RVALID,
    output wire                            M_AXIMM_1_RREADY,
    //AXI-MM pass-through interface 2
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_2_AWADDR,
    input wire [7:0]                      AP_AXIMM_2_AWLEN,
    input wire [2:0]                      AP_AXIMM_2_AWSIZE,
    input wire [1:0]                      AP_AXIMM_2_AWBURST,
    input wire [1:0]                      AP_AXIMM_2_AWLOCK,
    input wire [3:0]                      AP_AXIMM_2_AWCACHE,
    input wire [2:0]                      AP_AXIMM_2_AWPROT,
    input wire [3:0]                      AP_AXIMM_2_AWREGION,
    input wire [3:0]                      AP_AXIMM_2_AWQOS,
    input wire                            AP_AXIMM_2_AWVALID,
    output  wire                            AP_AXIMM_2_AWREADY,
    input wire [M_AXIMM_2_DATA_WIDTH-1:0]   AP_AXIMM_2_WDATA,
    input wire [M_AXIMM_2_DATA_WIDTH/8-1:0] AP_AXIMM_2_WSTRB,
    input wire                            AP_AXIMM_2_WLAST,
    input wire                            AP_AXIMM_2_WVALID,
    output  wire                            AP_AXIMM_2_WREADY,
    output  wire [1:0]                      AP_AXIMM_2_BRESP,
    output  wire                            AP_AXIMM_2_BVALID,
    input wire                            AP_AXIMM_2_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_2_ARADDR,
    input wire [7:0]                      AP_AXIMM_2_ARLEN,
    input wire [2:0]                      AP_AXIMM_2_ARSIZE,
    input wire [1:0]                      AP_AXIMM_2_ARBURST,
    input wire [1:0]                      AP_AXIMM_2_ARLOCK,
    input wire [3:0]                      AP_AXIMM_2_ARCACHE,
    input wire [2:0]                      AP_AXIMM_2_ARPROT,
    input wire [3:0]                      AP_AXIMM_2_ARREGION,
    input wire [3:0]                      AP_AXIMM_2_ARQOS,
    input wire                            AP_AXIMM_2_ARVALID,
    output  wire                            AP_AXIMM_2_ARREADY,
    output  wire [M_AXIMM_2_DATA_WIDTH-1:0]   AP_AXIMM_2_RDATA,
    output  wire [1:0]                      AP_AXIMM_2_RRESP,
    output  wire                            AP_AXIMM_2_RLAST,
    output  wire                            AP_AXIMM_2_RVALID,
    input  wire                            AP_AXIMM_2_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_2_AWADDR,
    output wire [7:0]                      M_AXIMM_2_AWLEN,
    output wire [2:0]                      M_AXIMM_2_AWSIZE,
    output wire [1:0]                      M_AXIMM_2_AWBURST,
    output wire [1:0]                      M_AXIMM_2_AWLOCK,
    output wire [3:0]                      M_AXIMM_2_AWCACHE,
    output wire [2:0]                      M_AXIMM_2_AWPROT,
    output wire [3:0]                      M_AXIMM_2_AWREGION,
    output wire [3:0]                      M_AXIMM_2_AWQOS,
    output wire                            M_AXIMM_2_AWVALID,
    input  wire                            M_AXIMM_2_AWREADY,
    output wire [M_AXIMM_2_DATA_WIDTH-1:0]   M_AXIMM_2_WDATA,
    output wire [M_AXIMM_2_DATA_WIDTH/8-1:0] M_AXIMM_2_WSTRB,
    output wire                            M_AXIMM_2_WLAST,
    output wire                            M_AXIMM_2_WVALID,
    input  wire                            M_AXIMM_2_WREADY,
    input  wire [1:0]                      M_AXIMM_2_BRESP,
    input  wire                            M_AXIMM_2_BVALID,
    output wire                            M_AXIMM_2_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_2_ARADDR,
    output wire [7:0]                      M_AXIMM_2_ARLEN,
    output wire [2:0]                      M_AXIMM_2_ARSIZE,
    output wire [1:0]                      M_AXIMM_2_ARBURST,
    output wire [1:0]                      M_AXIMM_2_ARLOCK,
    output wire [3:0]                      M_AXIMM_2_ARCACHE,
    output wire [2:0]                      M_AXIMM_2_ARPROT,
    output wire [3:0]                      M_AXIMM_2_ARREGION,
    output wire [3:0]                      M_AXIMM_2_ARQOS,
    output wire                            M_AXIMM_2_ARVALID,
    input  wire                            M_AXIMM_2_ARREADY,
    input  wire [M_AXIMM_2_DATA_WIDTH-1:0]   M_AXIMM_2_RDATA,
    input  wire [1:0]                      M_AXIMM_2_RRESP,
    input  wire                            M_AXIMM_2_RLAST,
    input  wire                            M_AXIMM_2_RVALID,
    output wire                            M_AXIMM_2_RREADY,
    //AXI-MM pass-through interface 3
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_3_AWADDR,
    input wire [7:0]                      AP_AXIMM_3_AWLEN,
    input wire [2:0]                      AP_AXIMM_3_AWSIZE,
    input wire [1:0]                      AP_AXIMM_3_AWBURST,
    input wire [1:0]                      AP_AXIMM_3_AWLOCK,
    input wire [3:0]                      AP_AXIMM_3_AWCACHE,
    input wire [2:0]                      AP_AXIMM_3_AWPROT,
    input wire [3:0]                      AP_AXIMM_3_AWREGION,
    input wire [3:0]                      AP_AXIMM_3_AWQOS,
    input wire                            AP_AXIMM_3_AWVALID,
    output  wire                            AP_AXIMM_3_AWREADY,
    input wire [M_AXIMM_3_DATA_WIDTH-1:0]   AP_AXIMM_3_WDATA,
    input wire [M_AXIMM_3_DATA_WIDTH/8-1:0] AP_AXIMM_3_WSTRB,
    input wire                            AP_AXIMM_3_WLAST,
    input wire                            AP_AXIMM_3_WVALID,
    output  wire                            AP_AXIMM_3_WREADY,
    output  wire [1:0]                      AP_AXIMM_3_BRESP,
    output  wire                            AP_AXIMM_3_BVALID,
    input wire                            AP_AXIMM_3_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_3_ARADDR,
    input wire [7:0]                      AP_AXIMM_3_ARLEN,
    input wire [2:0]                      AP_AXIMM_3_ARSIZE,
    input wire [1:0]                      AP_AXIMM_3_ARBURST,
    input wire [1:0]                      AP_AXIMM_3_ARLOCK,
    input wire [3:0]                      AP_AXIMM_3_ARCACHE,
    input wire [2:0]                      AP_AXIMM_3_ARPROT,
    input wire [3:0]                      AP_AXIMM_3_ARREGION,
    input wire [3:0]                      AP_AXIMM_3_ARQOS,
    input wire                            AP_AXIMM_3_ARVALID,
    output  wire                            AP_AXIMM_3_ARREADY,
    output  wire [M_AXIMM_3_DATA_WIDTH-1:0]   AP_AXIMM_3_RDATA,
    output  wire [1:0]                      AP_AXIMM_3_RRESP,
    output  wire                            AP_AXIMM_3_RLAST,
    output  wire                            AP_AXIMM_3_RVALID,
    input  wire                            AP_AXIMM_3_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_3_AWADDR,
    output wire [7:0]                      M_AXIMM_3_AWLEN,
    output wire [2:0]                      M_AXIMM_3_AWSIZE,
    output wire [1:0]                      M_AXIMM_3_AWBURST,
    output wire [1:0]                      M_AXIMM_3_AWLOCK,
    output wire [3:0]                      M_AXIMM_3_AWCACHE,
    output wire [2:0]                      M_AXIMM_3_AWPROT,
    output wire [3:0]                      M_AXIMM_3_AWREGION,
    output wire [3:0]                      M_AXIMM_3_AWQOS,
    output wire                            M_AXIMM_3_AWVALID,
    input  wire                            M_AXIMM_3_AWREADY,
    output wire [M_AXIMM_3_DATA_WIDTH-1:0]   M_AXIMM_3_WDATA,
    output wire [M_AXIMM_3_DATA_WIDTH/8-1:0] M_AXIMM_3_WSTRB,
    output wire                            M_AXIMM_3_WLAST,
    output wire                            M_AXIMM_3_WVALID,
    input  wire                            M_AXIMM_3_WREADY,
    input  wire [1:0]                      M_AXIMM_3_BRESP,
    input  wire                            M_AXIMM_3_BVALID,
    output wire                            M_AXIMM_3_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_3_ARADDR,
    output wire [7:0]                      M_AXIMM_3_ARLEN,
    output wire [2:0]                      M_AXIMM_3_ARSIZE,
    output wire [1:0]                      M_AXIMM_3_ARBURST,
    output wire [1:0]                      M_AXIMM_3_ARLOCK,
    output wire [3:0]                      M_AXIMM_3_ARCACHE,
    output wire [2:0]                      M_AXIMM_3_ARPROT,
    output wire [3:0]                      M_AXIMM_3_ARREGION,
    output wire [3:0]                      M_AXIMM_3_ARQOS,
    output wire                            M_AXIMM_3_ARVALID,
    input  wire                            M_AXIMM_3_ARREADY,
    input  wire [M_AXIMM_3_DATA_WIDTH-1:0]   M_AXIMM_3_RDATA,
    input  wire [1:0]                      M_AXIMM_3_RRESP,
    input  wire                            M_AXIMM_3_RLAST,
    input  wire                            M_AXIMM_3_RVALID,
    output wire                            M_AXIMM_3_RREADY,
    //AXI-MM pass-through interface 4
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_4_AWADDR,
    input wire [7:0]                      AP_AXIMM_4_AWLEN,
    input wire [2:0]                      AP_AXIMM_4_AWSIZE,
    input wire [1:0]                      AP_AXIMM_4_AWBURST,
    input wire [1:0]                      AP_AXIMM_4_AWLOCK,
    input wire [3:0]                      AP_AXIMM_4_AWCACHE,
    input wire [2:0]                      AP_AXIMM_4_AWPROT,
    input wire [3:0]                      AP_AXIMM_4_AWREGION,
    input wire [3:0]                      AP_AXIMM_4_AWQOS,
    input wire                            AP_AXIMM_4_AWVALID,
    output  wire                            AP_AXIMM_4_AWREADY,
    input wire [M_AXIMM_4_DATA_WIDTH-1:0]   AP_AXIMM_4_WDATA,
    input wire [M_AXIMM_4_DATA_WIDTH/8-1:0] AP_AXIMM_4_WSTRB,
    input wire                            AP_AXIMM_4_WLAST,
    input wire                            AP_AXIMM_4_WVALID,
    output  wire                            AP_AXIMM_4_WREADY,
    output  wire [1:0]                      AP_AXIMM_4_BRESP,
    output  wire                            AP_AXIMM_4_BVALID,
    input wire                            AP_AXIMM_4_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_4_ARADDR,
    input wire [7:0]                      AP_AXIMM_4_ARLEN,
    input wire [2:0]                      AP_AXIMM_4_ARSIZE,
    input wire [1:0]                      AP_AXIMM_4_ARBURST,
    input wire [1:0]                      AP_AXIMM_4_ARLOCK,
    input wire [3:0]                      AP_AXIMM_4_ARCACHE,
    input wire [2:0]                      AP_AXIMM_4_ARPROT,
    input wire [3:0]                      AP_AXIMM_4_ARREGION,
    input wire [3:0]                      AP_AXIMM_4_ARQOS,
    input wire                            AP_AXIMM_4_ARVALID,
    output  wire                            AP_AXIMM_4_ARREADY,
    output  wire [M_AXIMM_4_DATA_WIDTH-1:0]   AP_AXIMM_4_RDATA,
    output  wire [1:0]                      AP_AXIMM_4_RRESP,
    output  wire                            AP_AXIMM_4_RLAST,
    output  wire                            AP_AXIMM_4_RVALID,
    input  wire                            AP_AXIMM_4_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_4_AWADDR,
    output wire [7:0]                      M_AXIMM_4_AWLEN,
    output wire [2:0]                      M_AXIMM_4_AWSIZE,
    output wire [1:0]                      M_AXIMM_4_AWBURST,
    output wire [1:0]                      M_AXIMM_4_AWLOCK,
    output wire [3:0]                      M_AXIMM_4_AWCACHE,
    output wire [2:0]                      M_AXIMM_4_AWPROT,
    output wire [3:0]                      M_AXIMM_4_AWREGION,
    output wire [3:0]                      M_AXIMM_4_AWQOS,
    output wire                            M_AXIMM_4_AWVALID,
    input  wire                            M_AXIMM_4_AWREADY,
    output wire [M_AXIMM_4_DATA_WIDTH-1:0]   M_AXIMM_4_WDATA,
    output wire [M_AXIMM_4_DATA_WIDTH/8-1:0] M_AXIMM_4_WSTRB,
    output wire                            M_AXIMM_4_WLAST,
    output wire                            M_AXIMM_4_WVALID,
    input  wire                            M_AXIMM_4_WREADY,
    input  wire [1:0]                      M_AXIMM_4_BRESP,
    input  wire                            M_AXIMM_4_BVALID,
    output wire                            M_AXIMM_4_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_4_ARADDR,
    output wire [7:0]                      M_AXIMM_4_ARLEN,
    output wire [2:0]                      M_AXIMM_4_ARSIZE,
    output wire [1:0]                      M_AXIMM_4_ARBURST,
    output wire [1:0]                      M_AXIMM_4_ARLOCK,
    output wire [3:0]                      M_AXIMM_4_ARCACHE,
    output wire [2:0]                      M_AXIMM_4_ARPROT,
    output wire [3:0]                      M_AXIMM_4_ARREGION,
    output wire [3:0]                      M_AXIMM_4_ARQOS,
    output wire                            M_AXIMM_4_ARVALID,
    input  wire                            M_AXIMM_4_ARREADY,
    input  wire [M_AXIMM_4_DATA_WIDTH-1:0]   M_AXIMM_4_RDATA,
    input  wire [1:0]                      M_AXIMM_4_RRESP,
    input  wire                            M_AXIMM_4_RLAST,
    input  wire                            M_AXIMM_4_RVALID,
    output wire                            M_AXIMM_4_RREADY,
    //AXI-MM pass-through interface 5
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_5_AWADDR,
    input wire [7:0]                      AP_AXIMM_5_AWLEN,
    input wire [2:0]                      AP_AXIMM_5_AWSIZE,
    input wire [1:0]                      AP_AXIMM_5_AWBURST,
    input wire [1:0]                      AP_AXIMM_5_AWLOCK,
    input wire [3:0]                      AP_AXIMM_5_AWCACHE,
    input wire [2:0]                      AP_AXIMM_5_AWPROT,
    input wire [3:0]                      AP_AXIMM_5_AWREGION,
    input wire [3:0]                      AP_AXIMM_5_AWQOS,
    input wire                            AP_AXIMM_5_AWVALID,
    output  wire                            AP_AXIMM_5_AWREADY,
    input wire [M_AXIMM_5_DATA_WIDTH-1:0]   AP_AXIMM_5_WDATA,
    input wire [M_AXIMM_5_DATA_WIDTH/8-1:0] AP_AXIMM_5_WSTRB,
    input wire                            AP_AXIMM_5_WLAST,
    input wire                            AP_AXIMM_5_WVALID,
    output  wire                            AP_AXIMM_5_WREADY,
    output  wire [1:0]                      AP_AXIMM_5_BRESP,
    output  wire                            AP_AXIMM_5_BVALID,
    input wire                            AP_AXIMM_5_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_5_ARADDR,
    input wire [7:0]                      AP_AXIMM_5_ARLEN,
    input wire [2:0]                      AP_AXIMM_5_ARSIZE,
    input wire [1:0]                      AP_AXIMM_5_ARBURST,
    input wire [1:0]                      AP_AXIMM_5_ARLOCK,
    input wire [3:0]                      AP_AXIMM_5_ARCACHE,
    input wire [2:0]                      AP_AXIMM_5_ARPROT,
    input wire [3:0]                      AP_AXIMM_5_ARREGION,
    input wire [3:0]                      AP_AXIMM_5_ARQOS,
    input wire                            AP_AXIMM_5_ARVALID,
    output  wire                            AP_AXIMM_5_ARREADY,
    output  wire [M_AXIMM_5_DATA_WIDTH-1:0]   AP_AXIMM_5_RDATA,
    output  wire [1:0]                      AP_AXIMM_5_RRESP,
    output  wire                            AP_AXIMM_5_RLAST,
    output  wire                            AP_AXIMM_5_RVALID,
    input  wire                            AP_AXIMM_5_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_5_AWADDR,
    output wire [7:0]                      M_AXIMM_5_AWLEN,
    output wire [2:0]                      M_AXIMM_5_AWSIZE,
    output wire [1:0]                      M_AXIMM_5_AWBURST,
    output wire [1:0]                      M_AXIMM_5_AWLOCK,
    output wire [3:0]                      M_AXIMM_5_AWCACHE,
    output wire [2:0]                      M_AXIMM_5_AWPROT,
    output wire [3:0]                      M_AXIMM_5_AWREGION,
    output wire [3:0]                      M_AXIMM_5_AWQOS,
    output wire                            M_AXIMM_5_AWVALID,
    input  wire                            M_AXIMM_5_AWREADY,
    output wire [M_AXIMM_5_DATA_WIDTH-1:0]   M_AXIMM_5_WDATA,
    output wire [M_AXIMM_5_DATA_WIDTH/8-1:0] M_AXIMM_5_WSTRB,
    output wire                            M_AXIMM_5_WLAST,
    output wire                            M_AXIMM_5_WVALID,
    input  wire                            M_AXIMM_5_WREADY,
    input  wire [1:0]                      M_AXIMM_5_BRESP,
    input  wire                            M_AXIMM_5_BVALID,
    output wire                            M_AXIMM_5_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_5_ARADDR,
    output wire [7:0]                      M_AXIMM_5_ARLEN,
    output wire [2:0]                      M_AXIMM_5_ARSIZE,
    output wire [1:0]                      M_AXIMM_5_ARBURST,
    output wire [1:0]                      M_AXIMM_5_ARLOCK,
    output wire [3:0]                      M_AXIMM_5_ARCACHE,
    output wire [2:0]                      M_AXIMM_5_ARPROT,
    output wire [3:0]                      M_AXIMM_5_ARREGION,
    output wire [3:0]                      M_AXIMM_5_ARQOS,
    output wire                            M_AXIMM_5_ARVALID,
    input  wire                            M_AXIMM_5_ARREADY,
    input  wire [M_AXIMM_5_DATA_WIDTH-1:0]   M_AXIMM_5_RDATA,
    input  wire [1:0]                      M_AXIMM_5_RRESP,
    input  wire                            M_AXIMM_5_RLAST,
    input  wire                            M_AXIMM_5_RVALID,
    output wire                            M_AXIMM_5_RREADY,
    //AXI-MM pass-through interface 6
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_6_AWADDR,
    input wire [7:0]                      AP_AXIMM_6_AWLEN,
    input wire [2:0]                      AP_AXIMM_6_AWSIZE,
    input wire [1:0]                      AP_AXIMM_6_AWBURST,
    input wire [1:0]                      AP_AXIMM_6_AWLOCK,
    input wire [3:0]                      AP_AXIMM_6_AWCACHE,
    input wire [2:0]                      AP_AXIMM_6_AWPROT,
    input wire [3:0]                      AP_AXIMM_6_AWREGION,
    input wire [3:0]                      AP_AXIMM_6_AWQOS,
    input wire                            AP_AXIMM_6_AWVALID,
    output  wire                            AP_AXIMM_6_AWREADY,
    input wire [M_AXIMM_6_DATA_WIDTH-1:0]   AP_AXIMM_6_WDATA,
    input wire [M_AXIMM_6_DATA_WIDTH/8-1:0] AP_AXIMM_6_WSTRB,
    input wire                            AP_AXIMM_6_WLAST,
    input wire                            AP_AXIMM_6_WVALID,
    output  wire                            AP_AXIMM_6_WREADY,
    output  wire [1:0]                      AP_AXIMM_6_BRESP,
    output  wire                            AP_AXIMM_6_BVALID,
    input wire                            AP_AXIMM_6_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_6_ARADDR,
    input wire [7:0]                      AP_AXIMM_6_ARLEN,
    input wire [2:0]                      AP_AXIMM_6_ARSIZE,
    input wire [1:0]                      AP_AXIMM_6_ARBURST,
    input wire [1:0]                      AP_AXIMM_6_ARLOCK,
    input wire [3:0]                      AP_AXIMM_6_ARCACHE,
    input wire [2:0]                      AP_AXIMM_6_ARPROT,
    input wire [3:0]                      AP_AXIMM_6_ARREGION,
    input wire [3:0]                      AP_AXIMM_6_ARQOS,
    input wire                            AP_AXIMM_6_ARVALID,
    output  wire                            AP_AXIMM_6_ARREADY,
    output  wire [M_AXIMM_6_DATA_WIDTH-1:0]   AP_AXIMM_6_RDATA,
    output  wire [1:0]                      AP_AXIMM_6_RRESP,
    output  wire                            AP_AXIMM_6_RLAST,
    output  wire                            AP_AXIMM_6_RVALID,
    input  wire                            AP_AXIMM_6_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_6_AWADDR,
    output wire [7:0]                      M_AXIMM_6_AWLEN,
    output wire [2:0]                      M_AXIMM_6_AWSIZE,
    output wire [1:0]                      M_AXIMM_6_AWBURST,
    output wire [1:0]                      M_AXIMM_6_AWLOCK,
    output wire [3:0]                      M_AXIMM_6_AWCACHE,
    output wire [2:0]                      M_AXIMM_6_AWPROT,
    output wire [3:0]                      M_AXIMM_6_AWREGION,
    output wire [3:0]                      M_AXIMM_6_AWQOS,
    output wire                            M_AXIMM_6_AWVALID,
    input  wire                            M_AXIMM_6_AWREADY,
    output wire [M_AXIMM_6_DATA_WIDTH-1:0]   M_AXIMM_6_WDATA,
    output wire [M_AXIMM_6_DATA_WIDTH/8-1:0] M_AXIMM_6_WSTRB,
    output wire                            M_AXIMM_6_WLAST,
    output wire                            M_AXIMM_6_WVALID,
    input  wire                            M_AXIMM_6_WREADY,
    input  wire [1:0]                      M_AXIMM_6_BRESP,
    input  wire                            M_AXIMM_6_BVALID,
    output wire                            M_AXIMM_6_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_6_ARADDR,
    output wire [7:0]                      M_AXIMM_6_ARLEN,
    output wire [2:0]                      M_AXIMM_6_ARSIZE,
    output wire [1:0]                      M_AXIMM_6_ARBURST,
    output wire [1:0]                      M_AXIMM_6_ARLOCK,
    output wire [3:0]                      M_AXIMM_6_ARCACHE,
    output wire [2:0]                      M_AXIMM_6_ARPROT,
    output wire [3:0]                      M_AXIMM_6_ARREGION,
    output wire [3:0]                      M_AXIMM_6_ARQOS,
    output wire                            M_AXIMM_6_ARVALID,
    input  wire                            M_AXIMM_6_ARREADY,
    input  wire [M_AXIMM_6_DATA_WIDTH-1:0]   M_AXIMM_6_RDATA,
    input  wire [1:0]                      M_AXIMM_6_RRESP,
    input  wire                            M_AXIMM_6_RLAST,
    input  wire                            M_AXIMM_6_RVALID,
    output wire                            M_AXIMM_6_RREADY,
    //AXI-MM pass-through interface 7
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_7_AWADDR,
    input wire [7:0]                      AP_AXIMM_7_AWLEN,
    input wire [2:0]                      AP_AXIMM_7_AWSIZE,
    input wire [1:0]                      AP_AXIMM_7_AWBURST,
    input wire [1:0]                      AP_AXIMM_7_AWLOCK,
    input wire [3:0]                      AP_AXIMM_7_AWCACHE,
    input wire [2:0]                      AP_AXIMM_7_AWPROT,
    input wire [3:0]                      AP_AXIMM_7_AWREGION,
    input wire [3:0]                      AP_AXIMM_7_AWQOS,
    input wire                            AP_AXIMM_7_AWVALID,
    output  wire                            AP_AXIMM_7_AWREADY,
    input wire [M_AXIMM_7_DATA_WIDTH-1:0]   AP_AXIMM_7_WDATA,
    input wire [M_AXIMM_7_DATA_WIDTH/8-1:0] AP_AXIMM_7_WSTRB,
    input wire                            AP_AXIMM_7_WLAST,
    input wire                            AP_AXIMM_7_WVALID,
    output  wire                            AP_AXIMM_7_WREADY,
    output  wire [1:0]                      AP_AXIMM_7_BRESP,
    output  wire                            AP_AXIMM_7_BVALID,
    input wire                            AP_AXIMM_7_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_7_ARADDR,
    input wire [7:0]                      AP_AXIMM_7_ARLEN,
    input wire [2:0]                      AP_AXIMM_7_ARSIZE,
    input wire [1:0]                      AP_AXIMM_7_ARBURST,
    input wire [1:0]                      AP_AXIMM_7_ARLOCK,
    input wire [3:0]                      AP_AXIMM_7_ARCACHE,
    input wire [2:0]                      AP_AXIMM_7_ARPROT,
    input wire [3:0]                      AP_AXIMM_7_ARREGION,
    input wire [3:0]                      AP_AXIMM_7_ARQOS,
    input wire                            AP_AXIMM_7_ARVALID,
    output  wire                            AP_AXIMM_7_ARREADY,
    output  wire [M_AXIMM_7_DATA_WIDTH-1:0]   AP_AXIMM_7_RDATA,
    output  wire [1:0]                      AP_AXIMM_7_RRESP,
    output  wire                            AP_AXIMM_7_RLAST,
    output  wire                            AP_AXIMM_7_RVALID,
    input  wire                            AP_AXIMM_7_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_7_AWADDR,
    output wire [7:0]                      M_AXIMM_7_AWLEN,
    output wire [2:0]                      M_AXIMM_7_AWSIZE,
    output wire [1:0]                      M_AXIMM_7_AWBURST,
    output wire [1:0]                      M_AXIMM_7_AWLOCK,
    output wire [3:0]                      M_AXIMM_7_AWCACHE,
    output wire [2:0]                      M_AXIMM_7_AWPROT,
    output wire [3:0]                      M_AXIMM_7_AWREGION,
    output wire [3:0]                      M_AXIMM_7_AWQOS,
    output wire                            M_AXIMM_7_AWVALID,
    input  wire                            M_AXIMM_7_AWREADY,
    output wire [M_AXIMM_7_DATA_WIDTH-1:0]   M_AXIMM_7_WDATA,
    output wire [M_AXIMM_7_DATA_WIDTH/8-1:0] M_AXIMM_7_WSTRB,
    output wire                            M_AXIMM_7_WLAST,
    output wire                            M_AXIMM_7_WVALID,
    input  wire                            M_AXIMM_7_WREADY,
    input  wire [1:0]                      M_AXIMM_7_BRESP,
    input  wire                            M_AXIMM_7_BVALID,
    output wire                            M_AXIMM_7_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_7_ARADDR,
    output wire [7:0]                      M_AXIMM_7_ARLEN,
    output wire [2:0]                      M_AXIMM_7_ARSIZE,
    output wire [1:0]                      M_AXIMM_7_ARBURST,
    output wire [1:0]                      M_AXIMM_7_ARLOCK,
    output wire [3:0]                      M_AXIMM_7_ARCACHE,
    output wire [2:0]                      M_AXIMM_7_ARPROT,
    output wire [3:0]                      M_AXIMM_7_ARREGION,
    output wire [3:0]                      M_AXIMM_7_ARQOS,
    output wire                            M_AXIMM_7_ARVALID,
    input  wire                            M_AXIMM_7_ARREADY,
    input  wire [M_AXIMM_7_DATA_WIDTH-1:0]   M_AXIMM_7_RDATA,
    input  wire [1:0]                      M_AXIMM_7_RRESP,
    input  wire                            M_AXIMM_7_RLAST,
    input  wire                            M_AXIMM_7_RVALID,
    output wire                            M_AXIMM_7_RREADY,
    //AXI-MM pass-through interface 8
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_8_AWADDR,
    input wire [7:0]                      AP_AXIMM_8_AWLEN,
    input wire [2:0]                      AP_AXIMM_8_AWSIZE,
    input wire [1:0]                      AP_AXIMM_8_AWBURST,
    input wire [1:0]                      AP_AXIMM_8_AWLOCK,
    input wire [3:0]                      AP_AXIMM_8_AWCACHE,
    input wire [2:0]                      AP_AXIMM_8_AWPROT,
    input wire [3:0]                      AP_AXIMM_8_AWREGION,
    input wire [3:0]                      AP_AXIMM_8_AWQOS,
    input wire                            AP_AXIMM_8_AWVALID,
    output  wire                            AP_AXIMM_8_AWREADY,
    input wire [M_AXIMM_8_DATA_WIDTH-1:0]   AP_AXIMM_8_WDATA,
    input wire [M_AXIMM_8_DATA_WIDTH/8-1:0] AP_AXIMM_8_WSTRB,
    input wire                            AP_AXIMM_8_WLAST,
    input wire                            AP_AXIMM_8_WVALID,
    output  wire                            AP_AXIMM_8_WREADY,
    output  wire [1:0]                      AP_AXIMM_8_BRESP,
    output  wire                            AP_AXIMM_8_BVALID,
    input wire                            AP_AXIMM_8_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_8_ARADDR,
    input wire [7:0]                      AP_AXIMM_8_ARLEN,
    input wire [2:0]                      AP_AXIMM_8_ARSIZE,
    input wire [1:0]                      AP_AXIMM_8_ARBURST,
    input wire [1:0]                      AP_AXIMM_8_ARLOCK,
    input wire [3:0]                      AP_AXIMM_8_ARCACHE,
    input wire [2:0]                      AP_AXIMM_8_ARPROT,
    input wire [3:0]                      AP_AXIMM_8_ARREGION,
    input wire [3:0]                      AP_AXIMM_8_ARQOS,
    input wire                            AP_AXIMM_8_ARVALID,
    output  wire                            AP_AXIMM_8_ARREADY,
    output  wire [M_AXIMM_8_DATA_WIDTH-1:0]   AP_AXIMM_8_RDATA,
    output  wire [1:0]                      AP_AXIMM_8_RRESP,
    output  wire                            AP_AXIMM_8_RLAST,
    output  wire                            AP_AXIMM_8_RVALID,
    input  wire                            AP_AXIMM_8_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_8_AWADDR,
    output wire [7:0]                      M_AXIMM_8_AWLEN,
    output wire [2:0]                      M_AXIMM_8_AWSIZE,
    output wire [1:0]                      M_AXIMM_8_AWBURST,
    output wire [1:0]                      M_AXIMM_8_AWLOCK,
    output wire [3:0]                      M_AXIMM_8_AWCACHE,
    output wire [2:0]                      M_AXIMM_8_AWPROT,
    output wire [3:0]                      M_AXIMM_8_AWREGION,
    output wire [3:0]                      M_AXIMM_8_AWQOS,
    output wire                            M_AXIMM_8_AWVALID,
    input  wire                            M_AXIMM_8_AWREADY,
    output wire [M_AXIMM_8_DATA_WIDTH-1:0]   M_AXIMM_8_WDATA,
    output wire [M_AXIMM_8_DATA_WIDTH/8-1:0] M_AXIMM_8_WSTRB,
    output wire                            M_AXIMM_8_WLAST,
    output wire                            M_AXIMM_8_WVALID,
    input  wire                            M_AXIMM_8_WREADY,
    input  wire [1:0]                      M_AXIMM_8_BRESP,
    input  wire                            M_AXIMM_8_BVALID,
    output wire                            M_AXIMM_8_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_8_ARADDR,
    output wire [7:0]                      M_AXIMM_8_ARLEN,
    output wire [2:0]                      M_AXIMM_8_ARSIZE,
    output wire [1:0]                      M_AXIMM_8_ARBURST,
    output wire [1:0]                      M_AXIMM_8_ARLOCK,
    output wire [3:0]                      M_AXIMM_8_ARCACHE,
    output wire [2:0]                      M_AXIMM_8_ARPROT,
    output wire [3:0]                      M_AXIMM_8_ARREGION,
    output wire [3:0]                      M_AXIMM_8_ARQOS,
    output wire                            M_AXIMM_8_ARVALID,
    input  wire                            M_AXIMM_8_ARREADY,
    input  wire [M_AXIMM_8_DATA_WIDTH-1:0]   M_AXIMM_8_RDATA,
    input  wire [1:0]                      M_AXIMM_8_RRESP,
    input  wire                            M_AXIMM_8_RLAST,
    input  wire                            M_AXIMM_8_RVALID,
    output wire                            M_AXIMM_8_RREADY,
    //AXI-MM pass-through interface 9
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_9_AWADDR,
    input wire [7:0]                      AP_AXIMM_9_AWLEN,
    input wire [2:0]                      AP_AXIMM_9_AWSIZE,
    input wire [1:0]                      AP_AXIMM_9_AWBURST,
    input wire [1:0]                      AP_AXIMM_9_AWLOCK,
    input wire [3:0]                      AP_AXIMM_9_AWCACHE,
    input wire [2:0]                      AP_AXIMM_9_AWPROT,
    input wire [3:0]                      AP_AXIMM_9_AWREGION,
    input wire [3:0]                      AP_AXIMM_9_AWQOS,
    input wire                            AP_AXIMM_9_AWVALID,
    output  wire                            AP_AXIMM_9_AWREADY,
    input wire [M_AXIMM_9_DATA_WIDTH-1:0]   AP_AXIMM_9_WDATA,
    input wire [M_AXIMM_9_DATA_WIDTH/8-1:0] AP_AXIMM_9_WSTRB,
    input wire                            AP_AXIMM_9_WLAST,
    input wire                            AP_AXIMM_9_WVALID,
    output  wire                            AP_AXIMM_9_WREADY,
    output  wire [1:0]                      AP_AXIMM_9_BRESP,
    output  wire                            AP_AXIMM_9_BVALID,
    input wire                            AP_AXIMM_9_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_9_ARADDR,
    input wire [7:0]                      AP_AXIMM_9_ARLEN,
    input wire [2:0]                      AP_AXIMM_9_ARSIZE,
    input wire [1:0]                      AP_AXIMM_9_ARBURST,
    input wire [1:0]                      AP_AXIMM_9_ARLOCK,
    input wire [3:0]                      AP_AXIMM_9_ARCACHE,
    input wire [2:0]                      AP_AXIMM_9_ARPROT,
    input wire [3:0]                      AP_AXIMM_9_ARREGION,
    input wire [3:0]                      AP_AXIMM_9_ARQOS,
    input wire                            AP_AXIMM_9_ARVALID,
    output  wire                            AP_AXIMM_9_ARREADY,
    output  wire [M_AXIMM_9_DATA_WIDTH-1:0]   AP_AXIMM_9_RDATA,
    output  wire [1:0]                      AP_AXIMM_9_RRESP,
    output  wire                            AP_AXIMM_9_RLAST,
    output  wire                            AP_AXIMM_9_RVALID,
    input  wire                            AP_AXIMM_9_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_9_AWADDR,
    output wire [7:0]                      M_AXIMM_9_AWLEN,
    output wire [2:0]                      M_AXIMM_9_AWSIZE,
    output wire [1:0]                      M_AXIMM_9_AWBURST,
    output wire [1:0]                      M_AXIMM_9_AWLOCK,
    output wire [3:0]                      M_AXIMM_9_AWCACHE,
    output wire [2:0]                      M_AXIMM_9_AWPROT,
    output wire [3:0]                      M_AXIMM_9_AWREGION,
    output wire [3:0]                      M_AXIMM_9_AWQOS,
    output wire                            M_AXIMM_9_AWVALID,
    input  wire                            M_AXIMM_9_AWREADY,
    output wire [M_AXIMM_9_DATA_WIDTH-1:0]   M_AXIMM_9_WDATA,
    output wire [M_AXIMM_9_DATA_WIDTH/8-1:0] M_AXIMM_9_WSTRB,
    output wire                            M_AXIMM_9_WLAST,
    output wire                            M_AXIMM_9_WVALID,
    input  wire                            M_AXIMM_9_WREADY,
    input  wire [1:0]                      M_AXIMM_9_BRESP,
    input  wire                            M_AXIMM_9_BVALID,
    output wire                            M_AXIMM_9_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_9_ARADDR,
    output wire [7:0]                      M_AXIMM_9_ARLEN,
    output wire [2:0]                      M_AXIMM_9_ARSIZE,
    output wire [1:0]                      M_AXIMM_9_ARBURST,
    output wire [1:0]                      M_AXIMM_9_ARLOCK,
    output wire [3:0]                      M_AXIMM_9_ARCACHE,
    output wire [2:0]                      M_AXIMM_9_ARPROT,
    output wire [3:0]                      M_AXIMM_9_ARREGION,
    output wire [3:0]                      M_AXIMM_9_ARQOS,
    output wire                            M_AXIMM_9_ARVALID,
    input  wire                            M_AXIMM_9_ARREADY,
    input  wire [M_AXIMM_9_DATA_WIDTH-1:0]   M_AXIMM_9_RDATA,
    input  wire [1:0]                      M_AXIMM_9_RRESP,
    input  wire                            M_AXIMM_9_RLAST,
    input  wire                            M_AXIMM_9_RVALID,
    output wire                            M_AXIMM_9_RREADY,
    //AXI-MM pass-through interface 10
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_10_AWADDR,
    input wire [7:0]                      AP_AXIMM_10_AWLEN,
    input wire [2:0]                      AP_AXIMM_10_AWSIZE,
    input wire [1:0]                      AP_AXIMM_10_AWBURST,
    input wire [1:0]                      AP_AXIMM_10_AWLOCK,
    input wire [3:0]                      AP_AXIMM_10_AWCACHE,
    input wire [2:0]                      AP_AXIMM_10_AWPROT,
    input wire [3:0]                      AP_AXIMM_10_AWREGION,
    input wire [3:0]                      AP_AXIMM_10_AWQOS,
    input wire                            AP_AXIMM_10_AWVALID,
    output  wire                            AP_AXIMM_10_AWREADY,
    input wire [M_AXIMM_10_DATA_WIDTH-1:0]   AP_AXIMM_10_WDATA,
    input wire [M_AXIMM_10_DATA_WIDTH/8-1:0] AP_AXIMM_10_WSTRB,
    input wire                            AP_AXIMM_10_WLAST,
    input wire                            AP_AXIMM_10_WVALID,
    output  wire                            AP_AXIMM_10_WREADY,
    output  wire [1:0]                      AP_AXIMM_10_BRESP,
    output  wire                            AP_AXIMM_10_BVALID,
    input wire                            AP_AXIMM_10_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_10_ARADDR,
    input wire [7:0]                      AP_AXIMM_10_ARLEN,
    input wire [2:0]                      AP_AXIMM_10_ARSIZE,
    input wire [1:0]                      AP_AXIMM_10_ARBURST,
    input wire [1:0]                      AP_AXIMM_10_ARLOCK,
    input wire [3:0]                      AP_AXIMM_10_ARCACHE,
    input wire [2:0]                      AP_AXIMM_10_ARPROT,
    input wire [3:0]                      AP_AXIMM_10_ARREGION,
    input wire [3:0]                      AP_AXIMM_10_ARQOS,
    input wire                            AP_AXIMM_10_ARVALID,
    output  wire                            AP_AXIMM_10_ARREADY,
    output  wire [M_AXIMM_10_DATA_WIDTH-1:0]   AP_AXIMM_10_RDATA,
    output  wire [1:0]                      AP_AXIMM_10_RRESP,
    output  wire                            AP_AXIMM_10_RLAST,
    output  wire                            AP_AXIMM_10_RVALID,
    input  wire                            AP_AXIMM_10_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_10_AWADDR,
    output wire [7:0]                      M_AXIMM_10_AWLEN,
    output wire [2:0]                      M_AXIMM_10_AWSIZE,
    output wire [1:0]                      M_AXIMM_10_AWBURST,
    output wire [1:0]                      M_AXIMM_10_AWLOCK,
    output wire [3:0]                      M_AXIMM_10_AWCACHE,
    output wire [2:0]                      M_AXIMM_10_AWPROT,
    output wire [3:0]                      M_AXIMM_10_AWREGION,
    output wire [3:0]                      M_AXIMM_10_AWQOS,
    output wire                            M_AXIMM_10_AWVALID,
    input  wire                            M_AXIMM_10_AWREADY,
    output wire [M_AXIMM_10_DATA_WIDTH-1:0]   M_AXIMM_10_WDATA,
    output wire [M_AXIMM_10_DATA_WIDTH/8-1:0] M_AXIMM_10_WSTRB,
    output wire                            M_AXIMM_10_WLAST,
    output wire                            M_AXIMM_10_WVALID,
    input  wire                            M_AXIMM_10_WREADY,
    input  wire [1:0]                      M_AXIMM_10_BRESP,
    input  wire                            M_AXIMM_10_BVALID,
    output wire                            M_AXIMM_10_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_10_ARADDR,
    output wire [7:0]                      M_AXIMM_10_ARLEN,
    output wire [2:0]                      M_AXIMM_10_ARSIZE,
    output wire [1:0]                      M_AXIMM_10_ARBURST,
    output wire [1:0]                      M_AXIMM_10_ARLOCK,
    output wire [3:0]                      M_AXIMM_10_ARCACHE,
    output wire [2:0]                      M_AXIMM_10_ARPROT,
    output wire [3:0]                      M_AXIMM_10_ARREGION,
    output wire [3:0]                      M_AXIMM_10_ARQOS,
    output wire                            M_AXIMM_10_ARVALID,
    input  wire                            M_AXIMM_10_ARREADY,
    input  wire [M_AXIMM_10_DATA_WIDTH-1:0]   M_AXIMM_10_RDATA,
    input  wire [1:0]                      M_AXIMM_10_RRESP,
    input  wire                            M_AXIMM_10_RLAST,
    input  wire                            M_AXIMM_10_RVALID,
    output wire                            M_AXIMM_10_RREADY,
    //AXI-MM pass-through interface 11
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_11_AWADDR,
    input wire [7:0]                      AP_AXIMM_11_AWLEN,
    input wire [2:0]                      AP_AXIMM_11_AWSIZE,
    input wire [1:0]                      AP_AXIMM_11_AWBURST,
    input wire [1:0]                      AP_AXIMM_11_AWLOCK,
    input wire [3:0]                      AP_AXIMM_11_AWCACHE,
    input wire [2:0]                      AP_AXIMM_11_AWPROT,
    input wire [3:0]                      AP_AXIMM_11_AWREGION,
    input wire [3:0]                      AP_AXIMM_11_AWQOS,
    input wire                            AP_AXIMM_11_AWVALID,
    output  wire                            AP_AXIMM_11_AWREADY,
    input wire [M_AXIMM_11_DATA_WIDTH-1:0]   AP_AXIMM_11_WDATA,
    input wire [M_AXIMM_11_DATA_WIDTH/8-1:0] AP_AXIMM_11_WSTRB,
    input wire                            AP_AXIMM_11_WLAST,
    input wire                            AP_AXIMM_11_WVALID,
    output  wire                            AP_AXIMM_11_WREADY,
    output  wire [1:0]                      AP_AXIMM_11_BRESP,
    output  wire                            AP_AXIMM_11_BVALID,
    input wire                            AP_AXIMM_11_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_11_ARADDR,
    input wire [7:0]                      AP_AXIMM_11_ARLEN,
    input wire [2:0]                      AP_AXIMM_11_ARSIZE,
    input wire [1:0]                      AP_AXIMM_11_ARBURST,
    input wire [1:0]                      AP_AXIMM_11_ARLOCK,
    input wire [3:0]                      AP_AXIMM_11_ARCACHE,
    input wire [2:0]                      AP_AXIMM_11_ARPROT,
    input wire [3:0]                      AP_AXIMM_11_ARREGION,
    input wire [3:0]                      AP_AXIMM_11_ARQOS,
    input wire                            AP_AXIMM_11_ARVALID,
    output  wire                            AP_AXIMM_11_ARREADY,
    output  wire [M_AXIMM_11_DATA_WIDTH-1:0]   AP_AXIMM_11_RDATA,
    output  wire [1:0]                      AP_AXIMM_11_RRESP,
    output  wire                            AP_AXIMM_11_RLAST,
    output  wire                            AP_AXIMM_11_RVALID,
    input  wire                            AP_AXIMM_11_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_11_AWADDR,
    output wire [7:0]                      M_AXIMM_11_AWLEN,
    output wire [2:0]                      M_AXIMM_11_AWSIZE,
    output wire [1:0]                      M_AXIMM_11_AWBURST,
    output wire [1:0]                      M_AXIMM_11_AWLOCK,
    output wire [3:0]                      M_AXIMM_11_AWCACHE,
    output wire [2:0]                      M_AXIMM_11_AWPROT,
    output wire [3:0]                      M_AXIMM_11_AWREGION,
    output wire [3:0]                      M_AXIMM_11_AWQOS,
    output wire                            M_AXIMM_11_AWVALID,
    input  wire                            M_AXIMM_11_AWREADY,
    output wire [M_AXIMM_11_DATA_WIDTH-1:0]   M_AXIMM_11_WDATA,
    output wire [M_AXIMM_11_DATA_WIDTH/8-1:0] M_AXIMM_11_WSTRB,
    output wire                            M_AXIMM_11_WLAST,
    output wire                            M_AXIMM_11_WVALID,
    input  wire                            M_AXIMM_11_WREADY,
    input  wire [1:0]                      M_AXIMM_11_BRESP,
    input  wire                            M_AXIMM_11_BVALID,
    output wire                            M_AXIMM_11_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_11_ARADDR,
    output wire [7:0]                      M_AXIMM_11_ARLEN,
    output wire [2:0]                      M_AXIMM_11_ARSIZE,
    output wire [1:0]                      M_AXIMM_11_ARBURST,
    output wire [1:0]                      M_AXIMM_11_ARLOCK,
    output wire [3:0]                      M_AXIMM_11_ARCACHE,
    output wire [2:0]                      M_AXIMM_11_ARPROT,
    output wire [3:0]                      M_AXIMM_11_ARREGION,
    output wire [3:0]                      M_AXIMM_11_ARQOS,
    output wire                            M_AXIMM_11_ARVALID,
    input  wire                            M_AXIMM_11_ARREADY,
    input  wire [M_AXIMM_11_DATA_WIDTH-1:0]   M_AXIMM_11_RDATA,
    input  wire [1:0]                      M_AXIMM_11_RRESP,
    input  wire                            M_AXIMM_11_RLAST,
    input  wire                            M_AXIMM_11_RVALID,
    output wire                            M_AXIMM_11_RREADY,
    //AXI-MM pass-through interface 12
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_12_AWADDR,
    input wire [7:0]                      AP_AXIMM_12_AWLEN,
    input wire [2:0]                      AP_AXIMM_12_AWSIZE,
    input wire [1:0]                      AP_AXIMM_12_AWBURST,
    input wire [1:0]                      AP_AXIMM_12_AWLOCK,
    input wire [3:0]                      AP_AXIMM_12_AWCACHE,
    input wire [2:0]                      AP_AXIMM_12_AWPROT,
    input wire [3:0]                      AP_AXIMM_12_AWREGION,
    input wire [3:0]                      AP_AXIMM_12_AWQOS,
    input wire                            AP_AXIMM_12_AWVALID,
    output  wire                            AP_AXIMM_12_AWREADY,
    input wire [M_AXIMM_12_DATA_WIDTH-1:0]   AP_AXIMM_12_WDATA,
    input wire [M_AXIMM_12_DATA_WIDTH/8-1:0] AP_AXIMM_12_WSTRB,
    input wire                            AP_AXIMM_12_WLAST,
    input wire                            AP_AXIMM_12_WVALID,
    output  wire                            AP_AXIMM_12_WREADY,
    output  wire [1:0]                      AP_AXIMM_12_BRESP,
    output  wire                            AP_AXIMM_12_BVALID,
    input wire                            AP_AXIMM_12_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_12_ARADDR,
    input wire [7:0]                      AP_AXIMM_12_ARLEN,
    input wire [2:0]                      AP_AXIMM_12_ARSIZE,
    input wire [1:0]                      AP_AXIMM_12_ARBURST,
    input wire [1:0]                      AP_AXIMM_12_ARLOCK,
    input wire [3:0]                      AP_AXIMM_12_ARCACHE,
    input wire [2:0]                      AP_AXIMM_12_ARPROT,
    input wire [3:0]                      AP_AXIMM_12_ARREGION,
    input wire [3:0]                      AP_AXIMM_12_ARQOS,
    input wire                            AP_AXIMM_12_ARVALID,
    output  wire                            AP_AXIMM_12_ARREADY,
    output  wire [M_AXIMM_12_DATA_WIDTH-1:0]   AP_AXIMM_12_RDATA,
    output  wire [1:0]                      AP_AXIMM_12_RRESP,
    output  wire                            AP_AXIMM_12_RLAST,
    output  wire                            AP_AXIMM_12_RVALID,
    input  wire                            AP_AXIMM_12_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_12_AWADDR,
    output wire [7:0]                      M_AXIMM_12_AWLEN,
    output wire [2:0]                      M_AXIMM_12_AWSIZE,
    output wire [1:0]                      M_AXIMM_12_AWBURST,
    output wire [1:0]                      M_AXIMM_12_AWLOCK,
    output wire [3:0]                      M_AXIMM_12_AWCACHE,
    output wire [2:0]                      M_AXIMM_12_AWPROT,
    output wire [3:0]                      M_AXIMM_12_AWREGION,
    output wire [3:0]                      M_AXIMM_12_AWQOS,
    output wire                            M_AXIMM_12_AWVALID,
    input  wire                            M_AXIMM_12_AWREADY,
    output wire [M_AXIMM_12_DATA_WIDTH-1:0]   M_AXIMM_12_WDATA,
    output wire [M_AXIMM_12_DATA_WIDTH/8-1:0] M_AXIMM_12_WSTRB,
    output wire                            M_AXIMM_12_WLAST,
    output wire                            M_AXIMM_12_WVALID,
    input  wire                            M_AXIMM_12_WREADY,
    input  wire [1:0]                      M_AXIMM_12_BRESP,
    input  wire                            M_AXIMM_12_BVALID,
    output wire                            M_AXIMM_12_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_12_ARADDR,
    output wire [7:0]                      M_AXIMM_12_ARLEN,
    output wire [2:0]                      M_AXIMM_12_ARSIZE,
    output wire [1:0]                      M_AXIMM_12_ARBURST,
    output wire [1:0]                      M_AXIMM_12_ARLOCK,
    output wire [3:0]                      M_AXIMM_12_ARCACHE,
    output wire [2:0]                      M_AXIMM_12_ARPROT,
    output wire [3:0]                      M_AXIMM_12_ARREGION,
    output wire [3:0]                      M_AXIMM_12_ARQOS,
    output wire                            M_AXIMM_12_ARVALID,
    input  wire                            M_AXIMM_12_ARREADY,
    input  wire [M_AXIMM_12_DATA_WIDTH-1:0]   M_AXIMM_12_RDATA,
    input  wire [1:0]                      M_AXIMM_12_RRESP,
    input  wire                            M_AXIMM_12_RLAST,
    input  wire                            M_AXIMM_12_RVALID,
    output wire                            M_AXIMM_12_RREADY,
    //AXI-MM pass-through interface 13
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_13_AWADDR,
    input wire [7:0]                      AP_AXIMM_13_AWLEN,
    input wire [2:0]                      AP_AXIMM_13_AWSIZE,
    input wire [1:0]                      AP_AXIMM_13_AWBURST,
    input wire [1:0]                      AP_AXIMM_13_AWLOCK,
    input wire [3:0]                      AP_AXIMM_13_AWCACHE,
    input wire [2:0]                      AP_AXIMM_13_AWPROT,
    input wire [3:0]                      AP_AXIMM_13_AWREGION,
    input wire [3:0]                      AP_AXIMM_13_AWQOS,
    input wire                            AP_AXIMM_13_AWVALID,
    output  wire                            AP_AXIMM_13_AWREADY,
    input wire [M_AXIMM_13_DATA_WIDTH-1:0]   AP_AXIMM_13_WDATA,
    input wire [M_AXIMM_13_DATA_WIDTH/8-1:0] AP_AXIMM_13_WSTRB,
    input wire                            AP_AXIMM_13_WLAST,
    input wire                            AP_AXIMM_13_WVALID,
    output  wire                            AP_AXIMM_13_WREADY,
    output  wire [1:0]                      AP_AXIMM_13_BRESP,
    output  wire                            AP_AXIMM_13_BVALID,
    input wire                            AP_AXIMM_13_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_13_ARADDR,
    input wire [7:0]                      AP_AXIMM_13_ARLEN,
    input wire [2:0]                      AP_AXIMM_13_ARSIZE,
    input wire [1:0]                      AP_AXIMM_13_ARBURST,
    input wire [1:0]                      AP_AXIMM_13_ARLOCK,
    input wire [3:0]                      AP_AXIMM_13_ARCACHE,
    input wire [2:0]                      AP_AXIMM_13_ARPROT,
    input wire [3:0]                      AP_AXIMM_13_ARREGION,
    input wire [3:0]                      AP_AXIMM_13_ARQOS,
    input wire                            AP_AXIMM_13_ARVALID,
    output  wire                            AP_AXIMM_13_ARREADY,
    output  wire [M_AXIMM_13_DATA_WIDTH-1:0]   AP_AXIMM_13_RDATA,
    output  wire [1:0]                      AP_AXIMM_13_RRESP,
    output  wire                            AP_AXIMM_13_RLAST,
    output  wire                            AP_AXIMM_13_RVALID,
    input  wire                            AP_AXIMM_13_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_13_AWADDR,
    output wire [7:0]                      M_AXIMM_13_AWLEN,
    output wire [2:0]                      M_AXIMM_13_AWSIZE,
    output wire [1:0]                      M_AXIMM_13_AWBURST,
    output wire [1:0]                      M_AXIMM_13_AWLOCK,
    output wire [3:0]                      M_AXIMM_13_AWCACHE,
    output wire [2:0]                      M_AXIMM_13_AWPROT,
    output wire [3:0]                      M_AXIMM_13_AWREGION,
    output wire [3:0]                      M_AXIMM_13_AWQOS,
    output wire                            M_AXIMM_13_AWVALID,
    input  wire                            M_AXIMM_13_AWREADY,
    output wire [M_AXIMM_13_DATA_WIDTH-1:0]   M_AXIMM_13_WDATA,
    output wire [M_AXIMM_13_DATA_WIDTH/8-1:0] M_AXIMM_13_WSTRB,
    output wire                            M_AXIMM_13_WLAST,
    output wire                            M_AXIMM_13_WVALID,
    input  wire                            M_AXIMM_13_WREADY,
    input  wire [1:0]                      M_AXIMM_13_BRESP,
    input  wire                            M_AXIMM_13_BVALID,
    output wire                            M_AXIMM_13_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_13_ARADDR,
    output wire [7:0]                      M_AXIMM_13_ARLEN,
    output wire [2:0]                      M_AXIMM_13_ARSIZE,
    output wire [1:0]                      M_AXIMM_13_ARBURST,
    output wire [1:0]                      M_AXIMM_13_ARLOCK,
    output wire [3:0]                      M_AXIMM_13_ARCACHE,
    output wire [2:0]                      M_AXIMM_13_ARPROT,
    output wire [3:0]                      M_AXIMM_13_ARREGION,
    output wire [3:0]                      M_AXIMM_13_ARQOS,
    output wire                            M_AXIMM_13_ARVALID,
    input  wire                            M_AXIMM_13_ARREADY,
    input  wire [M_AXIMM_13_DATA_WIDTH-1:0]   M_AXIMM_13_RDATA,
    input  wire [1:0]                      M_AXIMM_13_RRESP,
    input  wire                            M_AXIMM_13_RLAST,
    input  wire                            M_AXIMM_13_RVALID,
    output wire                            M_AXIMM_13_RREADY,
    //AXI-MM pass-through interface 14
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_14_AWADDR,
    input wire [7:0]                      AP_AXIMM_14_AWLEN,
    input wire [2:0]                      AP_AXIMM_14_AWSIZE,
    input wire [1:0]                      AP_AXIMM_14_AWBURST,
    input wire [1:0]                      AP_AXIMM_14_AWLOCK,
    input wire [3:0]                      AP_AXIMM_14_AWCACHE,
    input wire [2:0]                      AP_AXIMM_14_AWPROT,
    input wire [3:0]                      AP_AXIMM_14_AWREGION,
    input wire [3:0]                      AP_AXIMM_14_AWQOS,
    input wire                            AP_AXIMM_14_AWVALID,
    output  wire                            AP_AXIMM_14_AWREADY,
    input wire [M_AXIMM_14_DATA_WIDTH-1:0]   AP_AXIMM_14_WDATA,
    input wire [M_AXIMM_14_DATA_WIDTH/8-1:0] AP_AXIMM_14_WSTRB,
    input wire                            AP_AXIMM_14_WLAST,
    input wire                            AP_AXIMM_14_WVALID,
    output  wire                            AP_AXIMM_14_WREADY,
    output  wire [1:0]                      AP_AXIMM_14_BRESP,
    output  wire                            AP_AXIMM_14_BVALID,
    input wire                            AP_AXIMM_14_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_14_ARADDR,
    input wire [7:0]                      AP_AXIMM_14_ARLEN,
    input wire [2:0]                      AP_AXIMM_14_ARSIZE,
    input wire [1:0]                      AP_AXIMM_14_ARBURST,
    input wire [1:0]                      AP_AXIMM_14_ARLOCK,
    input wire [3:0]                      AP_AXIMM_14_ARCACHE,
    input wire [2:0]                      AP_AXIMM_14_ARPROT,
    input wire [3:0]                      AP_AXIMM_14_ARREGION,
    input wire [3:0]                      AP_AXIMM_14_ARQOS,
    input wire                            AP_AXIMM_14_ARVALID,
    output  wire                            AP_AXIMM_14_ARREADY,
    output  wire [M_AXIMM_14_DATA_WIDTH-1:0]   AP_AXIMM_14_RDATA,
    output  wire [1:0]                      AP_AXIMM_14_RRESP,
    output  wire                            AP_AXIMM_14_RLAST,
    output  wire                            AP_AXIMM_14_RVALID,
    input  wire                            AP_AXIMM_14_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_14_AWADDR,
    output wire [7:0]                      M_AXIMM_14_AWLEN,
    output wire [2:0]                      M_AXIMM_14_AWSIZE,
    output wire [1:0]                      M_AXIMM_14_AWBURST,
    output wire [1:0]                      M_AXIMM_14_AWLOCK,
    output wire [3:0]                      M_AXIMM_14_AWCACHE,
    output wire [2:0]                      M_AXIMM_14_AWPROT,
    output wire [3:0]                      M_AXIMM_14_AWREGION,
    output wire [3:0]                      M_AXIMM_14_AWQOS,
    output wire                            M_AXIMM_14_AWVALID,
    input  wire                            M_AXIMM_14_AWREADY,
    output wire [M_AXIMM_14_DATA_WIDTH-1:0]   M_AXIMM_14_WDATA,
    output wire [M_AXIMM_14_DATA_WIDTH/8-1:0] M_AXIMM_14_WSTRB,
    output wire                            M_AXIMM_14_WLAST,
    output wire                            M_AXIMM_14_WVALID,
    input  wire                            M_AXIMM_14_WREADY,
    input  wire [1:0]                      M_AXIMM_14_BRESP,
    input  wire                            M_AXIMM_14_BVALID,
    output wire                            M_AXIMM_14_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_14_ARADDR,
    output wire [7:0]                      M_AXIMM_14_ARLEN,
    output wire [2:0]                      M_AXIMM_14_ARSIZE,
    output wire [1:0]                      M_AXIMM_14_ARBURST,
    output wire [1:0]                      M_AXIMM_14_ARLOCK,
    output wire [3:0]                      M_AXIMM_14_ARCACHE,
    output wire [2:0]                      M_AXIMM_14_ARPROT,
    output wire [3:0]                      M_AXIMM_14_ARREGION,
    output wire [3:0]                      M_AXIMM_14_ARQOS,
    output wire                            M_AXIMM_14_ARVALID,
    input  wire                            M_AXIMM_14_ARREADY,
    input  wire [M_AXIMM_14_DATA_WIDTH-1:0]   M_AXIMM_14_RDATA,
    input  wire [1:0]                      M_AXIMM_14_RRESP,
    input  wire                            M_AXIMM_14_RLAST,
    input  wire                            M_AXIMM_14_RVALID,
    output wire                            M_AXIMM_14_RREADY,
    //AXI-MM pass-through interface 15
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_15_AWADDR,
    input wire [7:0]                      AP_AXIMM_15_AWLEN,
    input wire [2:0]                      AP_AXIMM_15_AWSIZE,
    input wire [1:0]                      AP_AXIMM_15_AWBURST,
    input wire [1:0]                      AP_AXIMM_15_AWLOCK,
    input wire [3:0]                      AP_AXIMM_15_AWCACHE,
    input wire [2:0]                      AP_AXIMM_15_AWPROT,
    input wire [3:0]                      AP_AXIMM_15_AWREGION,
    input wire [3:0]                      AP_AXIMM_15_AWQOS,
    input wire                            AP_AXIMM_15_AWVALID,
    output  wire                            AP_AXIMM_15_AWREADY,
    input wire [M_AXIMM_15_DATA_WIDTH-1:0]   AP_AXIMM_15_WDATA,
    input wire [M_AXIMM_15_DATA_WIDTH/8-1:0] AP_AXIMM_15_WSTRB,
    input wire                            AP_AXIMM_15_WLAST,
    input wire                            AP_AXIMM_15_WVALID,
    output  wire                            AP_AXIMM_15_WREADY,
    output  wire [1:0]                      AP_AXIMM_15_BRESP,
    output  wire                            AP_AXIMM_15_BVALID,
    input wire                            AP_AXIMM_15_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_15_ARADDR,
    input wire [7:0]                      AP_AXIMM_15_ARLEN,
    input wire [2:0]                      AP_AXIMM_15_ARSIZE,
    input wire [1:0]                      AP_AXIMM_15_ARBURST,
    input wire [1:0]                      AP_AXIMM_15_ARLOCK,
    input wire [3:0]                      AP_AXIMM_15_ARCACHE,
    input wire [2:0]                      AP_AXIMM_15_ARPROT,
    input wire [3:0]                      AP_AXIMM_15_ARREGION,
    input wire [3:0]                      AP_AXIMM_15_ARQOS,
    input wire                            AP_AXIMM_15_ARVALID,
    output  wire                            AP_AXIMM_15_ARREADY,
    output  wire [M_AXIMM_15_DATA_WIDTH-1:0]   AP_AXIMM_15_RDATA,
    output  wire [1:0]                      AP_AXIMM_15_RRESP,
    output  wire                            AP_AXIMM_15_RLAST,
    output  wire                            AP_AXIMM_15_RVALID,
    input  wire                            AP_AXIMM_15_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_15_AWADDR,
    output wire [7:0]                      M_AXIMM_15_AWLEN,
    output wire [2:0]                      M_AXIMM_15_AWSIZE,
    output wire [1:0]                      M_AXIMM_15_AWBURST,
    output wire [1:0]                      M_AXIMM_15_AWLOCK,
    output wire [3:0]                      M_AXIMM_15_AWCACHE,
    output wire [2:0]                      M_AXIMM_15_AWPROT,
    output wire [3:0]                      M_AXIMM_15_AWREGION,
    output wire [3:0]                      M_AXIMM_15_AWQOS,
    output wire                            M_AXIMM_15_AWVALID,
    input  wire                            M_AXIMM_15_AWREADY,
    output wire [M_AXIMM_15_DATA_WIDTH-1:0]   M_AXIMM_15_WDATA,
    output wire [M_AXIMM_15_DATA_WIDTH/8-1:0] M_AXIMM_15_WSTRB,
    output wire                            M_AXIMM_15_WLAST,
    output wire                            M_AXIMM_15_WVALID,
    input  wire                            M_AXIMM_15_WREADY,
    input  wire [1:0]                      M_AXIMM_15_BRESP,
    input  wire                            M_AXIMM_15_BVALID,
    output wire                            M_AXIMM_15_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_15_ARADDR,
    output wire [7:0]                      M_AXIMM_15_ARLEN,
    output wire [2:0]                      M_AXIMM_15_ARSIZE,
    output wire [1:0]                      M_AXIMM_15_ARBURST,
    output wire [1:0]                      M_AXIMM_15_ARLOCK,
    output wire [3:0]                      M_AXIMM_15_ARCACHE,
    output wire [2:0]                      M_AXIMM_15_ARPROT,
    output wire [3:0]                      M_AXIMM_15_ARREGION,
    output wire [3:0]                      M_AXIMM_15_ARQOS,
    output wire                            M_AXIMM_15_ARVALID,
    input  wire                            M_AXIMM_15_ARREADY,
    input  wire [M_AXIMM_15_DATA_WIDTH-1:0]   M_AXIMM_15_RDATA,
    input  wire [1:0]                      M_AXIMM_15_RRESP,
    input  wire                            M_AXIMM_15_RLAST,
    input  wire                            M_AXIMM_15_RVALID,
    output wire                            M_AXIMM_15_RREADY,
    //AXI-MM pass-through interface 16
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_16_AWADDR,
    input wire [7:0]                      AP_AXIMM_16_AWLEN,
    input wire [2:0]                      AP_AXIMM_16_AWSIZE,
    input wire [1:0]                      AP_AXIMM_16_AWBURST,
    input wire [1:0]                      AP_AXIMM_16_AWLOCK,
    input wire [3:0]                      AP_AXIMM_16_AWCACHE,
    input wire [2:0]                      AP_AXIMM_16_AWPROT,
    input wire [3:0]                      AP_AXIMM_16_AWREGION,
    input wire [3:0]                      AP_AXIMM_16_AWQOS,
    input wire                            AP_AXIMM_16_AWVALID,
    output  wire                            AP_AXIMM_16_AWREADY,
    input wire [M_AXIMM_16_DATA_WIDTH-1:0]   AP_AXIMM_16_WDATA,
    input wire [M_AXIMM_16_DATA_WIDTH/8-1:0] AP_AXIMM_16_WSTRB,
    input wire                            AP_AXIMM_16_WLAST,
    input wire                            AP_AXIMM_16_WVALID,
    output  wire                            AP_AXIMM_16_WREADY,
    output  wire [1:0]                      AP_AXIMM_16_BRESP,
    output  wire                            AP_AXIMM_16_BVALID,
    input wire                            AP_AXIMM_16_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_16_ARADDR,
    input wire [7:0]                      AP_AXIMM_16_ARLEN,
    input wire [2:0]                      AP_AXIMM_16_ARSIZE,
    input wire [1:0]                      AP_AXIMM_16_ARBURST,
    input wire [1:0]                      AP_AXIMM_16_ARLOCK,
    input wire [3:0]                      AP_AXIMM_16_ARCACHE,
    input wire [2:0]                      AP_AXIMM_16_ARPROT,
    input wire [3:0]                      AP_AXIMM_16_ARREGION,
    input wire [3:0]                      AP_AXIMM_16_ARQOS,
    input wire                            AP_AXIMM_16_ARVALID,
    output  wire                            AP_AXIMM_16_ARREADY,
    output  wire [M_AXIMM_16_DATA_WIDTH-1:0]   AP_AXIMM_16_RDATA,
    output  wire [1:0]                      AP_AXIMM_16_RRESP,
    output  wire                            AP_AXIMM_16_RLAST,
    output  wire                            AP_AXIMM_16_RVALID,
    input  wire                            AP_AXIMM_16_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_16_AWADDR,
    output wire [7:0]                      M_AXIMM_16_AWLEN,
    output wire [2:0]                      M_AXIMM_16_AWSIZE,
    output wire [1:0]                      M_AXIMM_16_AWBURST,
    output wire [1:0]                      M_AXIMM_16_AWLOCK,
    output wire [3:0]                      M_AXIMM_16_AWCACHE,
    output wire [2:0]                      M_AXIMM_16_AWPROT,
    output wire [3:0]                      M_AXIMM_16_AWREGION,
    output wire [3:0]                      M_AXIMM_16_AWQOS,
    output wire                            M_AXIMM_16_AWVALID,
    input  wire                            M_AXIMM_16_AWREADY,
    output wire [M_AXIMM_16_DATA_WIDTH-1:0]   M_AXIMM_16_WDATA,
    output wire [M_AXIMM_16_DATA_WIDTH/8-1:0] M_AXIMM_16_WSTRB,
    output wire                            M_AXIMM_16_WLAST,
    output wire                            M_AXIMM_16_WVALID,
    input  wire                            M_AXIMM_16_WREADY,
    input  wire [1:0]                      M_AXIMM_16_BRESP,
    input  wire                            M_AXIMM_16_BVALID,
    output wire                            M_AXIMM_16_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_16_ARADDR,
    output wire [7:0]                      M_AXIMM_16_ARLEN,
    output wire [2:0]                      M_AXIMM_16_ARSIZE,
    output wire [1:0]                      M_AXIMM_16_ARBURST,
    output wire [1:0]                      M_AXIMM_16_ARLOCK,
    output wire [3:0]                      M_AXIMM_16_ARCACHE,
    output wire [2:0]                      M_AXIMM_16_ARPROT,
    output wire [3:0]                      M_AXIMM_16_ARREGION,
    output wire [3:0]                      M_AXIMM_16_ARQOS,
    output wire                            M_AXIMM_16_ARVALID,
    input  wire                            M_AXIMM_16_ARREADY,
    input  wire [M_AXIMM_16_DATA_WIDTH-1:0]   M_AXIMM_16_RDATA,
    input  wire [1:0]                      M_AXIMM_16_RRESP,
    input  wire                            M_AXIMM_16_RLAST,
    input  wire                            M_AXIMM_16_RVALID,
    output wire                            M_AXIMM_16_RREADY,
    //AXI-MM pass-through interface 17
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_17_AWADDR,
    input wire [7:0]                      AP_AXIMM_17_AWLEN,
    input wire [2:0]                      AP_AXIMM_17_AWSIZE,
    input wire [1:0]                      AP_AXIMM_17_AWBURST,
    input wire [1:0]                      AP_AXIMM_17_AWLOCK,
    input wire [3:0]                      AP_AXIMM_17_AWCACHE,
    input wire [2:0]                      AP_AXIMM_17_AWPROT,
    input wire [3:0]                      AP_AXIMM_17_AWREGION,
    input wire [3:0]                      AP_AXIMM_17_AWQOS,
    input wire                            AP_AXIMM_17_AWVALID,
    output  wire                            AP_AXIMM_17_AWREADY,
    input wire [M_AXIMM_17_DATA_WIDTH-1:0]   AP_AXIMM_17_WDATA,
    input wire [M_AXIMM_17_DATA_WIDTH/8-1:0] AP_AXIMM_17_WSTRB,
    input wire                            AP_AXIMM_17_WLAST,
    input wire                            AP_AXIMM_17_WVALID,
    output  wire                            AP_AXIMM_17_WREADY,
    output  wire [1:0]                      AP_AXIMM_17_BRESP,
    output  wire                            AP_AXIMM_17_BVALID,
    input wire                            AP_AXIMM_17_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_17_ARADDR,
    input wire [7:0]                      AP_AXIMM_17_ARLEN,
    input wire [2:0]                      AP_AXIMM_17_ARSIZE,
    input wire [1:0]                      AP_AXIMM_17_ARBURST,
    input wire [1:0]                      AP_AXIMM_17_ARLOCK,
    input wire [3:0]                      AP_AXIMM_17_ARCACHE,
    input wire [2:0]                      AP_AXIMM_17_ARPROT,
    input wire [3:0]                      AP_AXIMM_17_ARREGION,
    input wire [3:0]                      AP_AXIMM_17_ARQOS,
    input wire                            AP_AXIMM_17_ARVALID,
    output  wire                            AP_AXIMM_17_ARREADY,
    output  wire [M_AXIMM_17_DATA_WIDTH-1:0]   AP_AXIMM_17_RDATA,
    output  wire [1:0]                      AP_AXIMM_17_RRESP,
    output  wire                            AP_AXIMM_17_RLAST,
    output  wire                            AP_AXIMM_17_RVALID,
    input  wire                            AP_AXIMM_17_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_17_AWADDR,
    output wire [7:0]                      M_AXIMM_17_AWLEN,
    output wire [2:0]                      M_AXIMM_17_AWSIZE,
    output wire [1:0]                      M_AXIMM_17_AWBURST,
    output wire [1:0]                      M_AXIMM_17_AWLOCK,
    output wire [3:0]                      M_AXIMM_17_AWCACHE,
    output wire [2:0]                      M_AXIMM_17_AWPROT,
    output wire [3:0]                      M_AXIMM_17_AWREGION,
    output wire [3:0]                      M_AXIMM_17_AWQOS,
    output wire                            M_AXIMM_17_AWVALID,
    input  wire                            M_AXIMM_17_AWREADY,
    output wire [M_AXIMM_17_DATA_WIDTH-1:0]   M_AXIMM_17_WDATA,
    output wire [M_AXIMM_17_DATA_WIDTH/8-1:0] M_AXIMM_17_WSTRB,
    output wire                            M_AXIMM_17_WLAST,
    output wire                            M_AXIMM_17_WVALID,
    input  wire                            M_AXIMM_17_WREADY,
    input  wire [1:0]                      M_AXIMM_17_BRESP,
    input  wire                            M_AXIMM_17_BVALID,
    output wire                            M_AXIMM_17_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_17_ARADDR,
    output wire [7:0]                      M_AXIMM_17_ARLEN,
    output wire [2:0]                      M_AXIMM_17_ARSIZE,
    output wire [1:0]                      M_AXIMM_17_ARBURST,
    output wire [1:0]                      M_AXIMM_17_ARLOCK,
    output wire [3:0]                      M_AXIMM_17_ARCACHE,
    output wire [2:0]                      M_AXIMM_17_ARPROT,
    output wire [3:0]                      M_AXIMM_17_ARREGION,
    output wire [3:0]                      M_AXIMM_17_ARQOS,
    output wire                            M_AXIMM_17_ARVALID,
    input  wire                            M_AXIMM_17_ARREADY,
    input  wire [M_AXIMM_17_DATA_WIDTH-1:0]   M_AXIMM_17_RDATA,
    input  wire [1:0]                      M_AXIMM_17_RRESP,
    input  wire                            M_AXIMM_17_RLAST,
    input  wire                            M_AXIMM_17_RVALID,
    output wire                            M_AXIMM_17_RREADY,
    //AXI-MM pass-through interface 18
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_18_AWADDR,
    input wire [7:0]                      AP_AXIMM_18_AWLEN,
    input wire [2:0]                      AP_AXIMM_18_AWSIZE,
    input wire [1:0]                      AP_AXIMM_18_AWBURST,
    input wire [1:0]                      AP_AXIMM_18_AWLOCK,
    input wire [3:0]                      AP_AXIMM_18_AWCACHE,
    input wire [2:0]                      AP_AXIMM_18_AWPROT,
    input wire [3:0]                      AP_AXIMM_18_AWREGION,
    input wire [3:0]                      AP_AXIMM_18_AWQOS,
    input wire                            AP_AXIMM_18_AWVALID,
    output  wire                            AP_AXIMM_18_AWREADY,
    input wire [M_AXIMM_18_DATA_WIDTH-1:0]   AP_AXIMM_18_WDATA,
    input wire [M_AXIMM_18_DATA_WIDTH/8-1:0] AP_AXIMM_18_WSTRB,
    input wire                            AP_AXIMM_18_WLAST,
    input wire                            AP_AXIMM_18_WVALID,
    output  wire                            AP_AXIMM_18_WREADY,
    output  wire [1:0]                      AP_AXIMM_18_BRESP,
    output  wire                            AP_AXIMM_18_BVALID,
    input wire                            AP_AXIMM_18_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_18_ARADDR,
    input wire [7:0]                      AP_AXIMM_18_ARLEN,
    input wire [2:0]                      AP_AXIMM_18_ARSIZE,
    input wire [1:0]                      AP_AXIMM_18_ARBURST,
    input wire [1:0]                      AP_AXIMM_18_ARLOCK,
    input wire [3:0]                      AP_AXIMM_18_ARCACHE,
    input wire [2:0]                      AP_AXIMM_18_ARPROT,
    input wire [3:0]                      AP_AXIMM_18_ARREGION,
    input wire [3:0]                      AP_AXIMM_18_ARQOS,
    input wire                            AP_AXIMM_18_ARVALID,
    output  wire                            AP_AXIMM_18_ARREADY,
    output  wire [M_AXIMM_18_DATA_WIDTH-1:0]   AP_AXIMM_18_RDATA,
    output  wire [1:0]                      AP_AXIMM_18_RRESP,
    output  wire                            AP_AXIMM_18_RLAST,
    output  wire                            AP_AXIMM_18_RVALID,
    input  wire                            AP_AXIMM_18_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_18_AWADDR,
    output wire [7:0]                      M_AXIMM_18_AWLEN,
    output wire [2:0]                      M_AXIMM_18_AWSIZE,
    output wire [1:0]                      M_AXIMM_18_AWBURST,
    output wire [1:0]                      M_AXIMM_18_AWLOCK,
    output wire [3:0]                      M_AXIMM_18_AWCACHE,
    output wire [2:0]                      M_AXIMM_18_AWPROT,
    output wire [3:0]                      M_AXIMM_18_AWREGION,
    output wire [3:0]                      M_AXIMM_18_AWQOS,
    output wire                            M_AXIMM_18_AWVALID,
    input  wire                            M_AXIMM_18_AWREADY,
    output wire [M_AXIMM_18_DATA_WIDTH-1:0]   M_AXIMM_18_WDATA,
    output wire [M_AXIMM_18_DATA_WIDTH/8-1:0] M_AXIMM_18_WSTRB,
    output wire                            M_AXIMM_18_WLAST,
    output wire                            M_AXIMM_18_WVALID,
    input  wire                            M_AXIMM_18_WREADY,
    input  wire [1:0]                      M_AXIMM_18_BRESP,
    input  wire                            M_AXIMM_18_BVALID,
    output wire                            M_AXIMM_18_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_18_ARADDR,
    output wire [7:0]                      M_AXIMM_18_ARLEN,
    output wire [2:0]                      M_AXIMM_18_ARSIZE,
    output wire [1:0]                      M_AXIMM_18_ARBURST,
    output wire [1:0]                      M_AXIMM_18_ARLOCK,
    output wire [3:0]                      M_AXIMM_18_ARCACHE,
    output wire [2:0]                      M_AXIMM_18_ARPROT,
    output wire [3:0]                      M_AXIMM_18_ARREGION,
    output wire [3:0]                      M_AXIMM_18_ARQOS,
    output wire                            M_AXIMM_18_ARVALID,
    input  wire                            M_AXIMM_18_ARREADY,
    input  wire [M_AXIMM_18_DATA_WIDTH-1:0]   M_AXIMM_18_RDATA,
    input  wire [1:0]                      M_AXIMM_18_RRESP,
    input  wire                            M_AXIMM_18_RLAST,
    input  wire                            M_AXIMM_18_RVALID,
    output wire                            M_AXIMM_18_RREADY,
    //AXI-MM pass-through interface 19
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_19_AWADDR,
    input wire [7:0]                      AP_AXIMM_19_AWLEN,
    input wire [2:0]                      AP_AXIMM_19_AWSIZE,
    input wire [1:0]                      AP_AXIMM_19_AWBURST,
    input wire [1:0]                      AP_AXIMM_19_AWLOCK,
    input wire [3:0]                      AP_AXIMM_19_AWCACHE,
    input wire [2:0]                      AP_AXIMM_19_AWPROT,
    input wire [3:0]                      AP_AXIMM_19_AWREGION,
    input wire [3:0]                      AP_AXIMM_19_AWQOS,
    input wire                            AP_AXIMM_19_AWVALID,
    output  wire                            AP_AXIMM_19_AWREADY,
    input wire [M_AXIMM_19_DATA_WIDTH-1:0]   AP_AXIMM_19_WDATA,
    input wire [M_AXIMM_19_DATA_WIDTH/8-1:0] AP_AXIMM_19_WSTRB,
    input wire                            AP_AXIMM_19_WLAST,
    input wire                            AP_AXIMM_19_WVALID,
    output  wire                            AP_AXIMM_19_WREADY,
    output  wire [1:0]                      AP_AXIMM_19_BRESP,
    output  wire                            AP_AXIMM_19_BVALID,
    input wire                            AP_AXIMM_19_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_19_ARADDR,
    input wire [7:0]                      AP_AXIMM_19_ARLEN,
    input wire [2:0]                      AP_AXIMM_19_ARSIZE,
    input wire [1:0]                      AP_AXIMM_19_ARBURST,
    input wire [1:0]                      AP_AXIMM_19_ARLOCK,
    input wire [3:0]                      AP_AXIMM_19_ARCACHE,
    input wire [2:0]                      AP_AXIMM_19_ARPROT,
    input wire [3:0]                      AP_AXIMM_19_ARREGION,
    input wire [3:0]                      AP_AXIMM_19_ARQOS,
    input wire                            AP_AXIMM_19_ARVALID,
    output  wire                            AP_AXIMM_19_ARREADY,
    output  wire [M_AXIMM_19_DATA_WIDTH-1:0]   AP_AXIMM_19_RDATA,
    output  wire [1:0]                      AP_AXIMM_19_RRESP,
    output  wire                            AP_AXIMM_19_RLAST,
    output  wire                            AP_AXIMM_19_RVALID,
    input  wire                            AP_AXIMM_19_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_19_AWADDR,
    output wire [7:0]                      M_AXIMM_19_AWLEN,
    output wire [2:0]                      M_AXIMM_19_AWSIZE,
    output wire [1:0]                      M_AXIMM_19_AWBURST,
    output wire [1:0]                      M_AXIMM_19_AWLOCK,
    output wire [3:0]                      M_AXIMM_19_AWCACHE,
    output wire [2:0]                      M_AXIMM_19_AWPROT,
    output wire [3:0]                      M_AXIMM_19_AWREGION,
    output wire [3:0]                      M_AXIMM_19_AWQOS,
    output wire                            M_AXIMM_19_AWVALID,
    input  wire                            M_AXIMM_19_AWREADY,
    output wire [M_AXIMM_19_DATA_WIDTH-1:0]   M_AXIMM_19_WDATA,
    output wire [M_AXIMM_19_DATA_WIDTH/8-1:0] M_AXIMM_19_WSTRB,
    output wire                            M_AXIMM_19_WLAST,
    output wire                            M_AXIMM_19_WVALID,
    input  wire                            M_AXIMM_19_WREADY,
    input  wire [1:0]                      M_AXIMM_19_BRESP,
    input  wire                            M_AXIMM_19_BVALID,
    output wire                            M_AXIMM_19_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_19_ARADDR,
    output wire [7:0]                      M_AXIMM_19_ARLEN,
    output wire [2:0]                      M_AXIMM_19_ARSIZE,
    output wire [1:0]                      M_AXIMM_19_ARBURST,
    output wire [1:0]                      M_AXIMM_19_ARLOCK,
    output wire [3:0]                      M_AXIMM_19_ARCACHE,
    output wire [2:0]                      M_AXIMM_19_ARPROT,
    output wire [3:0]                      M_AXIMM_19_ARREGION,
    output wire [3:0]                      M_AXIMM_19_ARQOS,
    output wire                            M_AXIMM_19_ARVALID,
    input  wire                            M_AXIMM_19_ARREADY,
    input  wire [M_AXIMM_19_DATA_WIDTH-1:0]   M_AXIMM_19_RDATA,
    input  wire [1:0]                      M_AXIMM_19_RRESP,
    input  wire                            M_AXIMM_19_RLAST,
    input  wire                            M_AXIMM_19_RVALID,
    output wire                            M_AXIMM_19_RREADY,
    //AXI-MM pass-through interface 20
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_20_AWADDR,
    input wire [7:0]                      AP_AXIMM_20_AWLEN,
    input wire [2:0]                      AP_AXIMM_20_AWSIZE,
    input wire [1:0]                      AP_AXIMM_20_AWBURST,
    input wire [1:0]                      AP_AXIMM_20_AWLOCK,
    input wire [3:0]                      AP_AXIMM_20_AWCACHE,
    input wire [2:0]                      AP_AXIMM_20_AWPROT,
    input wire [3:0]                      AP_AXIMM_20_AWREGION,
    input wire [3:0]                      AP_AXIMM_20_AWQOS,
    input wire                            AP_AXIMM_20_AWVALID,
    output  wire                            AP_AXIMM_20_AWREADY,
    input wire [M_AXIMM_20_DATA_WIDTH-1:0]   AP_AXIMM_20_WDATA,
    input wire [M_AXIMM_20_DATA_WIDTH/8-1:0] AP_AXIMM_20_WSTRB,
    input wire                            AP_AXIMM_20_WLAST,
    input wire                            AP_AXIMM_20_WVALID,
    output  wire                            AP_AXIMM_20_WREADY,
    output  wire [1:0]                      AP_AXIMM_20_BRESP,
    output  wire                            AP_AXIMM_20_BVALID,
    input wire                            AP_AXIMM_20_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_20_ARADDR,
    input wire [7:0]                      AP_AXIMM_20_ARLEN,
    input wire [2:0]                      AP_AXIMM_20_ARSIZE,
    input wire [1:0]                      AP_AXIMM_20_ARBURST,
    input wire [1:0]                      AP_AXIMM_20_ARLOCK,
    input wire [3:0]                      AP_AXIMM_20_ARCACHE,
    input wire [2:0]                      AP_AXIMM_20_ARPROT,
    input wire [3:0]                      AP_AXIMM_20_ARREGION,
    input wire [3:0]                      AP_AXIMM_20_ARQOS,
    input wire                            AP_AXIMM_20_ARVALID,
    output  wire                            AP_AXIMM_20_ARREADY,
    output  wire [M_AXIMM_20_DATA_WIDTH-1:0]   AP_AXIMM_20_RDATA,
    output  wire [1:0]                      AP_AXIMM_20_RRESP,
    output  wire                            AP_AXIMM_20_RLAST,
    output  wire                            AP_AXIMM_20_RVALID,
    input  wire                            AP_AXIMM_20_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_20_AWADDR,
    output wire [7:0]                      M_AXIMM_20_AWLEN,
    output wire [2:0]                      M_AXIMM_20_AWSIZE,
    output wire [1:0]                      M_AXIMM_20_AWBURST,
    output wire [1:0]                      M_AXIMM_20_AWLOCK,
    output wire [3:0]                      M_AXIMM_20_AWCACHE,
    output wire [2:0]                      M_AXIMM_20_AWPROT,
    output wire [3:0]                      M_AXIMM_20_AWREGION,
    output wire [3:0]                      M_AXIMM_20_AWQOS,
    output wire                            M_AXIMM_20_AWVALID,
    input  wire                            M_AXIMM_20_AWREADY,
    output wire [M_AXIMM_20_DATA_WIDTH-1:0]   M_AXIMM_20_WDATA,
    output wire [M_AXIMM_20_DATA_WIDTH/8-1:0] M_AXIMM_20_WSTRB,
    output wire                            M_AXIMM_20_WLAST,
    output wire                            M_AXIMM_20_WVALID,
    input  wire                            M_AXIMM_20_WREADY,
    input  wire [1:0]                      M_AXIMM_20_BRESP,
    input  wire                            M_AXIMM_20_BVALID,
    output wire                            M_AXIMM_20_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_20_ARADDR,
    output wire [7:0]                      M_AXIMM_20_ARLEN,
    output wire [2:0]                      M_AXIMM_20_ARSIZE,
    output wire [1:0]                      M_AXIMM_20_ARBURST,
    output wire [1:0]                      M_AXIMM_20_ARLOCK,
    output wire [3:0]                      M_AXIMM_20_ARCACHE,
    output wire [2:0]                      M_AXIMM_20_ARPROT,
    output wire [3:0]                      M_AXIMM_20_ARREGION,
    output wire [3:0]                      M_AXIMM_20_ARQOS,
    output wire                            M_AXIMM_20_ARVALID,
    input  wire                            M_AXIMM_20_ARREADY,
    input  wire [M_AXIMM_20_DATA_WIDTH-1:0]   M_AXIMM_20_RDATA,
    input  wire [1:0]                      M_AXIMM_20_RRESP,
    input  wire                            M_AXIMM_20_RLAST,
    input  wire                            M_AXIMM_20_RVALID,
    output wire                            M_AXIMM_20_RREADY,
    //AXI-MM pass-through interface 21
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_21_AWADDR,
    input wire [7:0]                      AP_AXIMM_21_AWLEN,
    input wire [2:0]                      AP_AXIMM_21_AWSIZE,
    input wire [1:0]                      AP_AXIMM_21_AWBURST,
    input wire [1:0]                      AP_AXIMM_21_AWLOCK,
    input wire [3:0]                      AP_AXIMM_21_AWCACHE,
    input wire [2:0]                      AP_AXIMM_21_AWPROT,
    input wire [3:0]                      AP_AXIMM_21_AWREGION,
    input wire [3:0]                      AP_AXIMM_21_AWQOS,
    input wire                            AP_AXIMM_21_AWVALID,
    output  wire                            AP_AXIMM_21_AWREADY,
    input wire [M_AXIMM_21_DATA_WIDTH-1:0]   AP_AXIMM_21_WDATA,
    input wire [M_AXIMM_21_DATA_WIDTH/8-1:0] AP_AXIMM_21_WSTRB,
    input wire                            AP_AXIMM_21_WLAST,
    input wire                            AP_AXIMM_21_WVALID,
    output  wire                            AP_AXIMM_21_WREADY,
    output  wire [1:0]                      AP_AXIMM_21_BRESP,
    output  wire                            AP_AXIMM_21_BVALID,
    input wire                            AP_AXIMM_21_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_21_ARADDR,
    input wire [7:0]                      AP_AXIMM_21_ARLEN,
    input wire [2:0]                      AP_AXIMM_21_ARSIZE,
    input wire [1:0]                      AP_AXIMM_21_ARBURST,
    input wire [1:0]                      AP_AXIMM_21_ARLOCK,
    input wire [3:0]                      AP_AXIMM_21_ARCACHE,
    input wire [2:0]                      AP_AXIMM_21_ARPROT,
    input wire [3:0]                      AP_AXIMM_21_ARREGION,
    input wire [3:0]                      AP_AXIMM_21_ARQOS,
    input wire                            AP_AXIMM_21_ARVALID,
    output  wire                            AP_AXIMM_21_ARREADY,
    output  wire [M_AXIMM_21_DATA_WIDTH-1:0]   AP_AXIMM_21_RDATA,
    output  wire [1:0]                      AP_AXIMM_21_RRESP,
    output  wire                            AP_AXIMM_21_RLAST,
    output  wire                            AP_AXIMM_21_RVALID,
    input  wire                            AP_AXIMM_21_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_21_AWADDR,
    output wire [7:0]                      M_AXIMM_21_AWLEN,
    output wire [2:0]                      M_AXIMM_21_AWSIZE,
    output wire [1:0]                      M_AXIMM_21_AWBURST,
    output wire [1:0]                      M_AXIMM_21_AWLOCK,
    output wire [3:0]                      M_AXIMM_21_AWCACHE,
    output wire [2:0]                      M_AXIMM_21_AWPROT,
    output wire [3:0]                      M_AXIMM_21_AWREGION,
    output wire [3:0]                      M_AXIMM_21_AWQOS,
    output wire                            M_AXIMM_21_AWVALID,
    input  wire                            M_AXIMM_21_AWREADY,
    output wire [M_AXIMM_21_DATA_WIDTH-1:0]   M_AXIMM_21_WDATA,
    output wire [M_AXIMM_21_DATA_WIDTH/8-1:0] M_AXIMM_21_WSTRB,
    output wire                            M_AXIMM_21_WLAST,
    output wire                            M_AXIMM_21_WVALID,
    input  wire                            M_AXIMM_21_WREADY,
    input  wire [1:0]                      M_AXIMM_21_BRESP,
    input  wire                            M_AXIMM_21_BVALID,
    output wire                            M_AXIMM_21_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_21_ARADDR,
    output wire [7:0]                      M_AXIMM_21_ARLEN,
    output wire [2:0]                      M_AXIMM_21_ARSIZE,
    output wire [1:0]                      M_AXIMM_21_ARBURST,
    output wire [1:0]                      M_AXIMM_21_ARLOCK,
    output wire [3:0]                      M_AXIMM_21_ARCACHE,
    output wire [2:0]                      M_AXIMM_21_ARPROT,
    output wire [3:0]                      M_AXIMM_21_ARREGION,
    output wire [3:0]                      M_AXIMM_21_ARQOS,
    output wire                            M_AXIMM_21_ARVALID,
    input  wire                            M_AXIMM_21_ARREADY,
    input  wire [M_AXIMM_21_DATA_WIDTH-1:0]   M_AXIMM_21_RDATA,
    input  wire [1:0]                      M_AXIMM_21_RRESP,
    input  wire                            M_AXIMM_21_RLAST,
    input  wire                            M_AXIMM_21_RVALID,
    output wire                            M_AXIMM_21_RREADY,
    //AXI-MM pass-through interface 22
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_22_AWADDR,
    input wire [7:0]                      AP_AXIMM_22_AWLEN,
    input wire [2:0]                      AP_AXIMM_22_AWSIZE,
    input wire [1:0]                      AP_AXIMM_22_AWBURST,
    input wire [1:0]                      AP_AXIMM_22_AWLOCK,
    input wire [3:0]                      AP_AXIMM_22_AWCACHE,
    input wire [2:0]                      AP_AXIMM_22_AWPROT,
    input wire [3:0]                      AP_AXIMM_22_AWREGION,
    input wire [3:0]                      AP_AXIMM_22_AWQOS,
    input wire                            AP_AXIMM_22_AWVALID,
    output  wire                            AP_AXIMM_22_AWREADY,
    input wire [M_AXIMM_22_DATA_WIDTH-1:0]   AP_AXIMM_22_WDATA,
    input wire [M_AXIMM_22_DATA_WIDTH/8-1:0] AP_AXIMM_22_WSTRB,
    input wire                            AP_AXIMM_22_WLAST,
    input wire                            AP_AXIMM_22_WVALID,
    output  wire                            AP_AXIMM_22_WREADY,
    output  wire [1:0]                      AP_AXIMM_22_BRESP,
    output  wire                            AP_AXIMM_22_BVALID,
    input wire                            AP_AXIMM_22_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_22_ARADDR,
    input wire [7:0]                      AP_AXIMM_22_ARLEN,
    input wire [2:0]                      AP_AXIMM_22_ARSIZE,
    input wire [1:0]                      AP_AXIMM_22_ARBURST,
    input wire [1:0]                      AP_AXIMM_22_ARLOCK,
    input wire [3:0]                      AP_AXIMM_22_ARCACHE,
    input wire [2:0]                      AP_AXIMM_22_ARPROT,
    input wire [3:0]                      AP_AXIMM_22_ARREGION,
    input wire [3:0]                      AP_AXIMM_22_ARQOS,
    input wire                            AP_AXIMM_22_ARVALID,
    output  wire                            AP_AXIMM_22_ARREADY,
    output  wire [M_AXIMM_22_DATA_WIDTH-1:0]   AP_AXIMM_22_RDATA,
    output  wire [1:0]                      AP_AXIMM_22_RRESP,
    output  wire                            AP_AXIMM_22_RLAST,
    output  wire                            AP_AXIMM_22_RVALID,
    input  wire                            AP_AXIMM_22_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_22_AWADDR,
    output wire [7:0]                      M_AXIMM_22_AWLEN,
    output wire [2:0]                      M_AXIMM_22_AWSIZE,
    output wire [1:0]                      M_AXIMM_22_AWBURST,
    output wire [1:0]                      M_AXIMM_22_AWLOCK,
    output wire [3:0]                      M_AXIMM_22_AWCACHE,
    output wire [2:0]                      M_AXIMM_22_AWPROT,
    output wire [3:0]                      M_AXIMM_22_AWREGION,
    output wire [3:0]                      M_AXIMM_22_AWQOS,
    output wire                            M_AXIMM_22_AWVALID,
    input  wire                            M_AXIMM_22_AWREADY,
    output wire [M_AXIMM_22_DATA_WIDTH-1:0]   M_AXIMM_22_WDATA,
    output wire [M_AXIMM_22_DATA_WIDTH/8-1:0] M_AXIMM_22_WSTRB,
    output wire                            M_AXIMM_22_WLAST,
    output wire                            M_AXIMM_22_WVALID,
    input  wire                            M_AXIMM_22_WREADY,
    input  wire [1:0]                      M_AXIMM_22_BRESP,
    input  wire                            M_AXIMM_22_BVALID,
    output wire                            M_AXIMM_22_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_22_ARADDR,
    output wire [7:0]                      M_AXIMM_22_ARLEN,
    output wire [2:0]                      M_AXIMM_22_ARSIZE,
    output wire [1:0]                      M_AXIMM_22_ARBURST,
    output wire [1:0]                      M_AXIMM_22_ARLOCK,
    output wire [3:0]                      M_AXIMM_22_ARCACHE,
    output wire [2:0]                      M_AXIMM_22_ARPROT,
    output wire [3:0]                      M_AXIMM_22_ARREGION,
    output wire [3:0]                      M_AXIMM_22_ARQOS,
    output wire                            M_AXIMM_22_ARVALID,
    input  wire                            M_AXIMM_22_ARREADY,
    input  wire [M_AXIMM_22_DATA_WIDTH-1:0]   M_AXIMM_22_RDATA,
    input  wire [1:0]                      M_AXIMM_22_RRESP,
    input  wire                            M_AXIMM_22_RLAST,
    input  wire                            M_AXIMM_22_RVALID,
    output wire                            M_AXIMM_22_RREADY,
    //AXI-MM pass-through interface 23
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_23_AWADDR,
    input wire [7:0]                      AP_AXIMM_23_AWLEN,
    input wire [2:0]                      AP_AXIMM_23_AWSIZE,
    input wire [1:0]                      AP_AXIMM_23_AWBURST,
    input wire [1:0]                      AP_AXIMM_23_AWLOCK,
    input wire [3:0]                      AP_AXIMM_23_AWCACHE,
    input wire [2:0]                      AP_AXIMM_23_AWPROT,
    input wire [3:0]                      AP_AXIMM_23_AWREGION,
    input wire [3:0]                      AP_AXIMM_23_AWQOS,
    input wire                            AP_AXIMM_23_AWVALID,
    output  wire                            AP_AXIMM_23_AWREADY,
    input wire [M_AXIMM_23_DATA_WIDTH-1:0]   AP_AXIMM_23_WDATA,
    input wire [M_AXIMM_23_DATA_WIDTH/8-1:0] AP_AXIMM_23_WSTRB,
    input wire                            AP_AXIMM_23_WLAST,
    input wire                            AP_AXIMM_23_WVALID,
    output  wire                            AP_AXIMM_23_WREADY,
    output  wire [1:0]                      AP_AXIMM_23_BRESP,
    output  wire                            AP_AXIMM_23_BVALID,
    input wire                            AP_AXIMM_23_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_23_ARADDR,
    input wire [7:0]                      AP_AXIMM_23_ARLEN,
    input wire [2:0]                      AP_AXIMM_23_ARSIZE,
    input wire [1:0]                      AP_AXIMM_23_ARBURST,
    input wire [1:0]                      AP_AXIMM_23_ARLOCK,
    input wire [3:0]                      AP_AXIMM_23_ARCACHE,
    input wire [2:0]                      AP_AXIMM_23_ARPROT,
    input wire [3:0]                      AP_AXIMM_23_ARREGION,
    input wire [3:0]                      AP_AXIMM_23_ARQOS,
    input wire                            AP_AXIMM_23_ARVALID,
    output  wire                            AP_AXIMM_23_ARREADY,
    output  wire [M_AXIMM_23_DATA_WIDTH-1:0]   AP_AXIMM_23_RDATA,
    output  wire [1:0]                      AP_AXIMM_23_RRESP,
    output  wire                            AP_AXIMM_23_RLAST,
    output  wire                            AP_AXIMM_23_RVALID,
    input  wire                            AP_AXIMM_23_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_23_AWADDR,
    output wire [7:0]                      M_AXIMM_23_AWLEN,
    output wire [2:0]                      M_AXIMM_23_AWSIZE,
    output wire [1:0]                      M_AXIMM_23_AWBURST,
    output wire [1:0]                      M_AXIMM_23_AWLOCK,
    output wire [3:0]                      M_AXIMM_23_AWCACHE,
    output wire [2:0]                      M_AXIMM_23_AWPROT,
    output wire [3:0]                      M_AXIMM_23_AWREGION,
    output wire [3:0]                      M_AXIMM_23_AWQOS,
    output wire                            M_AXIMM_23_AWVALID,
    input  wire                            M_AXIMM_23_AWREADY,
    output wire [M_AXIMM_23_DATA_WIDTH-1:0]   M_AXIMM_23_WDATA,
    output wire [M_AXIMM_23_DATA_WIDTH/8-1:0] M_AXIMM_23_WSTRB,
    output wire                            M_AXIMM_23_WLAST,
    output wire                            M_AXIMM_23_WVALID,
    input  wire                            M_AXIMM_23_WREADY,
    input  wire [1:0]                      M_AXIMM_23_BRESP,
    input  wire                            M_AXIMM_23_BVALID,
    output wire                            M_AXIMM_23_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_23_ARADDR,
    output wire [7:0]                      M_AXIMM_23_ARLEN,
    output wire [2:0]                      M_AXIMM_23_ARSIZE,
    output wire [1:0]                      M_AXIMM_23_ARBURST,
    output wire [1:0]                      M_AXIMM_23_ARLOCK,
    output wire [3:0]                      M_AXIMM_23_ARCACHE,
    output wire [2:0]                      M_AXIMM_23_ARPROT,
    output wire [3:0]                      M_AXIMM_23_ARREGION,
    output wire [3:0]                      M_AXIMM_23_ARQOS,
    output wire                            M_AXIMM_23_ARVALID,
    input  wire                            M_AXIMM_23_ARREADY,
    input  wire [M_AXIMM_23_DATA_WIDTH-1:0]   M_AXIMM_23_RDATA,
    input  wire [1:0]                      M_AXIMM_23_RRESP,
    input  wire                            M_AXIMM_23_RLAST,
    input  wire                            M_AXIMM_23_RVALID,
    output wire                            M_AXIMM_23_RREADY,
    //AXI-MM pass-through interface 24
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_24_AWADDR,
    input wire [7:0]                      AP_AXIMM_24_AWLEN,
    input wire [2:0]                      AP_AXIMM_24_AWSIZE,
    input wire [1:0]                      AP_AXIMM_24_AWBURST,
    input wire [1:0]                      AP_AXIMM_24_AWLOCK,
    input wire [3:0]                      AP_AXIMM_24_AWCACHE,
    input wire [2:0]                      AP_AXIMM_24_AWPROT,
    input wire [3:0]                      AP_AXIMM_24_AWREGION,
    input wire [3:0]                      AP_AXIMM_24_AWQOS,
    input wire                            AP_AXIMM_24_AWVALID,
    output  wire                            AP_AXIMM_24_AWREADY,
    input wire [M_AXIMM_24_DATA_WIDTH-1:0]   AP_AXIMM_24_WDATA,
    input wire [M_AXIMM_24_DATA_WIDTH/8-1:0] AP_AXIMM_24_WSTRB,
    input wire                            AP_AXIMM_24_WLAST,
    input wire                            AP_AXIMM_24_WVALID,
    output  wire                            AP_AXIMM_24_WREADY,
    output  wire [1:0]                      AP_AXIMM_24_BRESP,
    output  wire                            AP_AXIMM_24_BVALID,
    input wire                            AP_AXIMM_24_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_24_ARADDR,
    input wire [7:0]                      AP_AXIMM_24_ARLEN,
    input wire [2:0]                      AP_AXIMM_24_ARSIZE,
    input wire [1:0]                      AP_AXIMM_24_ARBURST,
    input wire [1:0]                      AP_AXIMM_24_ARLOCK,
    input wire [3:0]                      AP_AXIMM_24_ARCACHE,
    input wire [2:0]                      AP_AXIMM_24_ARPROT,
    input wire [3:0]                      AP_AXIMM_24_ARREGION,
    input wire [3:0]                      AP_AXIMM_24_ARQOS,
    input wire                            AP_AXIMM_24_ARVALID,
    output  wire                            AP_AXIMM_24_ARREADY,
    output  wire [M_AXIMM_24_DATA_WIDTH-1:0]   AP_AXIMM_24_RDATA,
    output  wire [1:0]                      AP_AXIMM_24_RRESP,
    output  wire                            AP_AXIMM_24_RLAST,
    output  wire                            AP_AXIMM_24_RVALID,
    input  wire                            AP_AXIMM_24_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_24_AWADDR,
    output wire [7:0]                      M_AXIMM_24_AWLEN,
    output wire [2:0]                      M_AXIMM_24_AWSIZE,
    output wire [1:0]                      M_AXIMM_24_AWBURST,
    output wire [1:0]                      M_AXIMM_24_AWLOCK,
    output wire [3:0]                      M_AXIMM_24_AWCACHE,
    output wire [2:0]                      M_AXIMM_24_AWPROT,
    output wire [3:0]                      M_AXIMM_24_AWREGION,
    output wire [3:0]                      M_AXIMM_24_AWQOS,
    output wire                            M_AXIMM_24_AWVALID,
    input  wire                            M_AXIMM_24_AWREADY,
    output wire [M_AXIMM_24_DATA_WIDTH-1:0]   M_AXIMM_24_WDATA,
    output wire [M_AXIMM_24_DATA_WIDTH/8-1:0] M_AXIMM_24_WSTRB,
    output wire                            M_AXIMM_24_WLAST,
    output wire                            M_AXIMM_24_WVALID,
    input  wire                            M_AXIMM_24_WREADY,
    input  wire [1:0]                      M_AXIMM_24_BRESP,
    input  wire                            M_AXIMM_24_BVALID,
    output wire                            M_AXIMM_24_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_24_ARADDR,
    output wire [7:0]                      M_AXIMM_24_ARLEN,
    output wire [2:0]                      M_AXIMM_24_ARSIZE,
    output wire [1:0]                      M_AXIMM_24_ARBURST,
    output wire [1:0]                      M_AXIMM_24_ARLOCK,
    output wire [3:0]                      M_AXIMM_24_ARCACHE,
    output wire [2:0]                      M_AXIMM_24_ARPROT,
    output wire [3:0]                      M_AXIMM_24_ARREGION,
    output wire [3:0]                      M_AXIMM_24_ARQOS,
    output wire                            M_AXIMM_24_ARVALID,
    input  wire                            M_AXIMM_24_ARREADY,
    input  wire [M_AXIMM_24_DATA_WIDTH-1:0]   M_AXIMM_24_RDATA,
    input  wire [1:0]                      M_AXIMM_24_RRESP,
    input  wire                            M_AXIMM_24_RLAST,
    input  wire                            M_AXIMM_24_RVALID,
    output wire                            M_AXIMM_24_RREADY,
    //AXI-MM pass-through interface 25
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_25_AWADDR,
    input wire [7:0]                      AP_AXIMM_25_AWLEN,
    input wire [2:0]                      AP_AXIMM_25_AWSIZE,
    input wire [1:0]                      AP_AXIMM_25_AWBURST,
    input wire [1:0]                      AP_AXIMM_25_AWLOCK,
    input wire [3:0]                      AP_AXIMM_25_AWCACHE,
    input wire [2:0]                      AP_AXIMM_25_AWPROT,
    input wire [3:0]                      AP_AXIMM_25_AWREGION,
    input wire [3:0]                      AP_AXIMM_25_AWQOS,
    input wire                            AP_AXIMM_25_AWVALID,
    output  wire                            AP_AXIMM_25_AWREADY,
    input wire [M_AXIMM_25_DATA_WIDTH-1:0]   AP_AXIMM_25_WDATA,
    input wire [M_AXIMM_25_DATA_WIDTH/8-1:0] AP_AXIMM_25_WSTRB,
    input wire                            AP_AXIMM_25_WLAST,
    input wire                            AP_AXIMM_25_WVALID,
    output  wire                            AP_AXIMM_25_WREADY,
    output  wire [1:0]                      AP_AXIMM_25_BRESP,
    output  wire                            AP_AXIMM_25_BVALID,
    input wire                            AP_AXIMM_25_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_25_ARADDR,
    input wire [7:0]                      AP_AXIMM_25_ARLEN,
    input wire [2:0]                      AP_AXIMM_25_ARSIZE,
    input wire [1:0]                      AP_AXIMM_25_ARBURST,
    input wire [1:0]                      AP_AXIMM_25_ARLOCK,
    input wire [3:0]                      AP_AXIMM_25_ARCACHE,
    input wire [2:0]                      AP_AXIMM_25_ARPROT,
    input wire [3:0]                      AP_AXIMM_25_ARREGION,
    input wire [3:0]                      AP_AXIMM_25_ARQOS,
    input wire                            AP_AXIMM_25_ARVALID,
    output  wire                            AP_AXIMM_25_ARREADY,
    output  wire [M_AXIMM_25_DATA_WIDTH-1:0]   AP_AXIMM_25_RDATA,
    output  wire [1:0]                      AP_AXIMM_25_RRESP,
    output  wire                            AP_AXIMM_25_RLAST,
    output  wire                            AP_AXIMM_25_RVALID,
    input  wire                            AP_AXIMM_25_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_25_AWADDR,
    output wire [7:0]                      M_AXIMM_25_AWLEN,
    output wire [2:0]                      M_AXIMM_25_AWSIZE,
    output wire [1:0]                      M_AXIMM_25_AWBURST,
    output wire [1:0]                      M_AXIMM_25_AWLOCK,
    output wire [3:0]                      M_AXIMM_25_AWCACHE,
    output wire [2:0]                      M_AXIMM_25_AWPROT,
    output wire [3:0]                      M_AXIMM_25_AWREGION,
    output wire [3:0]                      M_AXIMM_25_AWQOS,
    output wire                            M_AXIMM_25_AWVALID,
    input  wire                            M_AXIMM_25_AWREADY,
    output wire [M_AXIMM_25_DATA_WIDTH-1:0]   M_AXIMM_25_WDATA,
    output wire [M_AXIMM_25_DATA_WIDTH/8-1:0] M_AXIMM_25_WSTRB,
    output wire                            M_AXIMM_25_WLAST,
    output wire                            M_AXIMM_25_WVALID,
    input  wire                            M_AXIMM_25_WREADY,
    input  wire [1:0]                      M_AXIMM_25_BRESP,
    input  wire                            M_AXIMM_25_BVALID,
    output wire                            M_AXIMM_25_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_25_ARADDR,
    output wire [7:0]                      M_AXIMM_25_ARLEN,
    output wire [2:0]                      M_AXIMM_25_ARSIZE,
    output wire [1:0]                      M_AXIMM_25_ARBURST,
    output wire [1:0]                      M_AXIMM_25_ARLOCK,
    output wire [3:0]                      M_AXIMM_25_ARCACHE,
    output wire [2:0]                      M_AXIMM_25_ARPROT,
    output wire [3:0]                      M_AXIMM_25_ARREGION,
    output wire [3:0]                      M_AXIMM_25_ARQOS,
    output wire                            M_AXIMM_25_ARVALID,
    input  wire                            M_AXIMM_25_ARREADY,
    input  wire [M_AXIMM_25_DATA_WIDTH-1:0]   M_AXIMM_25_RDATA,
    input  wire [1:0]                      M_AXIMM_25_RRESP,
    input  wire                            M_AXIMM_25_RLAST,
    input  wire                            M_AXIMM_25_RVALID,
    output wire                            M_AXIMM_25_RREADY,
    //AXI-MM pass-through interface 26
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_26_AWADDR,
    input wire [7:0]                      AP_AXIMM_26_AWLEN,
    input wire [2:0]                      AP_AXIMM_26_AWSIZE,
    input wire [1:0]                      AP_AXIMM_26_AWBURST,
    input wire [1:0]                      AP_AXIMM_26_AWLOCK,
    input wire [3:0]                      AP_AXIMM_26_AWCACHE,
    input wire [2:0]                      AP_AXIMM_26_AWPROT,
    input wire [3:0]                      AP_AXIMM_26_AWREGION,
    input wire [3:0]                      AP_AXIMM_26_AWQOS,
    input wire                            AP_AXIMM_26_AWVALID,
    output  wire                            AP_AXIMM_26_AWREADY,
    input wire [M_AXIMM_26_DATA_WIDTH-1:0]   AP_AXIMM_26_WDATA,
    input wire [M_AXIMM_26_DATA_WIDTH/8-1:0] AP_AXIMM_26_WSTRB,
    input wire                            AP_AXIMM_26_WLAST,
    input wire                            AP_AXIMM_26_WVALID,
    output  wire                            AP_AXIMM_26_WREADY,
    output  wire [1:0]                      AP_AXIMM_26_BRESP,
    output  wire                            AP_AXIMM_26_BVALID,
    input wire                            AP_AXIMM_26_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_26_ARADDR,
    input wire [7:0]                      AP_AXIMM_26_ARLEN,
    input wire [2:0]                      AP_AXIMM_26_ARSIZE,
    input wire [1:0]                      AP_AXIMM_26_ARBURST,
    input wire [1:0]                      AP_AXIMM_26_ARLOCK,
    input wire [3:0]                      AP_AXIMM_26_ARCACHE,
    input wire [2:0]                      AP_AXIMM_26_ARPROT,
    input wire [3:0]                      AP_AXIMM_26_ARREGION,
    input wire [3:0]                      AP_AXIMM_26_ARQOS,
    input wire                            AP_AXIMM_26_ARVALID,
    output  wire                            AP_AXIMM_26_ARREADY,
    output  wire [M_AXIMM_26_DATA_WIDTH-1:0]   AP_AXIMM_26_RDATA,
    output  wire [1:0]                      AP_AXIMM_26_RRESP,
    output  wire                            AP_AXIMM_26_RLAST,
    output  wire                            AP_AXIMM_26_RVALID,
    input  wire                            AP_AXIMM_26_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_26_AWADDR,
    output wire [7:0]                      M_AXIMM_26_AWLEN,
    output wire [2:0]                      M_AXIMM_26_AWSIZE,
    output wire [1:0]                      M_AXIMM_26_AWBURST,
    output wire [1:0]                      M_AXIMM_26_AWLOCK,
    output wire [3:0]                      M_AXIMM_26_AWCACHE,
    output wire [2:0]                      M_AXIMM_26_AWPROT,
    output wire [3:0]                      M_AXIMM_26_AWREGION,
    output wire [3:0]                      M_AXIMM_26_AWQOS,
    output wire                            M_AXIMM_26_AWVALID,
    input  wire                            M_AXIMM_26_AWREADY,
    output wire [M_AXIMM_26_DATA_WIDTH-1:0]   M_AXIMM_26_WDATA,
    output wire [M_AXIMM_26_DATA_WIDTH/8-1:0] M_AXIMM_26_WSTRB,
    output wire                            M_AXIMM_26_WLAST,
    output wire                            M_AXIMM_26_WVALID,
    input  wire                            M_AXIMM_26_WREADY,
    input  wire [1:0]                      M_AXIMM_26_BRESP,
    input  wire                            M_AXIMM_26_BVALID,
    output wire                            M_AXIMM_26_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_26_ARADDR,
    output wire [7:0]                      M_AXIMM_26_ARLEN,
    output wire [2:0]                      M_AXIMM_26_ARSIZE,
    output wire [1:0]                      M_AXIMM_26_ARBURST,
    output wire [1:0]                      M_AXIMM_26_ARLOCK,
    output wire [3:0]                      M_AXIMM_26_ARCACHE,
    output wire [2:0]                      M_AXIMM_26_ARPROT,
    output wire [3:0]                      M_AXIMM_26_ARREGION,
    output wire [3:0]                      M_AXIMM_26_ARQOS,
    output wire                            M_AXIMM_26_ARVALID,
    input  wire                            M_AXIMM_26_ARREADY,
    input  wire [M_AXIMM_26_DATA_WIDTH-1:0]   M_AXIMM_26_RDATA,
    input  wire [1:0]                      M_AXIMM_26_RRESP,
    input  wire                            M_AXIMM_26_RLAST,
    input  wire                            M_AXIMM_26_RVALID,
    output wire                            M_AXIMM_26_RREADY,
    //AXI-MM pass-through interface 27
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_27_AWADDR,
    input wire [7:0]                      AP_AXIMM_27_AWLEN,
    input wire [2:0]                      AP_AXIMM_27_AWSIZE,
    input wire [1:0]                      AP_AXIMM_27_AWBURST,
    input wire [1:0]                      AP_AXIMM_27_AWLOCK,
    input wire [3:0]                      AP_AXIMM_27_AWCACHE,
    input wire [2:0]                      AP_AXIMM_27_AWPROT,
    input wire [3:0]                      AP_AXIMM_27_AWREGION,
    input wire [3:0]                      AP_AXIMM_27_AWQOS,
    input wire                            AP_AXIMM_27_AWVALID,
    output  wire                            AP_AXIMM_27_AWREADY,
    input wire [M_AXIMM_27_DATA_WIDTH-1:0]   AP_AXIMM_27_WDATA,
    input wire [M_AXIMM_27_DATA_WIDTH/8-1:0] AP_AXIMM_27_WSTRB,
    input wire                            AP_AXIMM_27_WLAST,
    input wire                            AP_AXIMM_27_WVALID,
    output  wire                            AP_AXIMM_27_WREADY,
    output  wire [1:0]                      AP_AXIMM_27_BRESP,
    output  wire                            AP_AXIMM_27_BVALID,
    input wire                            AP_AXIMM_27_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_27_ARADDR,
    input wire [7:0]                      AP_AXIMM_27_ARLEN,
    input wire [2:0]                      AP_AXIMM_27_ARSIZE,
    input wire [1:0]                      AP_AXIMM_27_ARBURST,
    input wire [1:0]                      AP_AXIMM_27_ARLOCK,
    input wire [3:0]                      AP_AXIMM_27_ARCACHE,
    input wire [2:0]                      AP_AXIMM_27_ARPROT,
    input wire [3:0]                      AP_AXIMM_27_ARREGION,
    input wire [3:0]                      AP_AXIMM_27_ARQOS,
    input wire                            AP_AXIMM_27_ARVALID,
    output  wire                            AP_AXIMM_27_ARREADY,
    output  wire [M_AXIMM_27_DATA_WIDTH-1:0]   AP_AXIMM_27_RDATA,
    output  wire [1:0]                      AP_AXIMM_27_RRESP,
    output  wire                            AP_AXIMM_27_RLAST,
    output  wire                            AP_AXIMM_27_RVALID,
    input  wire                            AP_AXIMM_27_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_27_AWADDR,
    output wire [7:0]                      M_AXIMM_27_AWLEN,
    output wire [2:0]                      M_AXIMM_27_AWSIZE,
    output wire [1:0]                      M_AXIMM_27_AWBURST,
    output wire [1:0]                      M_AXIMM_27_AWLOCK,
    output wire [3:0]                      M_AXIMM_27_AWCACHE,
    output wire [2:0]                      M_AXIMM_27_AWPROT,
    output wire [3:0]                      M_AXIMM_27_AWREGION,
    output wire [3:0]                      M_AXIMM_27_AWQOS,
    output wire                            M_AXIMM_27_AWVALID,
    input  wire                            M_AXIMM_27_AWREADY,
    output wire [M_AXIMM_27_DATA_WIDTH-1:0]   M_AXIMM_27_WDATA,
    output wire [M_AXIMM_27_DATA_WIDTH/8-1:0] M_AXIMM_27_WSTRB,
    output wire                            M_AXIMM_27_WLAST,
    output wire                            M_AXIMM_27_WVALID,
    input  wire                            M_AXIMM_27_WREADY,
    input  wire [1:0]                      M_AXIMM_27_BRESP,
    input  wire                            M_AXIMM_27_BVALID,
    output wire                            M_AXIMM_27_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_27_ARADDR,
    output wire [7:0]                      M_AXIMM_27_ARLEN,
    output wire [2:0]                      M_AXIMM_27_ARSIZE,
    output wire [1:0]                      M_AXIMM_27_ARBURST,
    output wire [1:0]                      M_AXIMM_27_ARLOCK,
    output wire [3:0]                      M_AXIMM_27_ARCACHE,
    output wire [2:0]                      M_AXIMM_27_ARPROT,
    output wire [3:0]                      M_AXIMM_27_ARREGION,
    output wire [3:0]                      M_AXIMM_27_ARQOS,
    output wire                            M_AXIMM_27_ARVALID,
    input  wire                            M_AXIMM_27_ARREADY,
    input  wire [M_AXIMM_27_DATA_WIDTH-1:0]   M_AXIMM_27_RDATA,
    input  wire [1:0]                      M_AXIMM_27_RRESP,
    input  wire                            M_AXIMM_27_RLAST,
    input  wire                            M_AXIMM_27_RVALID,
    output wire                            M_AXIMM_27_RREADY,
    //AXI-MM pass-through interface 28
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_28_AWADDR,
    input wire [7:0]                      AP_AXIMM_28_AWLEN,
    input wire [2:0]                      AP_AXIMM_28_AWSIZE,
    input wire [1:0]                      AP_AXIMM_28_AWBURST,
    input wire [1:0]                      AP_AXIMM_28_AWLOCK,
    input wire [3:0]                      AP_AXIMM_28_AWCACHE,
    input wire [2:0]                      AP_AXIMM_28_AWPROT,
    input wire [3:0]                      AP_AXIMM_28_AWREGION,
    input wire [3:0]                      AP_AXIMM_28_AWQOS,
    input wire                            AP_AXIMM_28_AWVALID,
    output  wire                            AP_AXIMM_28_AWREADY,
    input wire [M_AXIMM_28_DATA_WIDTH-1:0]   AP_AXIMM_28_WDATA,
    input wire [M_AXIMM_28_DATA_WIDTH/8-1:0] AP_AXIMM_28_WSTRB,
    input wire                            AP_AXIMM_28_WLAST,
    input wire                            AP_AXIMM_28_WVALID,
    output  wire                            AP_AXIMM_28_WREADY,
    output  wire [1:0]                      AP_AXIMM_28_BRESP,
    output  wire                            AP_AXIMM_28_BVALID,
    input wire                            AP_AXIMM_28_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_28_ARADDR,
    input wire [7:0]                      AP_AXIMM_28_ARLEN,
    input wire [2:0]                      AP_AXIMM_28_ARSIZE,
    input wire [1:0]                      AP_AXIMM_28_ARBURST,
    input wire [1:0]                      AP_AXIMM_28_ARLOCK,
    input wire [3:0]                      AP_AXIMM_28_ARCACHE,
    input wire [2:0]                      AP_AXIMM_28_ARPROT,
    input wire [3:0]                      AP_AXIMM_28_ARREGION,
    input wire [3:0]                      AP_AXIMM_28_ARQOS,
    input wire                            AP_AXIMM_28_ARVALID,
    output  wire                            AP_AXIMM_28_ARREADY,
    output  wire [M_AXIMM_28_DATA_WIDTH-1:0]   AP_AXIMM_28_RDATA,
    output  wire [1:0]                      AP_AXIMM_28_RRESP,
    output  wire                            AP_AXIMM_28_RLAST,
    output  wire                            AP_AXIMM_28_RVALID,
    input  wire                            AP_AXIMM_28_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_28_AWADDR,
    output wire [7:0]                      M_AXIMM_28_AWLEN,
    output wire [2:0]                      M_AXIMM_28_AWSIZE,
    output wire [1:0]                      M_AXIMM_28_AWBURST,
    output wire [1:0]                      M_AXIMM_28_AWLOCK,
    output wire [3:0]                      M_AXIMM_28_AWCACHE,
    output wire [2:0]                      M_AXIMM_28_AWPROT,
    output wire [3:0]                      M_AXIMM_28_AWREGION,
    output wire [3:0]                      M_AXIMM_28_AWQOS,
    output wire                            M_AXIMM_28_AWVALID,
    input  wire                            M_AXIMM_28_AWREADY,
    output wire [M_AXIMM_28_DATA_WIDTH-1:0]   M_AXIMM_28_WDATA,
    output wire [M_AXIMM_28_DATA_WIDTH/8-1:0] M_AXIMM_28_WSTRB,
    output wire                            M_AXIMM_28_WLAST,
    output wire                            M_AXIMM_28_WVALID,
    input  wire                            M_AXIMM_28_WREADY,
    input  wire [1:0]                      M_AXIMM_28_BRESP,
    input  wire                            M_AXIMM_28_BVALID,
    output wire                            M_AXIMM_28_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_28_ARADDR,
    output wire [7:0]                      M_AXIMM_28_ARLEN,
    output wire [2:0]                      M_AXIMM_28_ARSIZE,
    output wire [1:0]                      M_AXIMM_28_ARBURST,
    output wire [1:0]                      M_AXIMM_28_ARLOCK,
    output wire [3:0]                      M_AXIMM_28_ARCACHE,
    output wire [2:0]                      M_AXIMM_28_ARPROT,
    output wire [3:0]                      M_AXIMM_28_ARREGION,
    output wire [3:0]                      M_AXIMM_28_ARQOS,
    output wire                            M_AXIMM_28_ARVALID,
    input  wire                            M_AXIMM_28_ARREADY,
    input  wire [M_AXIMM_28_DATA_WIDTH-1:0]   M_AXIMM_28_RDATA,
    input  wire [1:0]                      M_AXIMM_28_RRESP,
    input  wire                            M_AXIMM_28_RLAST,
    input  wire                            M_AXIMM_28_RVALID,
    output wire                            M_AXIMM_28_RREADY,
    //AXI-MM pass-through interface 29
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_29_AWADDR,
    input wire [7:0]                      AP_AXIMM_29_AWLEN,
    input wire [2:0]                      AP_AXIMM_29_AWSIZE,
    input wire [1:0]                      AP_AXIMM_29_AWBURST,
    input wire [1:0]                      AP_AXIMM_29_AWLOCK,
    input wire [3:0]                      AP_AXIMM_29_AWCACHE,
    input wire [2:0]                      AP_AXIMM_29_AWPROT,
    input wire [3:0]                      AP_AXIMM_29_AWREGION,
    input wire [3:0]                      AP_AXIMM_29_AWQOS,
    input wire                            AP_AXIMM_29_AWVALID,
    output  wire                            AP_AXIMM_29_AWREADY,
    input wire [M_AXIMM_29_DATA_WIDTH-1:0]   AP_AXIMM_29_WDATA,
    input wire [M_AXIMM_29_DATA_WIDTH/8-1:0] AP_AXIMM_29_WSTRB,
    input wire                            AP_AXIMM_29_WLAST,
    input wire                            AP_AXIMM_29_WVALID,
    output  wire                            AP_AXIMM_29_WREADY,
    output  wire [1:0]                      AP_AXIMM_29_BRESP,
    output  wire                            AP_AXIMM_29_BVALID,
    input wire                            AP_AXIMM_29_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_29_ARADDR,
    input wire [7:0]                      AP_AXIMM_29_ARLEN,
    input wire [2:0]                      AP_AXIMM_29_ARSIZE,
    input wire [1:0]                      AP_AXIMM_29_ARBURST,
    input wire [1:0]                      AP_AXIMM_29_ARLOCK,
    input wire [3:0]                      AP_AXIMM_29_ARCACHE,
    input wire [2:0]                      AP_AXIMM_29_ARPROT,
    input wire [3:0]                      AP_AXIMM_29_ARREGION,
    input wire [3:0]                      AP_AXIMM_29_ARQOS,
    input wire                            AP_AXIMM_29_ARVALID,
    output  wire                            AP_AXIMM_29_ARREADY,
    output  wire [M_AXIMM_29_DATA_WIDTH-1:0]   AP_AXIMM_29_RDATA,
    output  wire [1:0]                      AP_AXIMM_29_RRESP,
    output  wire                            AP_AXIMM_29_RLAST,
    output  wire                            AP_AXIMM_29_RVALID,
    input  wire                            AP_AXIMM_29_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_29_AWADDR,
    output wire [7:0]                      M_AXIMM_29_AWLEN,
    output wire [2:0]                      M_AXIMM_29_AWSIZE,
    output wire [1:0]                      M_AXIMM_29_AWBURST,
    output wire [1:0]                      M_AXIMM_29_AWLOCK,
    output wire [3:0]                      M_AXIMM_29_AWCACHE,
    output wire [2:0]                      M_AXIMM_29_AWPROT,
    output wire [3:0]                      M_AXIMM_29_AWREGION,
    output wire [3:0]                      M_AXIMM_29_AWQOS,
    output wire                            M_AXIMM_29_AWVALID,
    input  wire                            M_AXIMM_29_AWREADY,
    output wire [M_AXIMM_29_DATA_WIDTH-1:0]   M_AXIMM_29_WDATA,
    output wire [M_AXIMM_29_DATA_WIDTH/8-1:0] M_AXIMM_29_WSTRB,
    output wire                            M_AXIMM_29_WLAST,
    output wire                            M_AXIMM_29_WVALID,
    input  wire                            M_AXIMM_29_WREADY,
    input  wire [1:0]                      M_AXIMM_29_BRESP,
    input  wire                            M_AXIMM_29_BVALID,
    output wire                            M_AXIMM_29_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_29_ARADDR,
    output wire [7:0]                      M_AXIMM_29_ARLEN,
    output wire [2:0]                      M_AXIMM_29_ARSIZE,
    output wire [1:0]                      M_AXIMM_29_ARBURST,
    output wire [1:0]                      M_AXIMM_29_ARLOCK,
    output wire [3:0]                      M_AXIMM_29_ARCACHE,
    output wire [2:0]                      M_AXIMM_29_ARPROT,
    output wire [3:0]                      M_AXIMM_29_ARREGION,
    output wire [3:0]                      M_AXIMM_29_ARQOS,
    output wire                            M_AXIMM_29_ARVALID,
    input  wire                            M_AXIMM_29_ARREADY,
    input  wire [M_AXIMM_29_DATA_WIDTH-1:0]   M_AXIMM_29_RDATA,
    input  wire [1:0]                      M_AXIMM_29_RRESP,
    input  wire                            M_AXIMM_29_RLAST,
    input  wire                            M_AXIMM_29_RVALID,
    output wire                            M_AXIMM_29_RREADY,
    //AXI-MM pass-through interface 30
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_30_AWADDR,
    input wire [7:0]                      AP_AXIMM_30_AWLEN,
    input wire [2:0]                      AP_AXIMM_30_AWSIZE,
    input wire [1:0]                      AP_AXIMM_30_AWBURST,
    input wire [1:0]                      AP_AXIMM_30_AWLOCK,
    input wire [3:0]                      AP_AXIMM_30_AWCACHE,
    input wire [2:0]                      AP_AXIMM_30_AWPROT,
    input wire [3:0]                      AP_AXIMM_30_AWREGION,
    input wire [3:0]                      AP_AXIMM_30_AWQOS,
    input wire                            AP_AXIMM_30_AWVALID,
    output  wire                            AP_AXIMM_30_AWREADY,
    input wire [M_AXIMM_30_DATA_WIDTH-1:0]   AP_AXIMM_30_WDATA,
    input wire [M_AXIMM_30_DATA_WIDTH/8-1:0] AP_AXIMM_30_WSTRB,
    input wire                            AP_AXIMM_30_WLAST,
    input wire                            AP_AXIMM_30_WVALID,
    output  wire                            AP_AXIMM_30_WREADY,
    output  wire [1:0]                      AP_AXIMM_30_BRESP,
    output  wire                            AP_AXIMM_30_BVALID,
    input wire                            AP_AXIMM_30_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_30_ARADDR,
    input wire [7:0]                      AP_AXIMM_30_ARLEN,
    input wire [2:0]                      AP_AXIMM_30_ARSIZE,
    input wire [1:0]                      AP_AXIMM_30_ARBURST,
    input wire [1:0]                      AP_AXIMM_30_ARLOCK,
    input wire [3:0]                      AP_AXIMM_30_ARCACHE,
    input wire [2:0]                      AP_AXIMM_30_ARPROT,
    input wire [3:0]                      AP_AXIMM_30_ARREGION,
    input wire [3:0]                      AP_AXIMM_30_ARQOS,
    input wire                            AP_AXIMM_30_ARVALID,
    output  wire                            AP_AXIMM_30_ARREADY,
    output  wire [M_AXIMM_30_DATA_WIDTH-1:0]   AP_AXIMM_30_RDATA,
    output  wire [1:0]                      AP_AXIMM_30_RRESP,
    output  wire                            AP_AXIMM_30_RLAST,
    output  wire                            AP_AXIMM_30_RVALID,
    input  wire                            AP_AXIMM_30_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_30_AWADDR,
    output wire [7:0]                      M_AXIMM_30_AWLEN,
    output wire [2:0]                      M_AXIMM_30_AWSIZE,
    output wire [1:0]                      M_AXIMM_30_AWBURST,
    output wire [1:0]                      M_AXIMM_30_AWLOCK,
    output wire [3:0]                      M_AXIMM_30_AWCACHE,
    output wire [2:0]                      M_AXIMM_30_AWPROT,
    output wire [3:0]                      M_AXIMM_30_AWREGION,
    output wire [3:0]                      M_AXIMM_30_AWQOS,
    output wire                            M_AXIMM_30_AWVALID,
    input  wire                            M_AXIMM_30_AWREADY,
    output wire [M_AXIMM_30_DATA_WIDTH-1:0]   M_AXIMM_30_WDATA,
    output wire [M_AXIMM_30_DATA_WIDTH/8-1:0] M_AXIMM_30_WSTRB,
    output wire                            M_AXIMM_30_WLAST,
    output wire                            M_AXIMM_30_WVALID,
    input  wire                            M_AXIMM_30_WREADY,
    input  wire [1:0]                      M_AXIMM_30_BRESP,
    input  wire                            M_AXIMM_30_BVALID,
    output wire                            M_AXIMM_30_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_30_ARADDR,
    output wire [7:0]                      M_AXIMM_30_ARLEN,
    output wire [2:0]                      M_AXIMM_30_ARSIZE,
    output wire [1:0]                      M_AXIMM_30_ARBURST,
    output wire [1:0]                      M_AXIMM_30_ARLOCK,
    output wire [3:0]                      M_AXIMM_30_ARCACHE,
    output wire [2:0]                      M_AXIMM_30_ARPROT,
    output wire [3:0]                      M_AXIMM_30_ARREGION,
    output wire [3:0]                      M_AXIMM_30_ARQOS,
    output wire                            M_AXIMM_30_ARVALID,
    input  wire                            M_AXIMM_30_ARREADY,
    input  wire [M_AXIMM_30_DATA_WIDTH-1:0]   M_AXIMM_30_RDATA,
    input  wire [1:0]                      M_AXIMM_30_RRESP,
    input  wire                            M_AXIMM_30_RLAST,
    input  wire                            M_AXIMM_30_RVALID,
    output wire                            M_AXIMM_30_RREADY,
    //AXI-MM pass-through interface 31
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_31_AWADDR,
    input wire [7:0]                      AP_AXIMM_31_AWLEN,
    input wire [2:0]                      AP_AXIMM_31_AWSIZE,
    input wire [1:0]                      AP_AXIMM_31_AWBURST,
    input wire [1:0]                      AP_AXIMM_31_AWLOCK,
    input wire [3:0]                      AP_AXIMM_31_AWCACHE,
    input wire [2:0]                      AP_AXIMM_31_AWPROT,
    input wire [3:0]                      AP_AXIMM_31_AWREGION,
    input wire [3:0]                      AP_AXIMM_31_AWQOS,
    input wire                            AP_AXIMM_31_AWVALID,
    output  wire                            AP_AXIMM_31_AWREADY,
    input wire [M_AXIMM_31_DATA_WIDTH-1:0]   AP_AXIMM_31_WDATA,
    input wire [M_AXIMM_31_DATA_WIDTH/8-1:0] AP_AXIMM_31_WSTRB,
    input wire                            AP_AXIMM_31_WLAST,
    input wire                            AP_AXIMM_31_WVALID,
    output  wire                            AP_AXIMM_31_WREADY,
    output  wire [1:0]                      AP_AXIMM_31_BRESP,
    output  wire                            AP_AXIMM_31_BVALID,
    input wire                            AP_AXIMM_31_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_31_ARADDR,
    input wire [7:0]                      AP_AXIMM_31_ARLEN,
    input wire [2:0]                      AP_AXIMM_31_ARSIZE,
    input wire [1:0]                      AP_AXIMM_31_ARBURST,
    input wire [1:0]                      AP_AXIMM_31_ARLOCK,
    input wire [3:0]                      AP_AXIMM_31_ARCACHE,
    input wire [2:0]                      AP_AXIMM_31_ARPROT,
    input wire [3:0]                      AP_AXIMM_31_ARREGION,
    input wire [3:0]                      AP_AXIMM_31_ARQOS,
    input wire                            AP_AXIMM_31_ARVALID,
    output  wire                            AP_AXIMM_31_ARREADY,
    output  wire [M_AXIMM_31_DATA_WIDTH-1:0]   AP_AXIMM_31_RDATA,
    output  wire [1:0]                      AP_AXIMM_31_RRESP,
    output  wire                            AP_AXIMM_31_RLAST,
    output  wire                            AP_AXIMM_31_RVALID,
    input  wire                            AP_AXIMM_31_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_31_AWADDR,
    output wire [7:0]                      M_AXIMM_31_AWLEN,
    output wire [2:0]                      M_AXIMM_31_AWSIZE,
    output wire [1:0]                      M_AXIMM_31_AWBURST,
    output wire [1:0]                      M_AXIMM_31_AWLOCK,
    output wire [3:0]                      M_AXIMM_31_AWCACHE,
    output wire [2:0]                      M_AXIMM_31_AWPROT,
    output wire [3:0]                      M_AXIMM_31_AWREGION,
    output wire [3:0]                      M_AXIMM_31_AWQOS,
    output wire                            M_AXIMM_31_AWVALID,
    input  wire                            M_AXIMM_31_AWREADY,
    output wire [M_AXIMM_31_DATA_WIDTH-1:0]   M_AXIMM_31_WDATA,
    output wire [M_AXIMM_31_DATA_WIDTH/8-1:0] M_AXIMM_31_WSTRB,
    output wire                            M_AXIMM_31_WLAST,
    output wire                            M_AXIMM_31_WVALID,
    input  wire                            M_AXIMM_31_WREADY,
    input  wire [1:0]                      M_AXIMM_31_BRESP,
    input  wire                            M_AXIMM_31_BVALID,
    output wire                            M_AXIMM_31_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_31_ARADDR,
    output wire [7:0]                      M_AXIMM_31_ARLEN,
    output wire [2:0]                      M_AXIMM_31_ARSIZE,
    output wire [1:0]                      M_AXIMM_31_ARBURST,
    output wire [1:0]                      M_AXIMM_31_ARLOCK,
    output wire [3:0]                      M_AXIMM_31_ARCACHE,
    output wire [2:0]                      M_AXIMM_31_ARPROT,
    output wire [3:0]                      M_AXIMM_31_ARREGION,
    output wire [3:0]                      M_AXIMM_31_ARQOS,
    output wire                            M_AXIMM_31_ARVALID,
    input  wire                            M_AXIMM_31_ARREADY,
    input  wire [M_AXIMM_31_DATA_WIDTH-1:0]   M_AXIMM_31_RDATA,
    input  wire [1:0]                      M_AXIMM_31_RRESP,
    input  wire                            M_AXIMM_31_RLAST,
    input  wire                            M_AXIMM_31_RVALID,
    output wire                            M_AXIMM_31_RREADY,
    //AXI-MM pass-through interface 32
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_32_AWADDR,
    input wire [7:0]                      AP_AXIMM_32_AWLEN,
    input wire [2:0]                      AP_AXIMM_32_AWSIZE,
    input wire [1:0]                      AP_AXIMM_32_AWBURST,
    input wire [1:0]                      AP_AXIMM_32_AWLOCK,
    input wire [3:0]                      AP_AXIMM_32_AWCACHE,
    input wire [2:0]                      AP_AXIMM_32_AWPROT,
    input wire [3:0]                      AP_AXIMM_32_AWREGION,
    input wire [3:0]                      AP_AXIMM_32_AWQOS,
    input wire                            AP_AXIMM_32_AWVALID,
    output  wire                            AP_AXIMM_32_AWREADY,
    input wire [M_AXIMM_32_DATA_WIDTH-1:0]   AP_AXIMM_32_WDATA,
    input wire [M_AXIMM_32_DATA_WIDTH/8-1:0] AP_AXIMM_32_WSTRB,
    input wire                            AP_AXIMM_32_WLAST,
    input wire                            AP_AXIMM_32_WVALID,
    output  wire                            AP_AXIMM_32_WREADY,
    output  wire [1:0]                      AP_AXIMM_32_BRESP,
    output  wire                            AP_AXIMM_32_BVALID,
    input wire                            AP_AXIMM_32_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_32_ARADDR,
    input wire [7:0]                      AP_AXIMM_32_ARLEN,
    input wire [2:0]                      AP_AXIMM_32_ARSIZE,
    input wire [1:0]                      AP_AXIMM_32_ARBURST,
    input wire [1:0]                      AP_AXIMM_32_ARLOCK,
    input wire [3:0]                      AP_AXIMM_32_ARCACHE,
    input wire [2:0]                      AP_AXIMM_32_ARPROT,
    input wire [3:0]                      AP_AXIMM_32_ARREGION,
    input wire [3:0]                      AP_AXIMM_32_ARQOS,
    input wire                            AP_AXIMM_32_ARVALID,
    output  wire                            AP_AXIMM_32_ARREADY,
    output  wire [M_AXIMM_32_DATA_WIDTH-1:0]   AP_AXIMM_32_RDATA,
    output  wire [1:0]                      AP_AXIMM_32_RRESP,
    output  wire                            AP_AXIMM_32_RLAST,
    output  wire                            AP_AXIMM_32_RVALID,
    input  wire                            AP_AXIMM_32_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_32_AWADDR,
    output wire [7:0]                      M_AXIMM_32_AWLEN,
    output wire [2:0]                      M_AXIMM_32_AWSIZE,
    output wire [1:0]                      M_AXIMM_32_AWBURST,
    output wire [1:0]                      M_AXIMM_32_AWLOCK,
    output wire [3:0]                      M_AXIMM_32_AWCACHE,
    output wire [2:0]                      M_AXIMM_32_AWPROT,
    output wire [3:0]                      M_AXIMM_32_AWREGION,
    output wire [3:0]                      M_AXIMM_32_AWQOS,
    output wire                            M_AXIMM_32_AWVALID,
    input  wire                            M_AXIMM_32_AWREADY,
    output wire [M_AXIMM_32_DATA_WIDTH-1:0]   M_AXIMM_32_WDATA,
    output wire [M_AXIMM_32_DATA_WIDTH/8-1:0] M_AXIMM_32_WSTRB,
    output wire                            M_AXIMM_32_WLAST,
    output wire                            M_AXIMM_32_WVALID,
    input  wire                            M_AXIMM_32_WREADY,
    input  wire [1:0]                      M_AXIMM_32_BRESP,
    input  wire                            M_AXIMM_32_BVALID,
    output wire                            M_AXIMM_32_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_32_ARADDR,
    output wire [7:0]                      M_AXIMM_32_ARLEN,
    output wire [2:0]                      M_AXIMM_32_ARSIZE,
    output wire [1:0]                      M_AXIMM_32_ARBURST,
    output wire [1:0]                      M_AXIMM_32_ARLOCK,
    output wire [3:0]                      M_AXIMM_32_ARCACHE,
    output wire [2:0]                      M_AXIMM_32_ARPROT,
    output wire [3:0]                      M_AXIMM_32_ARREGION,
    output wire [3:0]                      M_AXIMM_32_ARQOS,
    output wire                            M_AXIMM_32_ARVALID,
    input  wire                            M_AXIMM_32_ARREADY,
    input  wire [M_AXIMM_32_DATA_WIDTH-1:0]   M_AXIMM_32_RDATA,
    input  wire [1:0]                      M_AXIMM_32_RRESP,
    input  wire                            M_AXIMM_32_RLAST,
    input  wire                            M_AXIMM_32_RVALID,
    output wire                            M_AXIMM_32_RREADY,
    //AXI-MM pass-through interface 33
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_33_AWADDR,
    input wire [7:0]                      AP_AXIMM_33_AWLEN,
    input wire [2:0]                      AP_AXIMM_33_AWSIZE,
    input wire [1:0]                      AP_AXIMM_33_AWBURST,
    input wire [1:0]                      AP_AXIMM_33_AWLOCK,
    input wire [3:0]                      AP_AXIMM_33_AWCACHE,
    input wire [2:0]                      AP_AXIMM_33_AWPROT,
    input wire [3:0]                      AP_AXIMM_33_AWREGION,
    input wire [3:0]                      AP_AXIMM_33_AWQOS,
    input wire                            AP_AXIMM_33_AWVALID,
    output  wire                            AP_AXIMM_33_AWREADY,
    input wire [M_AXIMM_33_DATA_WIDTH-1:0]   AP_AXIMM_33_WDATA,
    input wire [M_AXIMM_33_DATA_WIDTH/8-1:0] AP_AXIMM_33_WSTRB,
    input wire                            AP_AXIMM_33_WLAST,
    input wire                            AP_AXIMM_33_WVALID,
    output  wire                            AP_AXIMM_33_WREADY,
    output  wire [1:0]                      AP_AXIMM_33_BRESP,
    output  wire                            AP_AXIMM_33_BVALID,
    input wire                            AP_AXIMM_33_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_33_ARADDR,
    input wire [7:0]                      AP_AXIMM_33_ARLEN,
    input wire [2:0]                      AP_AXIMM_33_ARSIZE,
    input wire [1:0]                      AP_AXIMM_33_ARBURST,
    input wire [1:0]                      AP_AXIMM_33_ARLOCK,
    input wire [3:0]                      AP_AXIMM_33_ARCACHE,
    input wire [2:0]                      AP_AXIMM_33_ARPROT,
    input wire [3:0]                      AP_AXIMM_33_ARREGION,
    input wire [3:0]                      AP_AXIMM_33_ARQOS,
    input wire                            AP_AXIMM_33_ARVALID,
    output  wire                            AP_AXIMM_33_ARREADY,
    output  wire [M_AXIMM_33_DATA_WIDTH-1:0]   AP_AXIMM_33_RDATA,
    output  wire [1:0]                      AP_AXIMM_33_RRESP,
    output  wire                            AP_AXIMM_33_RLAST,
    output  wire                            AP_AXIMM_33_RVALID,
    input  wire                            AP_AXIMM_33_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_33_AWADDR,
    output wire [7:0]                      M_AXIMM_33_AWLEN,
    output wire [2:0]                      M_AXIMM_33_AWSIZE,
    output wire [1:0]                      M_AXIMM_33_AWBURST,
    output wire [1:0]                      M_AXIMM_33_AWLOCK,
    output wire [3:0]                      M_AXIMM_33_AWCACHE,
    output wire [2:0]                      M_AXIMM_33_AWPROT,
    output wire [3:0]                      M_AXIMM_33_AWREGION,
    output wire [3:0]                      M_AXIMM_33_AWQOS,
    output wire                            M_AXIMM_33_AWVALID,
    input  wire                            M_AXIMM_33_AWREADY,
    output wire [M_AXIMM_33_DATA_WIDTH-1:0]   M_AXIMM_33_WDATA,
    output wire [M_AXIMM_33_DATA_WIDTH/8-1:0] M_AXIMM_33_WSTRB,
    output wire                            M_AXIMM_33_WLAST,
    output wire                            M_AXIMM_33_WVALID,
    input  wire                            M_AXIMM_33_WREADY,
    input  wire [1:0]                      M_AXIMM_33_BRESP,
    input  wire                            M_AXIMM_33_BVALID,
    output wire                            M_AXIMM_33_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_33_ARADDR,
    output wire [7:0]                      M_AXIMM_33_ARLEN,
    output wire [2:0]                      M_AXIMM_33_ARSIZE,
    output wire [1:0]                      M_AXIMM_33_ARBURST,
    output wire [1:0]                      M_AXIMM_33_ARLOCK,
    output wire [3:0]                      M_AXIMM_33_ARCACHE,
    output wire [2:0]                      M_AXIMM_33_ARPROT,
    output wire [3:0]                      M_AXIMM_33_ARREGION,
    output wire [3:0]                      M_AXIMM_33_ARQOS,
    output wire                            M_AXIMM_33_ARVALID,
    input  wire                            M_AXIMM_33_ARREADY,
    input  wire [M_AXIMM_33_DATA_WIDTH-1:0]   M_AXIMM_33_RDATA,
    input  wire [1:0]                      M_AXIMM_33_RRESP,
    input  wire                            M_AXIMM_33_RLAST,
    input  wire                            M_AXIMM_33_RVALID,
    output wire                            M_AXIMM_33_RREADY,
    //AXI-MM pass-through interface 34
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_34_AWADDR,
    input wire [7:0]                      AP_AXIMM_34_AWLEN,
    input wire [2:0]                      AP_AXIMM_34_AWSIZE,
    input wire [1:0]                      AP_AXIMM_34_AWBURST,
    input wire [1:0]                      AP_AXIMM_34_AWLOCK,
    input wire [3:0]                      AP_AXIMM_34_AWCACHE,
    input wire [2:0]                      AP_AXIMM_34_AWPROT,
    input wire [3:0]                      AP_AXIMM_34_AWREGION,
    input wire [3:0]                      AP_AXIMM_34_AWQOS,
    input wire                            AP_AXIMM_34_AWVALID,
    output  wire                            AP_AXIMM_34_AWREADY,
    input wire [M_AXIMM_34_DATA_WIDTH-1:0]   AP_AXIMM_34_WDATA,
    input wire [M_AXIMM_34_DATA_WIDTH/8-1:0] AP_AXIMM_34_WSTRB,
    input wire                            AP_AXIMM_34_WLAST,
    input wire                            AP_AXIMM_34_WVALID,
    output  wire                            AP_AXIMM_34_WREADY,
    output  wire [1:0]                      AP_AXIMM_34_BRESP,
    output  wire                            AP_AXIMM_34_BVALID,
    input wire                            AP_AXIMM_34_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_34_ARADDR,
    input wire [7:0]                      AP_AXIMM_34_ARLEN,
    input wire [2:0]                      AP_AXIMM_34_ARSIZE,
    input wire [1:0]                      AP_AXIMM_34_ARBURST,
    input wire [1:0]                      AP_AXIMM_34_ARLOCK,
    input wire [3:0]                      AP_AXIMM_34_ARCACHE,
    input wire [2:0]                      AP_AXIMM_34_ARPROT,
    input wire [3:0]                      AP_AXIMM_34_ARREGION,
    input wire [3:0]                      AP_AXIMM_34_ARQOS,
    input wire                            AP_AXIMM_34_ARVALID,
    output  wire                            AP_AXIMM_34_ARREADY,
    output  wire [M_AXIMM_34_DATA_WIDTH-1:0]   AP_AXIMM_34_RDATA,
    output  wire [1:0]                      AP_AXIMM_34_RRESP,
    output  wire                            AP_AXIMM_34_RLAST,
    output  wire                            AP_AXIMM_34_RVALID,
    input  wire                            AP_AXIMM_34_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_34_AWADDR,
    output wire [7:0]                      M_AXIMM_34_AWLEN,
    output wire [2:0]                      M_AXIMM_34_AWSIZE,
    output wire [1:0]                      M_AXIMM_34_AWBURST,
    output wire [1:0]                      M_AXIMM_34_AWLOCK,
    output wire [3:0]                      M_AXIMM_34_AWCACHE,
    output wire [2:0]                      M_AXIMM_34_AWPROT,
    output wire [3:0]                      M_AXIMM_34_AWREGION,
    output wire [3:0]                      M_AXIMM_34_AWQOS,
    output wire                            M_AXIMM_34_AWVALID,
    input  wire                            M_AXIMM_34_AWREADY,
    output wire [M_AXIMM_34_DATA_WIDTH-1:0]   M_AXIMM_34_WDATA,
    output wire [M_AXIMM_34_DATA_WIDTH/8-1:0] M_AXIMM_34_WSTRB,
    output wire                            M_AXIMM_34_WLAST,
    output wire                            M_AXIMM_34_WVALID,
    input  wire                            M_AXIMM_34_WREADY,
    input  wire [1:0]                      M_AXIMM_34_BRESP,
    input  wire                            M_AXIMM_34_BVALID,
    output wire                            M_AXIMM_34_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_34_ARADDR,
    output wire [7:0]                      M_AXIMM_34_ARLEN,
    output wire [2:0]                      M_AXIMM_34_ARSIZE,
    output wire [1:0]                      M_AXIMM_34_ARBURST,
    output wire [1:0]                      M_AXIMM_34_ARLOCK,
    output wire [3:0]                      M_AXIMM_34_ARCACHE,
    output wire [2:0]                      M_AXIMM_34_ARPROT,
    output wire [3:0]                      M_AXIMM_34_ARREGION,
    output wire [3:0]                      M_AXIMM_34_ARQOS,
    output wire                            M_AXIMM_34_ARVALID,
    input  wire                            M_AXIMM_34_ARREADY,
    input  wire [M_AXIMM_34_DATA_WIDTH-1:0]   M_AXIMM_34_RDATA,
    input  wire [1:0]                      M_AXIMM_34_RRESP,
    input  wire                            M_AXIMM_34_RLAST,
    input  wire                            M_AXIMM_34_RVALID,
    output wire                            M_AXIMM_34_RREADY,
    //AXI-MM pass-through interface 35
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_35_AWADDR,
    input wire [7:0]                      AP_AXIMM_35_AWLEN,
    input wire [2:0]                      AP_AXIMM_35_AWSIZE,
    input wire [1:0]                      AP_AXIMM_35_AWBURST,
    input wire [1:0]                      AP_AXIMM_35_AWLOCK,
    input wire [3:0]                      AP_AXIMM_35_AWCACHE,
    input wire [2:0]                      AP_AXIMM_35_AWPROT,
    input wire [3:0]                      AP_AXIMM_35_AWREGION,
    input wire [3:0]                      AP_AXIMM_35_AWQOS,
    input wire                            AP_AXIMM_35_AWVALID,
    output  wire                            AP_AXIMM_35_AWREADY,
    input wire [M_AXIMM_35_DATA_WIDTH-1:0]   AP_AXIMM_35_WDATA,
    input wire [M_AXIMM_35_DATA_WIDTH/8-1:0] AP_AXIMM_35_WSTRB,
    input wire                            AP_AXIMM_35_WLAST,
    input wire                            AP_AXIMM_35_WVALID,
    output  wire                            AP_AXIMM_35_WREADY,
    output  wire [1:0]                      AP_AXIMM_35_BRESP,
    output  wire                            AP_AXIMM_35_BVALID,
    input wire                            AP_AXIMM_35_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_35_ARADDR,
    input wire [7:0]                      AP_AXIMM_35_ARLEN,
    input wire [2:0]                      AP_AXIMM_35_ARSIZE,
    input wire [1:0]                      AP_AXIMM_35_ARBURST,
    input wire [1:0]                      AP_AXIMM_35_ARLOCK,
    input wire [3:0]                      AP_AXIMM_35_ARCACHE,
    input wire [2:0]                      AP_AXIMM_35_ARPROT,
    input wire [3:0]                      AP_AXIMM_35_ARREGION,
    input wire [3:0]                      AP_AXIMM_35_ARQOS,
    input wire                            AP_AXIMM_35_ARVALID,
    output  wire                            AP_AXIMM_35_ARREADY,
    output  wire [M_AXIMM_35_DATA_WIDTH-1:0]   AP_AXIMM_35_RDATA,
    output  wire [1:0]                      AP_AXIMM_35_RRESP,
    output  wire                            AP_AXIMM_35_RLAST,
    output  wire                            AP_AXIMM_35_RVALID,
    input  wire                            AP_AXIMM_35_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_35_AWADDR,
    output wire [7:0]                      M_AXIMM_35_AWLEN,
    output wire [2:0]                      M_AXIMM_35_AWSIZE,
    output wire [1:0]                      M_AXIMM_35_AWBURST,
    output wire [1:0]                      M_AXIMM_35_AWLOCK,
    output wire [3:0]                      M_AXIMM_35_AWCACHE,
    output wire [2:0]                      M_AXIMM_35_AWPROT,
    output wire [3:0]                      M_AXIMM_35_AWREGION,
    output wire [3:0]                      M_AXIMM_35_AWQOS,
    output wire                            M_AXIMM_35_AWVALID,
    input  wire                            M_AXIMM_35_AWREADY,
    output wire [M_AXIMM_35_DATA_WIDTH-1:0]   M_AXIMM_35_WDATA,
    output wire [M_AXIMM_35_DATA_WIDTH/8-1:0] M_AXIMM_35_WSTRB,
    output wire                            M_AXIMM_35_WLAST,
    output wire                            M_AXIMM_35_WVALID,
    input  wire                            M_AXIMM_35_WREADY,
    input  wire [1:0]                      M_AXIMM_35_BRESP,
    input  wire                            M_AXIMM_35_BVALID,
    output wire                            M_AXIMM_35_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_35_ARADDR,
    output wire [7:0]                      M_AXIMM_35_ARLEN,
    output wire [2:0]                      M_AXIMM_35_ARSIZE,
    output wire [1:0]                      M_AXIMM_35_ARBURST,
    output wire [1:0]                      M_AXIMM_35_ARLOCK,
    output wire [3:0]                      M_AXIMM_35_ARCACHE,
    output wire [2:0]                      M_AXIMM_35_ARPROT,
    output wire [3:0]                      M_AXIMM_35_ARREGION,
    output wire [3:0]                      M_AXIMM_35_ARQOS,
    output wire                            M_AXIMM_35_ARVALID,
    input  wire                            M_AXIMM_35_ARREADY,
    input  wire [M_AXIMM_35_DATA_WIDTH-1:0]   M_AXIMM_35_RDATA,
    input  wire [1:0]                      M_AXIMM_35_RRESP,
    input  wire                            M_AXIMM_35_RLAST,
    input  wire                            M_AXIMM_35_RVALID,
    output wire                            M_AXIMM_35_RREADY,
    //AXI-MM pass-through interface 36
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_36_AWADDR,
    input wire [7:0]                      AP_AXIMM_36_AWLEN,
    input wire [2:0]                      AP_AXIMM_36_AWSIZE,
    input wire [1:0]                      AP_AXIMM_36_AWBURST,
    input wire [1:0]                      AP_AXIMM_36_AWLOCK,
    input wire [3:0]                      AP_AXIMM_36_AWCACHE,
    input wire [2:0]                      AP_AXIMM_36_AWPROT,
    input wire [3:0]                      AP_AXIMM_36_AWREGION,
    input wire [3:0]                      AP_AXIMM_36_AWQOS,
    input wire                            AP_AXIMM_36_AWVALID,
    output  wire                            AP_AXIMM_36_AWREADY,
    input wire [M_AXIMM_36_DATA_WIDTH-1:0]   AP_AXIMM_36_WDATA,
    input wire [M_AXIMM_36_DATA_WIDTH/8-1:0] AP_AXIMM_36_WSTRB,
    input wire                            AP_AXIMM_36_WLAST,
    input wire                            AP_AXIMM_36_WVALID,
    output  wire                            AP_AXIMM_36_WREADY,
    output  wire [1:0]                      AP_AXIMM_36_BRESP,
    output  wire                            AP_AXIMM_36_BVALID,
    input wire                            AP_AXIMM_36_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_36_ARADDR,
    input wire [7:0]                      AP_AXIMM_36_ARLEN,
    input wire [2:0]                      AP_AXIMM_36_ARSIZE,
    input wire [1:0]                      AP_AXIMM_36_ARBURST,
    input wire [1:0]                      AP_AXIMM_36_ARLOCK,
    input wire [3:0]                      AP_AXIMM_36_ARCACHE,
    input wire [2:0]                      AP_AXIMM_36_ARPROT,
    input wire [3:0]                      AP_AXIMM_36_ARREGION,
    input wire [3:0]                      AP_AXIMM_36_ARQOS,
    input wire                            AP_AXIMM_36_ARVALID,
    output  wire                            AP_AXIMM_36_ARREADY,
    output  wire [M_AXIMM_36_DATA_WIDTH-1:0]   AP_AXIMM_36_RDATA,
    output  wire [1:0]                      AP_AXIMM_36_RRESP,
    output  wire                            AP_AXIMM_36_RLAST,
    output  wire                            AP_AXIMM_36_RVALID,
    input  wire                            AP_AXIMM_36_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_36_AWADDR,
    output wire [7:0]                      M_AXIMM_36_AWLEN,
    output wire [2:0]                      M_AXIMM_36_AWSIZE,
    output wire [1:0]                      M_AXIMM_36_AWBURST,
    output wire [1:0]                      M_AXIMM_36_AWLOCK,
    output wire [3:0]                      M_AXIMM_36_AWCACHE,
    output wire [2:0]                      M_AXIMM_36_AWPROT,
    output wire [3:0]                      M_AXIMM_36_AWREGION,
    output wire [3:0]                      M_AXIMM_36_AWQOS,
    output wire                            M_AXIMM_36_AWVALID,
    input  wire                            M_AXIMM_36_AWREADY,
    output wire [M_AXIMM_36_DATA_WIDTH-1:0]   M_AXIMM_36_WDATA,
    output wire [M_AXIMM_36_DATA_WIDTH/8-1:0] M_AXIMM_36_WSTRB,
    output wire                            M_AXIMM_36_WLAST,
    output wire                            M_AXIMM_36_WVALID,
    input  wire                            M_AXIMM_36_WREADY,
    input  wire [1:0]                      M_AXIMM_36_BRESP,
    input  wire                            M_AXIMM_36_BVALID,
    output wire                            M_AXIMM_36_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_36_ARADDR,
    output wire [7:0]                      M_AXIMM_36_ARLEN,
    output wire [2:0]                      M_AXIMM_36_ARSIZE,
    output wire [1:0]                      M_AXIMM_36_ARBURST,
    output wire [1:0]                      M_AXIMM_36_ARLOCK,
    output wire [3:0]                      M_AXIMM_36_ARCACHE,
    output wire [2:0]                      M_AXIMM_36_ARPROT,
    output wire [3:0]                      M_AXIMM_36_ARREGION,
    output wire [3:0]                      M_AXIMM_36_ARQOS,
    output wire                            M_AXIMM_36_ARVALID,
    input  wire                            M_AXIMM_36_ARREADY,
    input  wire [M_AXIMM_36_DATA_WIDTH-1:0]   M_AXIMM_36_RDATA,
    input  wire [1:0]                      M_AXIMM_36_RRESP,
    input  wire                            M_AXIMM_36_RLAST,
    input  wire                            M_AXIMM_36_RVALID,
    output wire                            M_AXIMM_36_RREADY,
    //AXI-MM pass-through interface 37
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_37_AWADDR,
    input wire [7:0]                      AP_AXIMM_37_AWLEN,
    input wire [2:0]                      AP_AXIMM_37_AWSIZE,
    input wire [1:0]                      AP_AXIMM_37_AWBURST,
    input wire [1:0]                      AP_AXIMM_37_AWLOCK,
    input wire [3:0]                      AP_AXIMM_37_AWCACHE,
    input wire [2:0]                      AP_AXIMM_37_AWPROT,
    input wire [3:0]                      AP_AXIMM_37_AWREGION,
    input wire [3:0]                      AP_AXIMM_37_AWQOS,
    input wire                            AP_AXIMM_37_AWVALID,
    output  wire                            AP_AXIMM_37_AWREADY,
    input wire [M_AXIMM_37_DATA_WIDTH-1:0]   AP_AXIMM_37_WDATA,
    input wire [M_AXIMM_37_DATA_WIDTH/8-1:0] AP_AXIMM_37_WSTRB,
    input wire                            AP_AXIMM_37_WLAST,
    input wire                            AP_AXIMM_37_WVALID,
    output  wire                            AP_AXIMM_37_WREADY,
    output  wire [1:0]                      AP_AXIMM_37_BRESP,
    output  wire                            AP_AXIMM_37_BVALID,
    input wire                            AP_AXIMM_37_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_37_ARADDR,
    input wire [7:0]                      AP_AXIMM_37_ARLEN,
    input wire [2:0]                      AP_AXIMM_37_ARSIZE,
    input wire [1:0]                      AP_AXIMM_37_ARBURST,
    input wire [1:0]                      AP_AXIMM_37_ARLOCK,
    input wire [3:0]                      AP_AXIMM_37_ARCACHE,
    input wire [2:0]                      AP_AXIMM_37_ARPROT,
    input wire [3:0]                      AP_AXIMM_37_ARREGION,
    input wire [3:0]                      AP_AXIMM_37_ARQOS,
    input wire                            AP_AXIMM_37_ARVALID,
    output  wire                            AP_AXIMM_37_ARREADY,
    output  wire [M_AXIMM_37_DATA_WIDTH-1:0]   AP_AXIMM_37_RDATA,
    output  wire [1:0]                      AP_AXIMM_37_RRESP,
    output  wire                            AP_AXIMM_37_RLAST,
    output  wire                            AP_AXIMM_37_RVALID,
    input  wire                            AP_AXIMM_37_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_37_AWADDR,
    output wire [7:0]                      M_AXIMM_37_AWLEN,
    output wire [2:0]                      M_AXIMM_37_AWSIZE,
    output wire [1:0]                      M_AXIMM_37_AWBURST,
    output wire [1:0]                      M_AXIMM_37_AWLOCK,
    output wire [3:0]                      M_AXIMM_37_AWCACHE,
    output wire [2:0]                      M_AXIMM_37_AWPROT,
    output wire [3:0]                      M_AXIMM_37_AWREGION,
    output wire [3:0]                      M_AXIMM_37_AWQOS,
    output wire                            M_AXIMM_37_AWVALID,
    input  wire                            M_AXIMM_37_AWREADY,
    output wire [M_AXIMM_37_DATA_WIDTH-1:0]   M_AXIMM_37_WDATA,
    output wire [M_AXIMM_37_DATA_WIDTH/8-1:0] M_AXIMM_37_WSTRB,
    output wire                            M_AXIMM_37_WLAST,
    output wire                            M_AXIMM_37_WVALID,
    input  wire                            M_AXIMM_37_WREADY,
    input  wire [1:0]                      M_AXIMM_37_BRESP,
    input  wire                            M_AXIMM_37_BVALID,
    output wire                            M_AXIMM_37_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_37_ARADDR,
    output wire [7:0]                      M_AXIMM_37_ARLEN,
    output wire [2:0]                      M_AXIMM_37_ARSIZE,
    output wire [1:0]                      M_AXIMM_37_ARBURST,
    output wire [1:0]                      M_AXIMM_37_ARLOCK,
    output wire [3:0]                      M_AXIMM_37_ARCACHE,
    output wire [2:0]                      M_AXIMM_37_ARPROT,
    output wire [3:0]                      M_AXIMM_37_ARREGION,
    output wire [3:0]                      M_AXIMM_37_ARQOS,
    output wire                            M_AXIMM_37_ARVALID,
    input  wire                            M_AXIMM_37_ARREADY,
    input  wire [M_AXIMM_37_DATA_WIDTH-1:0]   M_AXIMM_37_RDATA,
    input  wire [1:0]                      M_AXIMM_37_RRESP,
    input  wire                            M_AXIMM_37_RLAST,
    input  wire                            M_AXIMM_37_RVALID,
    output wire                            M_AXIMM_37_RREADY,
    //AXI-MM pass-through interface 38
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_38_AWADDR,
    input wire [7:0]                      AP_AXIMM_38_AWLEN,
    input wire [2:0]                      AP_AXIMM_38_AWSIZE,
    input wire [1:0]                      AP_AXIMM_38_AWBURST,
    input wire [1:0]                      AP_AXIMM_38_AWLOCK,
    input wire [3:0]                      AP_AXIMM_38_AWCACHE,
    input wire [2:0]                      AP_AXIMM_38_AWPROT,
    input wire [3:0]                      AP_AXIMM_38_AWREGION,
    input wire [3:0]                      AP_AXIMM_38_AWQOS,
    input wire                            AP_AXIMM_38_AWVALID,
    output  wire                            AP_AXIMM_38_AWREADY,
    input wire [M_AXIMM_38_DATA_WIDTH-1:0]   AP_AXIMM_38_WDATA,
    input wire [M_AXIMM_38_DATA_WIDTH/8-1:0] AP_AXIMM_38_WSTRB,
    input wire                            AP_AXIMM_38_WLAST,
    input wire                            AP_AXIMM_38_WVALID,
    output  wire                            AP_AXIMM_38_WREADY,
    output  wire [1:0]                      AP_AXIMM_38_BRESP,
    output  wire                            AP_AXIMM_38_BVALID,
    input wire                            AP_AXIMM_38_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_38_ARADDR,
    input wire [7:0]                      AP_AXIMM_38_ARLEN,
    input wire [2:0]                      AP_AXIMM_38_ARSIZE,
    input wire [1:0]                      AP_AXIMM_38_ARBURST,
    input wire [1:0]                      AP_AXIMM_38_ARLOCK,
    input wire [3:0]                      AP_AXIMM_38_ARCACHE,
    input wire [2:0]                      AP_AXIMM_38_ARPROT,
    input wire [3:0]                      AP_AXIMM_38_ARREGION,
    input wire [3:0]                      AP_AXIMM_38_ARQOS,
    input wire                            AP_AXIMM_38_ARVALID,
    output  wire                            AP_AXIMM_38_ARREADY,
    output  wire [M_AXIMM_38_DATA_WIDTH-1:0]   AP_AXIMM_38_RDATA,
    output  wire [1:0]                      AP_AXIMM_38_RRESP,
    output  wire                            AP_AXIMM_38_RLAST,
    output  wire                            AP_AXIMM_38_RVALID,
    input  wire                            AP_AXIMM_38_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_38_AWADDR,
    output wire [7:0]                      M_AXIMM_38_AWLEN,
    output wire [2:0]                      M_AXIMM_38_AWSIZE,
    output wire [1:0]                      M_AXIMM_38_AWBURST,
    output wire [1:0]                      M_AXIMM_38_AWLOCK,
    output wire [3:0]                      M_AXIMM_38_AWCACHE,
    output wire [2:0]                      M_AXIMM_38_AWPROT,
    output wire [3:0]                      M_AXIMM_38_AWREGION,
    output wire [3:0]                      M_AXIMM_38_AWQOS,
    output wire                            M_AXIMM_38_AWVALID,
    input  wire                            M_AXIMM_38_AWREADY,
    output wire [M_AXIMM_38_DATA_WIDTH-1:0]   M_AXIMM_38_WDATA,
    output wire [M_AXIMM_38_DATA_WIDTH/8-1:0] M_AXIMM_38_WSTRB,
    output wire                            M_AXIMM_38_WLAST,
    output wire                            M_AXIMM_38_WVALID,
    input  wire                            M_AXIMM_38_WREADY,
    input  wire [1:0]                      M_AXIMM_38_BRESP,
    input  wire                            M_AXIMM_38_BVALID,
    output wire                            M_AXIMM_38_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_38_ARADDR,
    output wire [7:0]                      M_AXIMM_38_ARLEN,
    output wire [2:0]                      M_AXIMM_38_ARSIZE,
    output wire [1:0]                      M_AXIMM_38_ARBURST,
    output wire [1:0]                      M_AXIMM_38_ARLOCK,
    output wire [3:0]                      M_AXIMM_38_ARCACHE,
    output wire [2:0]                      M_AXIMM_38_ARPROT,
    output wire [3:0]                      M_AXIMM_38_ARREGION,
    output wire [3:0]                      M_AXIMM_38_ARQOS,
    output wire                            M_AXIMM_38_ARVALID,
    input  wire                            M_AXIMM_38_ARREADY,
    input  wire [M_AXIMM_38_DATA_WIDTH-1:0]   M_AXIMM_38_RDATA,
    input  wire [1:0]                      M_AXIMM_38_RRESP,
    input  wire                            M_AXIMM_38_RLAST,
    input  wire                            M_AXIMM_38_RVALID,
    output wire                            M_AXIMM_38_RREADY,
    //AXI-MM pass-through interface 39
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_39_AWADDR,
    input wire [7:0]                      AP_AXIMM_39_AWLEN,
    input wire [2:0]                      AP_AXIMM_39_AWSIZE,
    input wire [1:0]                      AP_AXIMM_39_AWBURST,
    input wire [1:0]                      AP_AXIMM_39_AWLOCK,
    input wire [3:0]                      AP_AXIMM_39_AWCACHE,
    input wire [2:0]                      AP_AXIMM_39_AWPROT,
    input wire [3:0]                      AP_AXIMM_39_AWREGION,
    input wire [3:0]                      AP_AXIMM_39_AWQOS,
    input wire                            AP_AXIMM_39_AWVALID,
    output  wire                            AP_AXIMM_39_AWREADY,
    input wire [M_AXIMM_39_DATA_WIDTH-1:0]   AP_AXIMM_39_WDATA,
    input wire [M_AXIMM_39_DATA_WIDTH/8-1:0] AP_AXIMM_39_WSTRB,
    input wire                            AP_AXIMM_39_WLAST,
    input wire                            AP_AXIMM_39_WVALID,
    output  wire                            AP_AXIMM_39_WREADY,
    output  wire [1:0]                      AP_AXIMM_39_BRESP,
    output  wire                            AP_AXIMM_39_BVALID,
    input wire                            AP_AXIMM_39_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_39_ARADDR,
    input wire [7:0]                      AP_AXIMM_39_ARLEN,
    input wire [2:0]                      AP_AXIMM_39_ARSIZE,
    input wire [1:0]                      AP_AXIMM_39_ARBURST,
    input wire [1:0]                      AP_AXIMM_39_ARLOCK,
    input wire [3:0]                      AP_AXIMM_39_ARCACHE,
    input wire [2:0]                      AP_AXIMM_39_ARPROT,
    input wire [3:0]                      AP_AXIMM_39_ARREGION,
    input wire [3:0]                      AP_AXIMM_39_ARQOS,
    input wire                            AP_AXIMM_39_ARVALID,
    output  wire                            AP_AXIMM_39_ARREADY,
    output  wire [M_AXIMM_39_DATA_WIDTH-1:0]   AP_AXIMM_39_RDATA,
    output  wire [1:0]                      AP_AXIMM_39_RRESP,
    output  wire                            AP_AXIMM_39_RLAST,
    output  wire                            AP_AXIMM_39_RVALID,
    input  wire                            AP_AXIMM_39_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_39_AWADDR,
    output wire [7:0]                      M_AXIMM_39_AWLEN,
    output wire [2:0]                      M_AXIMM_39_AWSIZE,
    output wire [1:0]                      M_AXIMM_39_AWBURST,
    output wire [1:0]                      M_AXIMM_39_AWLOCK,
    output wire [3:0]                      M_AXIMM_39_AWCACHE,
    output wire [2:0]                      M_AXIMM_39_AWPROT,
    output wire [3:0]                      M_AXIMM_39_AWREGION,
    output wire [3:0]                      M_AXIMM_39_AWQOS,
    output wire                            M_AXIMM_39_AWVALID,
    input  wire                            M_AXIMM_39_AWREADY,
    output wire [M_AXIMM_39_DATA_WIDTH-1:0]   M_AXIMM_39_WDATA,
    output wire [M_AXIMM_39_DATA_WIDTH/8-1:0] M_AXIMM_39_WSTRB,
    output wire                            M_AXIMM_39_WLAST,
    output wire                            M_AXIMM_39_WVALID,
    input  wire                            M_AXIMM_39_WREADY,
    input  wire [1:0]                      M_AXIMM_39_BRESP,
    input  wire                            M_AXIMM_39_BVALID,
    output wire                            M_AXIMM_39_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_39_ARADDR,
    output wire [7:0]                      M_AXIMM_39_ARLEN,
    output wire [2:0]                      M_AXIMM_39_ARSIZE,
    output wire [1:0]                      M_AXIMM_39_ARBURST,
    output wire [1:0]                      M_AXIMM_39_ARLOCK,
    output wire [3:0]                      M_AXIMM_39_ARCACHE,
    output wire [2:0]                      M_AXIMM_39_ARPROT,
    output wire [3:0]                      M_AXIMM_39_ARREGION,
    output wire [3:0]                      M_AXIMM_39_ARQOS,
    output wire                            M_AXIMM_39_ARVALID,
    input  wire                            M_AXIMM_39_ARREADY,
    input  wire [M_AXIMM_39_DATA_WIDTH-1:0]   M_AXIMM_39_RDATA,
    input  wire [1:0]                      M_AXIMM_39_RRESP,
    input  wire                            M_AXIMM_39_RLAST,
    input  wire                            M_AXIMM_39_RVALID,
    output wire                            M_AXIMM_39_RREADY,
    //AXI-MM pass-through interface 40
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_40_AWADDR,
    input wire [7:0]                      AP_AXIMM_40_AWLEN,
    input wire [2:0]                      AP_AXIMM_40_AWSIZE,
    input wire [1:0]                      AP_AXIMM_40_AWBURST,
    input wire [1:0]                      AP_AXIMM_40_AWLOCK,
    input wire [3:0]                      AP_AXIMM_40_AWCACHE,
    input wire [2:0]                      AP_AXIMM_40_AWPROT,
    input wire [3:0]                      AP_AXIMM_40_AWREGION,
    input wire [3:0]                      AP_AXIMM_40_AWQOS,
    input wire                            AP_AXIMM_40_AWVALID,
    output  wire                            AP_AXIMM_40_AWREADY,
    input wire [M_AXIMM_40_DATA_WIDTH-1:0]   AP_AXIMM_40_WDATA,
    input wire [M_AXIMM_40_DATA_WIDTH/8-1:0] AP_AXIMM_40_WSTRB,
    input wire                            AP_AXIMM_40_WLAST,
    input wire                            AP_AXIMM_40_WVALID,
    output  wire                            AP_AXIMM_40_WREADY,
    output  wire [1:0]                      AP_AXIMM_40_BRESP,
    output  wire                            AP_AXIMM_40_BVALID,
    input wire                            AP_AXIMM_40_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_40_ARADDR,
    input wire [7:0]                      AP_AXIMM_40_ARLEN,
    input wire [2:0]                      AP_AXIMM_40_ARSIZE,
    input wire [1:0]                      AP_AXIMM_40_ARBURST,
    input wire [1:0]                      AP_AXIMM_40_ARLOCK,
    input wire [3:0]                      AP_AXIMM_40_ARCACHE,
    input wire [2:0]                      AP_AXIMM_40_ARPROT,
    input wire [3:0]                      AP_AXIMM_40_ARREGION,
    input wire [3:0]                      AP_AXIMM_40_ARQOS,
    input wire                            AP_AXIMM_40_ARVALID,
    output  wire                            AP_AXIMM_40_ARREADY,
    output  wire [M_AXIMM_40_DATA_WIDTH-1:0]   AP_AXIMM_40_RDATA,
    output  wire [1:0]                      AP_AXIMM_40_RRESP,
    output  wire                            AP_AXIMM_40_RLAST,
    output  wire                            AP_AXIMM_40_RVALID,
    input  wire                            AP_AXIMM_40_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_40_AWADDR,
    output wire [7:0]                      M_AXIMM_40_AWLEN,
    output wire [2:0]                      M_AXIMM_40_AWSIZE,
    output wire [1:0]                      M_AXIMM_40_AWBURST,
    output wire [1:0]                      M_AXIMM_40_AWLOCK,
    output wire [3:0]                      M_AXIMM_40_AWCACHE,
    output wire [2:0]                      M_AXIMM_40_AWPROT,
    output wire [3:0]                      M_AXIMM_40_AWREGION,
    output wire [3:0]                      M_AXIMM_40_AWQOS,
    output wire                            M_AXIMM_40_AWVALID,
    input  wire                            M_AXIMM_40_AWREADY,
    output wire [M_AXIMM_40_DATA_WIDTH-1:0]   M_AXIMM_40_WDATA,
    output wire [M_AXIMM_40_DATA_WIDTH/8-1:0] M_AXIMM_40_WSTRB,
    output wire                            M_AXIMM_40_WLAST,
    output wire                            M_AXIMM_40_WVALID,
    input  wire                            M_AXIMM_40_WREADY,
    input  wire [1:0]                      M_AXIMM_40_BRESP,
    input  wire                            M_AXIMM_40_BVALID,
    output wire                            M_AXIMM_40_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_40_ARADDR,
    output wire [7:0]                      M_AXIMM_40_ARLEN,
    output wire [2:0]                      M_AXIMM_40_ARSIZE,
    output wire [1:0]                      M_AXIMM_40_ARBURST,
    output wire [1:0]                      M_AXIMM_40_ARLOCK,
    output wire [3:0]                      M_AXIMM_40_ARCACHE,
    output wire [2:0]                      M_AXIMM_40_ARPROT,
    output wire [3:0]                      M_AXIMM_40_ARREGION,
    output wire [3:0]                      M_AXIMM_40_ARQOS,
    output wire                            M_AXIMM_40_ARVALID,
    input  wire                            M_AXIMM_40_ARREADY,
    input  wire [M_AXIMM_40_DATA_WIDTH-1:0]   M_AXIMM_40_RDATA,
    input  wire [1:0]                      M_AXIMM_40_RRESP,
    input  wire                            M_AXIMM_40_RLAST,
    input  wire                            M_AXIMM_40_RVALID,
    output wire                            M_AXIMM_40_RREADY,
    //AXI-MM pass-through interface 41
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_41_AWADDR,
    input wire [7:0]                      AP_AXIMM_41_AWLEN,
    input wire [2:0]                      AP_AXIMM_41_AWSIZE,
    input wire [1:0]                      AP_AXIMM_41_AWBURST,
    input wire [1:0]                      AP_AXIMM_41_AWLOCK,
    input wire [3:0]                      AP_AXIMM_41_AWCACHE,
    input wire [2:0]                      AP_AXIMM_41_AWPROT,
    input wire [3:0]                      AP_AXIMM_41_AWREGION,
    input wire [3:0]                      AP_AXIMM_41_AWQOS,
    input wire                            AP_AXIMM_41_AWVALID,
    output  wire                            AP_AXIMM_41_AWREADY,
    input wire [M_AXIMM_41_DATA_WIDTH-1:0]   AP_AXIMM_41_WDATA,
    input wire [M_AXIMM_41_DATA_WIDTH/8-1:0] AP_AXIMM_41_WSTRB,
    input wire                            AP_AXIMM_41_WLAST,
    input wire                            AP_AXIMM_41_WVALID,
    output  wire                            AP_AXIMM_41_WREADY,
    output  wire [1:0]                      AP_AXIMM_41_BRESP,
    output  wire                            AP_AXIMM_41_BVALID,
    input wire                            AP_AXIMM_41_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_41_ARADDR,
    input wire [7:0]                      AP_AXIMM_41_ARLEN,
    input wire [2:0]                      AP_AXIMM_41_ARSIZE,
    input wire [1:0]                      AP_AXIMM_41_ARBURST,
    input wire [1:0]                      AP_AXIMM_41_ARLOCK,
    input wire [3:0]                      AP_AXIMM_41_ARCACHE,
    input wire [2:0]                      AP_AXIMM_41_ARPROT,
    input wire [3:0]                      AP_AXIMM_41_ARREGION,
    input wire [3:0]                      AP_AXIMM_41_ARQOS,
    input wire                            AP_AXIMM_41_ARVALID,
    output  wire                            AP_AXIMM_41_ARREADY,
    output  wire [M_AXIMM_41_DATA_WIDTH-1:0]   AP_AXIMM_41_RDATA,
    output  wire [1:0]                      AP_AXIMM_41_RRESP,
    output  wire                            AP_AXIMM_41_RLAST,
    output  wire                            AP_AXIMM_41_RVALID,
    input  wire                            AP_AXIMM_41_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_41_AWADDR,
    output wire [7:0]                      M_AXIMM_41_AWLEN,
    output wire [2:0]                      M_AXIMM_41_AWSIZE,
    output wire [1:0]                      M_AXIMM_41_AWBURST,
    output wire [1:0]                      M_AXIMM_41_AWLOCK,
    output wire [3:0]                      M_AXIMM_41_AWCACHE,
    output wire [2:0]                      M_AXIMM_41_AWPROT,
    output wire [3:0]                      M_AXIMM_41_AWREGION,
    output wire [3:0]                      M_AXIMM_41_AWQOS,
    output wire                            M_AXIMM_41_AWVALID,
    input  wire                            M_AXIMM_41_AWREADY,
    output wire [M_AXIMM_41_DATA_WIDTH-1:0]   M_AXIMM_41_WDATA,
    output wire [M_AXIMM_41_DATA_WIDTH/8-1:0] M_AXIMM_41_WSTRB,
    output wire                            M_AXIMM_41_WLAST,
    output wire                            M_AXIMM_41_WVALID,
    input  wire                            M_AXIMM_41_WREADY,
    input  wire [1:0]                      M_AXIMM_41_BRESP,
    input  wire                            M_AXIMM_41_BVALID,
    output wire                            M_AXIMM_41_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_41_ARADDR,
    output wire [7:0]                      M_AXIMM_41_ARLEN,
    output wire [2:0]                      M_AXIMM_41_ARSIZE,
    output wire [1:0]                      M_AXIMM_41_ARBURST,
    output wire [1:0]                      M_AXIMM_41_ARLOCK,
    output wire [3:0]                      M_AXIMM_41_ARCACHE,
    output wire [2:0]                      M_AXIMM_41_ARPROT,
    output wire [3:0]                      M_AXIMM_41_ARREGION,
    output wire [3:0]                      M_AXIMM_41_ARQOS,
    output wire                            M_AXIMM_41_ARVALID,
    input  wire                            M_AXIMM_41_ARREADY,
    input  wire [M_AXIMM_41_DATA_WIDTH-1:0]   M_AXIMM_41_RDATA,
    input  wire [1:0]                      M_AXIMM_41_RRESP,
    input  wire                            M_AXIMM_41_RLAST,
    input  wire                            M_AXIMM_41_RVALID,
    output wire                            M_AXIMM_41_RREADY,
    //AXI-MM pass-through interface 42
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_42_AWADDR,
    input wire [7:0]                      AP_AXIMM_42_AWLEN,
    input wire [2:0]                      AP_AXIMM_42_AWSIZE,
    input wire [1:0]                      AP_AXIMM_42_AWBURST,
    input wire [1:0]                      AP_AXIMM_42_AWLOCK,
    input wire [3:0]                      AP_AXIMM_42_AWCACHE,
    input wire [2:0]                      AP_AXIMM_42_AWPROT,
    input wire [3:0]                      AP_AXIMM_42_AWREGION,
    input wire [3:0]                      AP_AXIMM_42_AWQOS,
    input wire                            AP_AXIMM_42_AWVALID,
    output  wire                            AP_AXIMM_42_AWREADY,
    input wire [M_AXIMM_42_DATA_WIDTH-1:0]   AP_AXIMM_42_WDATA,
    input wire [M_AXIMM_42_DATA_WIDTH/8-1:0] AP_AXIMM_42_WSTRB,
    input wire                            AP_AXIMM_42_WLAST,
    input wire                            AP_AXIMM_42_WVALID,
    output  wire                            AP_AXIMM_42_WREADY,
    output  wire [1:0]                      AP_AXIMM_42_BRESP,
    output  wire                            AP_AXIMM_42_BVALID,
    input wire                            AP_AXIMM_42_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_42_ARADDR,
    input wire [7:0]                      AP_AXIMM_42_ARLEN,
    input wire [2:0]                      AP_AXIMM_42_ARSIZE,
    input wire [1:0]                      AP_AXIMM_42_ARBURST,
    input wire [1:0]                      AP_AXIMM_42_ARLOCK,
    input wire [3:0]                      AP_AXIMM_42_ARCACHE,
    input wire [2:0]                      AP_AXIMM_42_ARPROT,
    input wire [3:0]                      AP_AXIMM_42_ARREGION,
    input wire [3:0]                      AP_AXIMM_42_ARQOS,
    input wire                            AP_AXIMM_42_ARVALID,
    output  wire                            AP_AXIMM_42_ARREADY,
    output  wire [M_AXIMM_42_DATA_WIDTH-1:0]   AP_AXIMM_42_RDATA,
    output  wire [1:0]                      AP_AXIMM_42_RRESP,
    output  wire                            AP_AXIMM_42_RLAST,
    output  wire                            AP_AXIMM_42_RVALID,
    input  wire                            AP_AXIMM_42_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_42_AWADDR,
    output wire [7:0]                      M_AXIMM_42_AWLEN,
    output wire [2:0]                      M_AXIMM_42_AWSIZE,
    output wire [1:0]                      M_AXIMM_42_AWBURST,
    output wire [1:0]                      M_AXIMM_42_AWLOCK,
    output wire [3:0]                      M_AXIMM_42_AWCACHE,
    output wire [2:0]                      M_AXIMM_42_AWPROT,
    output wire [3:0]                      M_AXIMM_42_AWREGION,
    output wire [3:0]                      M_AXIMM_42_AWQOS,
    output wire                            M_AXIMM_42_AWVALID,
    input  wire                            M_AXIMM_42_AWREADY,
    output wire [M_AXIMM_42_DATA_WIDTH-1:0]   M_AXIMM_42_WDATA,
    output wire [M_AXIMM_42_DATA_WIDTH/8-1:0] M_AXIMM_42_WSTRB,
    output wire                            M_AXIMM_42_WLAST,
    output wire                            M_AXIMM_42_WVALID,
    input  wire                            M_AXIMM_42_WREADY,
    input  wire [1:0]                      M_AXIMM_42_BRESP,
    input  wire                            M_AXIMM_42_BVALID,
    output wire                            M_AXIMM_42_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_42_ARADDR,
    output wire [7:0]                      M_AXIMM_42_ARLEN,
    output wire [2:0]                      M_AXIMM_42_ARSIZE,
    output wire [1:0]                      M_AXIMM_42_ARBURST,
    output wire [1:0]                      M_AXIMM_42_ARLOCK,
    output wire [3:0]                      M_AXIMM_42_ARCACHE,
    output wire [2:0]                      M_AXIMM_42_ARPROT,
    output wire [3:0]                      M_AXIMM_42_ARREGION,
    output wire [3:0]                      M_AXIMM_42_ARQOS,
    output wire                            M_AXIMM_42_ARVALID,
    input  wire                            M_AXIMM_42_ARREADY,
    input  wire [M_AXIMM_42_DATA_WIDTH-1:0]   M_AXIMM_42_RDATA,
    input  wire [1:0]                      M_AXIMM_42_RRESP,
    input  wire                            M_AXIMM_42_RLAST,
    input  wire                            M_AXIMM_42_RVALID,
    output wire                            M_AXIMM_42_RREADY,
    //AXI-MM pass-through interface 43
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_43_AWADDR,
    input wire [7:0]                      AP_AXIMM_43_AWLEN,
    input wire [2:0]                      AP_AXIMM_43_AWSIZE,
    input wire [1:0]                      AP_AXIMM_43_AWBURST,
    input wire [1:0]                      AP_AXIMM_43_AWLOCK,
    input wire [3:0]                      AP_AXIMM_43_AWCACHE,
    input wire [2:0]                      AP_AXIMM_43_AWPROT,
    input wire [3:0]                      AP_AXIMM_43_AWREGION,
    input wire [3:0]                      AP_AXIMM_43_AWQOS,
    input wire                            AP_AXIMM_43_AWVALID,
    output  wire                            AP_AXIMM_43_AWREADY,
    input wire [M_AXIMM_43_DATA_WIDTH-1:0]   AP_AXIMM_43_WDATA,
    input wire [M_AXIMM_43_DATA_WIDTH/8-1:0] AP_AXIMM_43_WSTRB,
    input wire                            AP_AXIMM_43_WLAST,
    input wire                            AP_AXIMM_43_WVALID,
    output  wire                            AP_AXIMM_43_WREADY,
    output  wire [1:0]                      AP_AXIMM_43_BRESP,
    output  wire                            AP_AXIMM_43_BVALID,
    input wire                            AP_AXIMM_43_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_43_ARADDR,
    input wire [7:0]                      AP_AXIMM_43_ARLEN,
    input wire [2:0]                      AP_AXIMM_43_ARSIZE,
    input wire [1:0]                      AP_AXIMM_43_ARBURST,
    input wire [1:0]                      AP_AXIMM_43_ARLOCK,
    input wire [3:0]                      AP_AXIMM_43_ARCACHE,
    input wire [2:0]                      AP_AXIMM_43_ARPROT,
    input wire [3:0]                      AP_AXIMM_43_ARREGION,
    input wire [3:0]                      AP_AXIMM_43_ARQOS,
    input wire                            AP_AXIMM_43_ARVALID,
    output  wire                            AP_AXIMM_43_ARREADY,
    output  wire [M_AXIMM_43_DATA_WIDTH-1:0]   AP_AXIMM_43_RDATA,
    output  wire [1:0]                      AP_AXIMM_43_RRESP,
    output  wire                            AP_AXIMM_43_RLAST,
    output  wire                            AP_AXIMM_43_RVALID,
    input  wire                            AP_AXIMM_43_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_43_AWADDR,
    output wire [7:0]                      M_AXIMM_43_AWLEN,
    output wire [2:0]                      M_AXIMM_43_AWSIZE,
    output wire [1:0]                      M_AXIMM_43_AWBURST,
    output wire [1:0]                      M_AXIMM_43_AWLOCK,
    output wire [3:0]                      M_AXIMM_43_AWCACHE,
    output wire [2:0]                      M_AXIMM_43_AWPROT,
    output wire [3:0]                      M_AXIMM_43_AWREGION,
    output wire [3:0]                      M_AXIMM_43_AWQOS,
    output wire                            M_AXIMM_43_AWVALID,
    input  wire                            M_AXIMM_43_AWREADY,
    output wire [M_AXIMM_43_DATA_WIDTH-1:0]   M_AXIMM_43_WDATA,
    output wire [M_AXIMM_43_DATA_WIDTH/8-1:0] M_AXIMM_43_WSTRB,
    output wire                            M_AXIMM_43_WLAST,
    output wire                            M_AXIMM_43_WVALID,
    input  wire                            M_AXIMM_43_WREADY,
    input  wire [1:0]                      M_AXIMM_43_BRESP,
    input  wire                            M_AXIMM_43_BVALID,
    output wire                            M_AXIMM_43_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_43_ARADDR,
    output wire [7:0]                      M_AXIMM_43_ARLEN,
    output wire [2:0]                      M_AXIMM_43_ARSIZE,
    output wire [1:0]                      M_AXIMM_43_ARBURST,
    output wire [1:0]                      M_AXIMM_43_ARLOCK,
    output wire [3:0]                      M_AXIMM_43_ARCACHE,
    output wire [2:0]                      M_AXIMM_43_ARPROT,
    output wire [3:0]                      M_AXIMM_43_ARREGION,
    output wire [3:0]                      M_AXIMM_43_ARQOS,
    output wire                            M_AXIMM_43_ARVALID,
    input  wire                            M_AXIMM_43_ARREADY,
    input  wire [M_AXIMM_43_DATA_WIDTH-1:0]   M_AXIMM_43_RDATA,
    input  wire [1:0]                      M_AXIMM_43_RRESP,
    input  wire                            M_AXIMM_43_RLAST,
    input  wire                            M_AXIMM_43_RVALID,
    output wire                            M_AXIMM_43_RREADY,
    //AXI-MM pass-through interface 44
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_44_AWADDR,
    input wire [7:0]                      AP_AXIMM_44_AWLEN,
    input wire [2:0]                      AP_AXIMM_44_AWSIZE,
    input wire [1:0]                      AP_AXIMM_44_AWBURST,
    input wire [1:0]                      AP_AXIMM_44_AWLOCK,
    input wire [3:0]                      AP_AXIMM_44_AWCACHE,
    input wire [2:0]                      AP_AXIMM_44_AWPROT,
    input wire [3:0]                      AP_AXIMM_44_AWREGION,
    input wire [3:0]                      AP_AXIMM_44_AWQOS,
    input wire                            AP_AXIMM_44_AWVALID,
    output  wire                            AP_AXIMM_44_AWREADY,
    input wire [M_AXIMM_44_DATA_WIDTH-1:0]   AP_AXIMM_44_WDATA,
    input wire [M_AXIMM_44_DATA_WIDTH/8-1:0] AP_AXIMM_44_WSTRB,
    input wire                            AP_AXIMM_44_WLAST,
    input wire                            AP_AXIMM_44_WVALID,
    output  wire                            AP_AXIMM_44_WREADY,
    output  wire [1:0]                      AP_AXIMM_44_BRESP,
    output  wire                            AP_AXIMM_44_BVALID,
    input wire                            AP_AXIMM_44_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_44_ARADDR,
    input wire [7:0]                      AP_AXIMM_44_ARLEN,
    input wire [2:0]                      AP_AXIMM_44_ARSIZE,
    input wire [1:0]                      AP_AXIMM_44_ARBURST,
    input wire [1:0]                      AP_AXIMM_44_ARLOCK,
    input wire [3:0]                      AP_AXIMM_44_ARCACHE,
    input wire [2:0]                      AP_AXIMM_44_ARPROT,
    input wire [3:0]                      AP_AXIMM_44_ARREGION,
    input wire [3:0]                      AP_AXIMM_44_ARQOS,
    input wire                            AP_AXIMM_44_ARVALID,
    output  wire                            AP_AXIMM_44_ARREADY,
    output  wire [M_AXIMM_44_DATA_WIDTH-1:0]   AP_AXIMM_44_RDATA,
    output  wire [1:0]                      AP_AXIMM_44_RRESP,
    output  wire                            AP_AXIMM_44_RLAST,
    output  wire                            AP_AXIMM_44_RVALID,
    input  wire                            AP_AXIMM_44_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_44_AWADDR,
    output wire [7:0]                      M_AXIMM_44_AWLEN,
    output wire [2:0]                      M_AXIMM_44_AWSIZE,
    output wire [1:0]                      M_AXIMM_44_AWBURST,
    output wire [1:0]                      M_AXIMM_44_AWLOCK,
    output wire [3:0]                      M_AXIMM_44_AWCACHE,
    output wire [2:0]                      M_AXIMM_44_AWPROT,
    output wire [3:0]                      M_AXIMM_44_AWREGION,
    output wire [3:0]                      M_AXIMM_44_AWQOS,
    output wire                            M_AXIMM_44_AWVALID,
    input  wire                            M_AXIMM_44_AWREADY,
    output wire [M_AXIMM_44_DATA_WIDTH-1:0]   M_AXIMM_44_WDATA,
    output wire [M_AXIMM_44_DATA_WIDTH/8-1:0] M_AXIMM_44_WSTRB,
    output wire                            M_AXIMM_44_WLAST,
    output wire                            M_AXIMM_44_WVALID,
    input  wire                            M_AXIMM_44_WREADY,
    input  wire [1:0]                      M_AXIMM_44_BRESP,
    input  wire                            M_AXIMM_44_BVALID,
    output wire                            M_AXIMM_44_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_44_ARADDR,
    output wire [7:0]                      M_AXIMM_44_ARLEN,
    output wire [2:0]                      M_AXIMM_44_ARSIZE,
    output wire [1:0]                      M_AXIMM_44_ARBURST,
    output wire [1:0]                      M_AXIMM_44_ARLOCK,
    output wire [3:0]                      M_AXIMM_44_ARCACHE,
    output wire [2:0]                      M_AXIMM_44_ARPROT,
    output wire [3:0]                      M_AXIMM_44_ARREGION,
    output wire [3:0]                      M_AXIMM_44_ARQOS,
    output wire                            M_AXIMM_44_ARVALID,
    input  wire                            M_AXIMM_44_ARREADY,
    input  wire [M_AXIMM_44_DATA_WIDTH-1:0]   M_AXIMM_44_RDATA,
    input  wire [1:0]                      M_AXIMM_44_RRESP,
    input  wire                            M_AXIMM_44_RLAST,
    input  wire                            M_AXIMM_44_RVALID,
    output wire                            M_AXIMM_44_RREADY,
    //AXI-MM pass-through interface 45
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_45_AWADDR,
    input wire [7:0]                      AP_AXIMM_45_AWLEN,
    input wire [2:0]                      AP_AXIMM_45_AWSIZE,
    input wire [1:0]                      AP_AXIMM_45_AWBURST,
    input wire [1:0]                      AP_AXIMM_45_AWLOCK,
    input wire [3:0]                      AP_AXIMM_45_AWCACHE,
    input wire [2:0]                      AP_AXIMM_45_AWPROT,
    input wire [3:0]                      AP_AXIMM_45_AWREGION,
    input wire [3:0]                      AP_AXIMM_45_AWQOS,
    input wire                            AP_AXIMM_45_AWVALID,
    output  wire                            AP_AXIMM_45_AWREADY,
    input wire [M_AXIMM_45_DATA_WIDTH-1:0]   AP_AXIMM_45_WDATA,
    input wire [M_AXIMM_45_DATA_WIDTH/8-1:0] AP_AXIMM_45_WSTRB,
    input wire                            AP_AXIMM_45_WLAST,
    input wire                            AP_AXIMM_45_WVALID,
    output  wire                            AP_AXIMM_45_WREADY,
    output  wire [1:0]                      AP_AXIMM_45_BRESP,
    output  wire                            AP_AXIMM_45_BVALID,
    input wire                            AP_AXIMM_45_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_45_ARADDR,
    input wire [7:0]                      AP_AXIMM_45_ARLEN,
    input wire [2:0]                      AP_AXIMM_45_ARSIZE,
    input wire [1:0]                      AP_AXIMM_45_ARBURST,
    input wire [1:0]                      AP_AXIMM_45_ARLOCK,
    input wire [3:0]                      AP_AXIMM_45_ARCACHE,
    input wire [2:0]                      AP_AXIMM_45_ARPROT,
    input wire [3:0]                      AP_AXIMM_45_ARREGION,
    input wire [3:0]                      AP_AXIMM_45_ARQOS,
    input wire                            AP_AXIMM_45_ARVALID,
    output  wire                            AP_AXIMM_45_ARREADY,
    output  wire [M_AXIMM_45_DATA_WIDTH-1:0]   AP_AXIMM_45_RDATA,
    output  wire [1:0]                      AP_AXIMM_45_RRESP,
    output  wire                            AP_AXIMM_45_RLAST,
    output  wire                            AP_AXIMM_45_RVALID,
    input  wire                            AP_AXIMM_45_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_45_AWADDR,
    output wire [7:0]                      M_AXIMM_45_AWLEN,
    output wire [2:0]                      M_AXIMM_45_AWSIZE,
    output wire [1:0]                      M_AXIMM_45_AWBURST,
    output wire [1:0]                      M_AXIMM_45_AWLOCK,
    output wire [3:0]                      M_AXIMM_45_AWCACHE,
    output wire [2:0]                      M_AXIMM_45_AWPROT,
    output wire [3:0]                      M_AXIMM_45_AWREGION,
    output wire [3:0]                      M_AXIMM_45_AWQOS,
    output wire                            M_AXIMM_45_AWVALID,
    input  wire                            M_AXIMM_45_AWREADY,
    output wire [M_AXIMM_45_DATA_WIDTH-1:0]   M_AXIMM_45_WDATA,
    output wire [M_AXIMM_45_DATA_WIDTH/8-1:0] M_AXIMM_45_WSTRB,
    output wire                            M_AXIMM_45_WLAST,
    output wire                            M_AXIMM_45_WVALID,
    input  wire                            M_AXIMM_45_WREADY,
    input  wire [1:0]                      M_AXIMM_45_BRESP,
    input  wire                            M_AXIMM_45_BVALID,
    output wire                            M_AXIMM_45_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_45_ARADDR,
    output wire [7:0]                      M_AXIMM_45_ARLEN,
    output wire [2:0]                      M_AXIMM_45_ARSIZE,
    output wire [1:0]                      M_AXIMM_45_ARBURST,
    output wire [1:0]                      M_AXIMM_45_ARLOCK,
    output wire [3:0]                      M_AXIMM_45_ARCACHE,
    output wire [2:0]                      M_AXIMM_45_ARPROT,
    output wire [3:0]                      M_AXIMM_45_ARREGION,
    output wire [3:0]                      M_AXIMM_45_ARQOS,
    output wire                            M_AXIMM_45_ARVALID,
    input  wire                            M_AXIMM_45_ARREADY,
    input  wire [M_AXIMM_45_DATA_WIDTH-1:0]   M_AXIMM_45_RDATA,
    input  wire [1:0]                      M_AXIMM_45_RRESP,
    input  wire                            M_AXIMM_45_RLAST,
    input  wire                            M_AXIMM_45_RVALID,
    output wire                            M_AXIMM_45_RREADY,
    //AXI-MM pass-through interface 46
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_46_AWADDR,
    input wire [7:0]                      AP_AXIMM_46_AWLEN,
    input wire [2:0]                      AP_AXIMM_46_AWSIZE,
    input wire [1:0]                      AP_AXIMM_46_AWBURST,
    input wire [1:0]                      AP_AXIMM_46_AWLOCK,
    input wire [3:0]                      AP_AXIMM_46_AWCACHE,
    input wire [2:0]                      AP_AXIMM_46_AWPROT,
    input wire [3:0]                      AP_AXIMM_46_AWREGION,
    input wire [3:0]                      AP_AXIMM_46_AWQOS,
    input wire                            AP_AXIMM_46_AWVALID,
    output  wire                            AP_AXIMM_46_AWREADY,
    input wire [M_AXIMM_46_DATA_WIDTH-1:0]   AP_AXIMM_46_WDATA,
    input wire [M_AXIMM_46_DATA_WIDTH/8-1:0] AP_AXIMM_46_WSTRB,
    input wire                            AP_AXIMM_46_WLAST,
    input wire                            AP_AXIMM_46_WVALID,
    output  wire                            AP_AXIMM_46_WREADY,
    output  wire [1:0]                      AP_AXIMM_46_BRESP,
    output  wire                            AP_AXIMM_46_BVALID,
    input wire                            AP_AXIMM_46_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_46_ARADDR,
    input wire [7:0]                      AP_AXIMM_46_ARLEN,
    input wire [2:0]                      AP_AXIMM_46_ARSIZE,
    input wire [1:0]                      AP_AXIMM_46_ARBURST,
    input wire [1:0]                      AP_AXIMM_46_ARLOCK,
    input wire [3:0]                      AP_AXIMM_46_ARCACHE,
    input wire [2:0]                      AP_AXIMM_46_ARPROT,
    input wire [3:0]                      AP_AXIMM_46_ARREGION,
    input wire [3:0]                      AP_AXIMM_46_ARQOS,
    input wire                            AP_AXIMM_46_ARVALID,
    output  wire                            AP_AXIMM_46_ARREADY,
    output  wire [M_AXIMM_46_DATA_WIDTH-1:0]   AP_AXIMM_46_RDATA,
    output  wire [1:0]                      AP_AXIMM_46_RRESP,
    output  wire                            AP_AXIMM_46_RLAST,
    output  wire                            AP_AXIMM_46_RVALID,
    input  wire                            AP_AXIMM_46_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_46_AWADDR,
    output wire [7:0]                      M_AXIMM_46_AWLEN,
    output wire [2:0]                      M_AXIMM_46_AWSIZE,
    output wire [1:0]                      M_AXIMM_46_AWBURST,
    output wire [1:0]                      M_AXIMM_46_AWLOCK,
    output wire [3:0]                      M_AXIMM_46_AWCACHE,
    output wire [2:0]                      M_AXIMM_46_AWPROT,
    output wire [3:0]                      M_AXIMM_46_AWREGION,
    output wire [3:0]                      M_AXIMM_46_AWQOS,
    output wire                            M_AXIMM_46_AWVALID,
    input  wire                            M_AXIMM_46_AWREADY,
    output wire [M_AXIMM_46_DATA_WIDTH-1:0]   M_AXIMM_46_WDATA,
    output wire [M_AXIMM_46_DATA_WIDTH/8-1:0] M_AXIMM_46_WSTRB,
    output wire                            M_AXIMM_46_WLAST,
    output wire                            M_AXIMM_46_WVALID,
    input  wire                            M_AXIMM_46_WREADY,
    input  wire [1:0]                      M_AXIMM_46_BRESP,
    input  wire                            M_AXIMM_46_BVALID,
    output wire                            M_AXIMM_46_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_46_ARADDR,
    output wire [7:0]                      M_AXIMM_46_ARLEN,
    output wire [2:0]                      M_AXIMM_46_ARSIZE,
    output wire [1:0]                      M_AXIMM_46_ARBURST,
    output wire [1:0]                      M_AXIMM_46_ARLOCK,
    output wire [3:0]                      M_AXIMM_46_ARCACHE,
    output wire [2:0]                      M_AXIMM_46_ARPROT,
    output wire [3:0]                      M_AXIMM_46_ARREGION,
    output wire [3:0]                      M_AXIMM_46_ARQOS,
    output wire                            M_AXIMM_46_ARVALID,
    input  wire                            M_AXIMM_46_ARREADY,
    input  wire [M_AXIMM_46_DATA_WIDTH-1:0]   M_AXIMM_46_RDATA,
    input  wire [1:0]                      M_AXIMM_46_RRESP,
    input  wire                            M_AXIMM_46_RLAST,
    input  wire                            M_AXIMM_46_RVALID,
    output wire                            M_AXIMM_46_RREADY,
    //AXI-MM pass-through interface 47
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_47_AWADDR,
    input wire [7:0]                      AP_AXIMM_47_AWLEN,
    input wire [2:0]                      AP_AXIMM_47_AWSIZE,
    input wire [1:0]                      AP_AXIMM_47_AWBURST,
    input wire [1:0]                      AP_AXIMM_47_AWLOCK,
    input wire [3:0]                      AP_AXIMM_47_AWCACHE,
    input wire [2:0]                      AP_AXIMM_47_AWPROT,
    input wire [3:0]                      AP_AXIMM_47_AWREGION,
    input wire [3:0]                      AP_AXIMM_47_AWQOS,
    input wire                            AP_AXIMM_47_AWVALID,
    output  wire                            AP_AXIMM_47_AWREADY,
    input wire [M_AXIMM_47_DATA_WIDTH-1:0]   AP_AXIMM_47_WDATA,
    input wire [M_AXIMM_47_DATA_WIDTH/8-1:0] AP_AXIMM_47_WSTRB,
    input wire                            AP_AXIMM_47_WLAST,
    input wire                            AP_AXIMM_47_WVALID,
    output  wire                            AP_AXIMM_47_WREADY,
    output  wire [1:0]                      AP_AXIMM_47_BRESP,
    output  wire                            AP_AXIMM_47_BVALID,
    input wire                            AP_AXIMM_47_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_47_ARADDR,
    input wire [7:0]                      AP_AXIMM_47_ARLEN,
    input wire [2:0]                      AP_AXIMM_47_ARSIZE,
    input wire [1:0]                      AP_AXIMM_47_ARBURST,
    input wire [1:0]                      AP_AXIMM_47_ARLOCK,
    input wire [3:0]                      AP_AXIMM_47_ARCACHE,
    input wire [2:0]                      AP_AXIMM_47_ARPROT,
    input wire [3:0]                      AP_AXIMM_47_ARREGION,
    input wire [3:0]                      AP_AXIMM_47_ARQOS,
    input wire                            AP_AXIMM_47_ARVALID,
    output  wire                            AP_AXIMM_47_ARREADY,
    output  wire [M_AXIMM_47_DATA_WIDTH-1:0]   AP_AXIMM_47_RDATA,
    output  wire [1:0]                      AP_AXIMM_47_RRESP,
    output  wire                            AP_AXIMM_47_RLAST,
    output  wire                            AP_AXIMM_47_RVALID,
    input  wire                            AP_AXIMM_47_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_47_AWADDR,
    output wire [7:0]                      M_AXIMM_47_AWLEN,
    output wire [2:0]                      M_AXIMM_47_AWSIZE,
    output wire [1:0]                      M_AXIMM_47_AWBURST,
    output wire [1:0]                      M_AXIMM_47_AWLOCK,
    output wire [3:0]                      M_AXIMM_47_AWCACHE,
    output wire [2:0]                      M_AXIMM_47_AWPROT,
    output wire [3:0]                      M_AXIMM_47_AWREGION,
    output wire [3:0]                      M_AXIMM_47_AWQOS,
    output wire                            M_AXIMM_47_AWVALID,
    input  wire                            M_AXIMM_47_AWREADY,
    output wire [M_AXIMM_47_DATA_WIDTH-1:0]   M_AXIMM_47_WDATA,
    output wire [M_AXIMM_47_DATA_WIDTH/8-1:0] M_AXIMM_47_WSTRB,
    output wire                            M_AXIMM_47_WLAST,
    output wire                            M_AXIMM_47_WVALID,
    input  wire                            M_AXIMM_47_WREADY,
    input  wire [1:0]                      M_AXIMM_47_BRESP,
    input  wire                            M_AXIMM_47_BVALID,
    output wire                            M_AXIMM_47_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_47_ARADDR,
    output wire [7:0]                      M_AXIMM_47_ARLEN,
    output wire [2:0]                      M_AXIMM_47_ARSIZE,
    output wire [1:0]                      M_AXIMM_47_ARBURST,
    output wire [1:0]                      M_AXIMM_47_ARLOCK,
    output wire [3:0]                      M_AXIMM_47_ARCACHE,
    output wire [2:0]                      M_AXIMM_47_ARPROT,
    output wire [3:0]                      M_AXIMM_47_ARREGION,
    output wire [3:0]                      M_AXIMM_47_ARQOS,
    output wire                            M_AXIMM_47_ARVALID,
    input  wire                            M_AXIMM_47_ARREADY,
    input  wire [M_AXIMM_47_DATA_WIDTH-1:0]   M_AXIMM_47_RDATA,
    input  wire [1:0]                      M_AXIMM_47_RRESP,
    input  wire                            M_AXIMM_47_RLAST,
    input  wire                            M_AXIMM_47_RVALID,
    output wire                            M_AXIMM_47_RREADY,
    //AXI-MM pass-through interface 48
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_48_AWADDR,
    input wire [7:0]                      AP_AXIMM_48_AWLEN,
    input wire [2:0]                      AP_AXIMM_48_AWSIZE,
    input wire [1:0]                      AP_AXIMM_48_AWBURST,
    input wire [1:0]                      AP_AXIMM_48_AWLOCK,
    input wire [3:0]                      AP_AXIMM_48_AWCACHE,
    input wire [2:0]                      AP_AXIMM_48_AWPROT,
    input wire [3:0]                      AP_AXIMM_48_AWREGION,
    input wire [3:0]                      AP_AXIMM_48_AWQOS,
    input wire                            AP_AXIMM_48_AWVALID,
    output  wire                            AP_AXIMM_48_AWREADY,
    input wire [M_AXIMM_48_DATA_WIDTH-1:0]   AP_AXIMM_48_WDATA,
    input wire [M_AXIMM_48_DATA_WIDTH/8-1:0] AP_AXIMM_48_WSTRB,
    input wire                            AP_AXIMM_48_WLAST,
    input wire                            AP_AXIMM_48_WVALID,
    output  wire                            AP_AXIMM_48_WREADY,
    output  wire [1:0]                      AP_AXIMM_48_BRESP,
    output  wire                            AP_AXIMM_48_BVALID,
    input wire                            AP_AXIMM_48_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_48_ARADDR,
    input wire [7:0]                      AP_AXIMM_48_ARLEN,
    input wire [2:0]                      AP_AXIMM_48_ARSIZE,
    input wire [1:0]                      AP_AXIMM_48_ARBURST,
    input wire [1:0]                      AP_AXIMM_48_ARLOCK,
    input wire [3:0]                      AP_AXIMM_48_ARCACHE,
    input wire [2:0]                      AP_AXIMM_48_ARPROT,
    input wire [3:0]                      AP_AXIMM_48_ARREGION,
    input wire [3:0]                      AP_AXIMM_48_ARQOS,
    input wire                            AP_AXIMM_48_ARVALID,
    output  wire                            AP_AXIMM_48_ARREADY,
    output  wire [M_AXIMM_48_DATA_WIDTH-1:0]   AP_AXIMM_48_RDATA,
    output  wire [1:0]                      AP_AXIMM_48_RRESP,
    output  wire                            AP_AXIMM_48_RLAST,
    output  wire                            AP_AXIMM_48_RVALID,
    input  wire                            AP_AXIMM_48_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_48_AWADDR,
    output wire [7:0]                      M_AXIMM_48_AWLEN,
    output wire [2:0]                      M_AXIMM_48_AWSIZE,
    output wire [1:0]                      M_AXIMM_48_AWBURST,
    output wire [1:0]                      M_AXIMM_48_AWLOCK,
    output wire [3:0]                      M_AXIMM_48_AWCACHE,
    output wire [2:0]                      M_AXIMM_48_AWPROT,
    output wire [3:0]                      M_AXIMM_48_AWREGION,
    output wire [3:0]                      M_AXIMM_48_AWQOS,
    output wire                            M_AXIMM_48_AWVALID,
    input  wire                            M_AXIMM_48_AWREADY,
    output wire [M_AXIMM_48_DATA_WIDTH-1:0]   M_AXIMM_48_WDATA,
    output wire [M_AXIMM_48_DATA_WIDTH/8-1:0] M_AXIMM_48_WSTRB,
    output wire                            M_AXIMM_48_WLAST,
    output wire                            M_AXIMM_48_WVALID,
    input  wire                            M_AXIMM_48_WREADY,
    input  wire [1:0]                      M_AXIMM_48_BRESP,
    input  wire                            M_AXIMM_48_BVALID,
    output wire                            M_AXIMM_48_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_48_ARADDR,
    output wire [7:0]                      M_AXIMM_48_ARLEN,
    output wire [2:0]                      M_AXIMM_48_ARSIZE,
    output wire [1:0]                      M_AXIMM_48_ARBURST,
    output wire [1:0]                      M_AXIMM_48_ARLOCK,
    output wire [3:0]                      M_AXIMM_48_ARCACHE,
    output wire [2:0]                      M_AXIMM_48_ARPROT,
    output wire [3:0]                      M_AXIMM_48_ARREGION,
    output wire [3:0]                      M_AXIMM_48_ARQOS,
    output wire                            M_AXIMM_48_ARVALID,
    input  wire                            M_AXIMM_48_ARREADY,
    input  wire [M_AXIMM_48_DATA_WIDTH-1:0]   M_AXIMM_48_RDATA,
    input  wire [1:0]                      M_AXIMM_48_RRESP,
    input  wire                            M_AXIMM_48_RLAST,
    input  wire                            M_AXIMM_48_RVALID,
    output wire                            M_AXIMM_48_RREADY,
    //AXI-MM pass-through interface 49
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_49_AWADDR,
    input wire [7:0]                      AP_AXIMM_49_AWLEN,
    input wire [2:0]                      AP_AXIMM_49_AWSIZE,
    input wire [1:0]                      AP_AXIMM_49_AWBURST,
    input wire [1:0]                      AP_AXIMM_49_AWLOCK,
    input wire [3:0]                      AP_AXIMM_49_AWCACHE,
    input wire [2:0]                      AP_AXIMM_49_AWPROT,
    input wire [3:0]                      AP_AXIMM_49_AWREGION,
    input wire [3:0]                      AP_AXIMM_49_AWQOS,
    input wire                            AP_AXIMM_49_AWVALID,
    output  wire                            AP_AXIMM_49_AWREADY,
    input wire [M_AXIMM_49_DATA_WIDTH-1:0]   AP_AXIMM_49_WDATA,
    input wire [M_AXIMM_49_DATA_WIDTH/8-1:0] AP_AXIMM_49_WSTRB,
    input wire                            AP_AXIMM_49_WLAST,
    input wire                            AP_AXIMM_49_WVALID,
    output  wire                            AP_AXIMM_49_WREADY,
    output  wire [1:0]                      AP_AXIMM_49_BRESP,
    output  wire                            AP_AXIMM_49_BVALID,
    input wire                            AP_AXIMM_49_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_49_ARADDR,
    input wire [7:0]                      AP_AXIMM_49_ARLEN,
    input wire [2:0]                      AP_AXIMM_49_ARSIZE,
    input wire [1:0]                      AP_AXIMM_49_ARBURST,
    input wire [1:0]                      AP_AXIMM_49_ARLOCK,
    input wire [3:0]                      AP_AXIMM_49_ARCACHE,
    input wire [2:0]                      AP_AXIMM_49_ARPROT,
    input wire [3:0]                      AP_AXIMM_49_ARREGION,
    input wire [3:0]                      AP_AXIMM_49_ARQOS,
    input wire                            AP_AXIMM_49_ARVALID,
    output  wire                            AP_AXIMM_49_ARREADY,
    output  wire [M_AXIMM_49_DATA_WIDTH-1:0]   AP_AXIMM_49_RDATA,
    output  wire [1:0]                      AP_AXIMM_49_RRESP,
    output  wire                            AP_AXIMM_49_RLAST,
    output  wire                            AP_AXIMM_49_RVALID,
    input  wire                            AP_AXIMM_49_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_49_AWADDR,
    output wire [7:0]                      M_AXIMM_49_AWLEN,
    output wire [2:0]                      M_AXIMM_49_AWSIZE,
    output wire [1:0]                      M_AXIMM_49_AWBURST,
    output wire [1:0]                      M_AXIMM_49_AWLOCK,
    output wire [3:0]                      M_AXIMM_49_AWCACHE,
    output wire [2:0]                      M_AXIMM_49_AWPROT,
    output wire [3:0]                      M_AXIMM_49_AWREGION,
    output wire [3:0]                      M_AXIMM_49_AWQOS,
    output wire                            M_AXIMM_49_AWVALID,
    input  wire                            M_AXIMM_49_AWREADY,
    output wire [M_AXIMM_49_DATA_WIDTH-1:0]   M_AXIMM_49_WDATA,
    output wire [M_AXIMM_49_DATA_WIDTH/8-1:0] M_AXIMM_49_WSTRB,
    output wire                            M_AXIMM_49_WLAST,
    output wire                            M_AXIMM_49_WVALID,
    input  wire                            M_AXIMM_49_WREADY,
    input  wire [1:0]                      M_AXIMM_49_BRESP,
    input  wire                            M_AXIMM_49_BVALID,
    output wire                            M_AXIMM_49_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_49_ARADDR,
    output wire [7:0]                      M_AXIMM_49_ARLEN,
    output wire [2:0]                      M_AXIMM_49_ARSIZE,
    output wire [1:0]                      M_AXIMM_49_ARBURST,
    output wire [1:0]                      M_AXIMM_49_ARLOCK,
    output wire [3:0]                      M_AXIMM_49_ARCACHE,
    output wire [2:0]                      M_AXIMM_49_ARPROT,
    output wire [3:0]                      M_AXIMM_49_ARREGION,
    output wire [3:0]                      M_AXIMM_49_ARQOS,
    output wire                            M_AXIMM_49_ARVALID,
    input  wire                            M_AXIMM_49_ARREADY,
    input  wire [M_AXIMM_49_DATA_WIDTH-1:0]   M_AXIMM_49_RDATA,
    input  wire [1:0]                      M_AXIMM_49_RRESP,
    input  wire                            M_AXIMM_49_RLAST,
    input  wire                            M_AXIMM_49_RVALID,
    output wire                            M_AXIMM_49_RREADY,
    //AXI-MM pass-through interface 50
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_50_AWADDR,
    input wire [7:0]                      AP_AXIMM_50_AWLEN,
    input wire [2:0]                      AP_AXIMM_50_AWSIZE,
    input wire [1:0]                      AP_AXIMM_50_AWBURST,
    input wire [1:0]                      AP_AXIMM_50_AWLOCK,
    input wire [3:0]                      AP_AXIMM_50_AWCACHE,
    input wire [2:0]                      AP_AXIMM_50_AWPROT,
    input wire [3:0]                      AP_AXIMM_50_AWREGION,
    input wire [3:0]                      AP_AXIMM_50_AWQOS,
    input wire                            AP_AXIMM_50_AWVALID,
    output  wire                            AP_AXIMM_50_AWREADY,
    input wire [M_AXIMM_50_DATA_WIDTH-1:0]   AP_AXIMM_50_WDATA,
    input wire [M_AXIMM_50_DATA_WIDTH/8-1:0] AP_AXIMM_50_WSTRB,
    input wire                            AP_AXIMM_50_WLAST,
    input wire                            AP_AXIMM_50_WVALID,
    output  wire                            AP_AXIMM_50_WREADY,
    output  wire [1:0]                      AP_AXIMM_50_BRESP,
    output  wire                            AP_AXIMM_50_BVALID,
    input wire                            AP_AXIMM_50_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_50_ARADDR,
    input wire [7:0]                      AP_AXIMM_50_ARLEN,
    input wire [2:0]                      AP_AXIMM_50_ARSIZE,
    input wire [1:0]                      AP_AXIMM_50_ARBURST,
    input wire [1:0]                      AP_AXIMM_50_ARLOCK,
    input wire [3:0]                      AP_AXIMM_50_ARCACHE,
    input wire [2:0]                      AP_AXIMM_50_ARPROT,
    input wire [3:0]                      AP_AXIMM_50_ARREGION,
    input wire [3:0]                      AP_AXIMM_50_ARQOS,
    input wire                            AP_AXIMM_50_ARVALID,
    output  wire                            AP_AXIMM_50_ARREADY,
    output  wire [M_AXIMM_50_DATA_WIDTH-1:0]   AP_AXIMM_50_RDATA,
    output  wire [1:0]                      AP_AXIMM_50_RRESP,
    output  wire                            AP_AXIMM_50_RLAST,
    output  wire                            AP_AXIMM_50_RVALID,
    input  wire                            AP_AXIMM_50_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_50_AWADDR,
    output wire [7:0]                      M_AXIMM_50_AWLEN,
    output wire [2:0]                      M_AXIMM_50_AWSIZE,
    output wire [1:0]                      M_AXIMM_50_AWBURST,
    output wire [1:0]                      M_AXIMM_50_AWLOCK,
    output wire [3:0]                      M_AXIMM_50_AWCACHE,
    output wire [2:0]                      M_AXIMM_50_AWPROT,
    output wire [3:0]                      M_AXIMM_50_AWREGION,
    output wire [3:0]                      M_AXIMM_50_AWQOS,
    output wire                            M_AXIMM_50_AWVALID,
    input  wire                            M_AXIMM_50_AWREADY,
    output wire [M_AXIMM_50_DATA_WIDTH-1:0]   M_AXIMM_50_WDATA,
    output wire [M_AXIMM_50_DATA_WIDTH/8-1:0] M_AXIMM_50_WSTRB,
    output wire                            M_AXIMM_50_WLAST,
    output wire                            M_AXIMM_50_WVALID,
    input  wire                            M_AXIMM_50_WREADY,
    input  wire [1:0]                      M_AXIMM_50_BRESP,
    input  wire                            M_AXIMM_50_BVALID,
    output wire                            M_AXIMM_50_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_50_ARADDR,
    output wire [7:0]                      M_AXIMM_50_ARLEN,
    output wire [2:0]                      M_AXIMM_50_ARSIZE,
    output wire [1:0]                      M_AXIMM_50_ARBURST,
    output wire [1:0]                      M_AXIMM_50_ARLOCK,
    output wire [3:0]                      M_AXIMM_50_ARCACHE,
    output wire [2:0]                      M_AXIMM_50_ARPROT,
    output wire [3:0]                      M_AXIMM_50_ARREGION,
    output wire [3:0]                      M_AXIMM_50_ARQOS,
    output wire                            M_AXIMM_50_ARVALID,
    input  wire                            M_AXIMM_50_ARREADY,
    input  wire [M_AXIMM_50_DATA_WIDTH-1:0]   M_AXIMM_50_RDATA,
    input  wire [1:0]                      M_AXIMM_50_RRESP,
    input  wire                            M_AXIMM_50_RLAST,
    input  wire                            M_AXIMM_50_RVALID,
    output wire                            M_AXIMM_50_RREADY,
    //AXI-MM pass-through interface 51
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_51_AWADDR,
    input wire [7:0]                      AP_AXIMM_51_AWLEN,
    input wire [2:0]                      AP_AXIMM_51_AWSIZE,
    input wire [1:0]                      AP_AXIMM_51_AWBURST,
    input wire [1:0]                      AP_AXIMM_51_AWLOCK,
    input wire [3:0]                      AP_AXIMM_51_AWCACHE,
    input wire [2:0]                      AP_AXIMM_51_AWPROT,
    input wire [3:0]                      AP_AXIMM_51_AWREGION,
    input wire [3:0]                      AP_AXIMM_51_AWQOS,
    input wire                            AP_AXIMM_51_AWVALID,
    output  wire                            AP_AXIMM_51_AWREADY,
    input wire [M_AXIMM_51_DATA_WIDTH-1:0]   AP_AXIMM_51_WDATA,
    input wire [M_AXIMM_51_DATA_WIDTH/8-1:0] AP_AXIMM_51_WSTRB,
    input wire                            AP_AXIMM_51_WLAST,
    input wire                            AP_AXIMM_51_WVALID,
    output  wire                            AP_AXIMM_51_WREADY,
    output  wire [1:0]                      AP_AXIMM_51_BRESP,
    output  wire                            AP_AXIMM_51_BVALID,
    input wire                            AP_AXIMM_51_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_51_ARADDR,
    input wire [7:0]                      AP_AXIMM_51_ARLEN,
    input wire [2:0]                      AP_AXIMM_51_ARSIZE,
    input wire [1:0]                      AP_AXIMM_51_ARBURST,
    input wire [1:0]                      AP_AXIMM_51_ARLOCK,
    input wire [3:0]                      AP_AXIMM_51_ARCACHE,
    input wire [2:0]                      AP_AXIMM_51_ARPROT,
    input wire [3:0]                      AP_AXIMM_51_ARREGION,
    input wire [3:0]                      AP_AXIMM_51_ARQOS,
    input wire                            AP_AXIMM_51_ARVALID,
    output  wire                            AP_AXIMM_51_ARREADY,
    output  wire [M_AXIMM_51_DATA_WIDTH-1:0]   AP_AXIMM_51_RDATA,
    output  wire [1:0]                      AP_AXIMM_51_RRESP,
    output  wire                            AP_AXIMM_51_RLAST,
    output  wire                            AP_AXIMM_51_RVALID,
    input  wire                            AP_AXIMM_51_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_51_AWADDR,
    output wire [7:0]                      M_AXIMM_51_AWLEN,
    output wire [2:0]                      M_AXIMM_51_AWSIZE,
    output wire [1:0]                      M_AXIMM_51_AWBURST,
    output wire [1:0]                      M_AXIMM_51_AWLOCK,
    output wire [3:0]                      M_AXIMM_51_AWCACHE,
    output wire [2:0]                      M_AXIMM_51_AWPROT,
    output wire [3:0]                      M_AXIMM_51_AWREGION,
    output wire [3:0]                      M_AXIMM_51_AWQOS,
    output wire                            M_AXIMM_51_AWVALID,
    input  wire                            M_AXIMM_51_AWREADY,
    output wire [M_AXIMM_51_DATA_WIDTH-1:0]   M_AXIMM_51_WDATA,
    output wire [M_AXIMM_51_DATA_WIDTH/8-1:0] M_AXIMM_51_WSTRB,
    output wire                            M_AXIMM_51_WLAST,
    output wire                            M_AXIMM_51_WVALID,
    input  wire                            M_AXIMM_51_WREADY,
    input  wire [1:0]                      M_AXIMM_51_BRESP,
    input  wire                            M_AXIMM_51_BVALID,
    output wire                            M_AXIMM_51_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_51_ARADDR,
    output wire [7:0]                      M_AXIMM_51_ARLEN,
    output wire [2:0]                      M_AXIMM_51_ARSIZE,
    output wire [1:0]                      M_AXIMM_51_ARBURST,
    output wire [1:0]                      M_AXIMM_51_ARLOCK,
    output wire [3:0]                      M_AXIMM_51_ARCACHE,
    output wire [2:0]                      M_AXIMM_51_ARPROT,
    output wire [3:0]                      M_AXIMM_51_ARREGION,
    output wire [3:0]                      M_AXIMM_51_ARQOS,
    output wire                            M_AXIMM_51_ARVALID,
    input  wire                            M_AXIMM_51_ARREADY,
    input  wire [M_AXIMM_51_DATA_WIDTH-1:0]   M_AXIMM_51_RDATA,
    input  wire [1:0]                      M_AXIMM_51_RRESP,
    input  wire                            M_AXIMM_51_RLAST,
    input  wire                            M_AXIMM_51_RVALID,
    output wire                            M_AXIMM_51_RREADY,
    //AXI-MM pass-through interface 52
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_52_AWADDR,
    input wire [7:0]                      AP_AXIMM_52_AWLEN,
    input wire [2:0]                      AP_AXIMM_52_AWSIZE,
    input wire [1:0]                      AP_AXIMM_52_AWBURST,
    input wire [1:0]                      AP_AXIMM_52_AWLOCK,
    input wire [3:0]                      AP_AXIMM_52_AWCACHE,
    input wire [2:0]                      AP_AXIMM_52_AWPROT,
    input wire [3:0]                      AP_AXIMM_52_AWREGION,
    input wire [3:0]                      AP_AXIMM_52_AWQOS,
    input wire                            AP_AXIMM_52_AWVALID,
    output  wire                            AP_AXIMM_52_AWREADY,
    input wire [M_AXIMM_52_DATA_WIDTH-1:0]   AP_AXIMM_52_WDATA,
    input wire [M_AXIMM_52_DATA_WIDTH/8-1:0] AP_AXIMM_52_WSTRB,
    input wire                            AP_AXIMM_52_WLAST,
    input wire                            AP_AXIMM_52_WVALID,
    output  wire                            AP_AXIMM_52_WREADY,
    output  wire [1:0]                      AP_AXIMM_52_BRESP,
    output  wire                            AP_AXIMM_52_BVALID,
    input wire                            AP_AXIMM_52_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_52_ARADDR,
    input wire [7:0]                      AP_AXIMM_52_ARLEN,
    input wire [2:0]                      AP_AXIMM_52_ARSIZE,
    input wire [1:0]                      AP_AXIMM_52_ARBURST,
    input wire [1:0]                      AP_AXIMM_52_ARLOCK,
    input wire [3:0]                      AP_AXIMM_52_ARCACHE,
    input wire [2:0]                      AP_AXIMM_52_ARPROT,
    input wire [3:0]                      AP_AXIMM_52_ARREGION,
    input wire [3:0]                      AP_AXIMM_52_ARQOS,
    input wire                            AP_AXIMM_52_ARVALID,
    output  wire                            AP_AXIMM_52_ARREADY,
    output  wire [M_AXIMM_52_DATA_WIDTH-1:0]   AP_AXIMM_52_RDATA,
    output  wire [1:0]                      AP_AXIMM_52_RRESP,
    output  wire                            AP_AXIMM_52_RLAST,
    output  wire                            AP_AXIMM_52_RVALID,
    input  wire                            AP_AXIMM_52_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_52_AWADDR,
    output wire [7:0]                      M_AXIMM_52_AWLEN,
    output wire [2:0]                      M_AXIMM_52_AWSIZE,
    output wire [1:0]                      M_AXIMM_52_AWBURST,
    output wire [1:0]                      M_AXIMM_52_AWLOCK,
    output wire [3:0]                      M_AXIMM_52_AWCACHE,
    output wire [2:0]                      M_AXIMM_52_AWPROT,
    output wire [3:0]                      M_AXIMM_52_AWREGION,
    output wire [3:0]                      M_AXIMM_52_AWQOS,
    output wire                            M_AXIMM_52_AWVALID,
    input  wire                            M_AXIMM_52_AWREADY,
    output wire [M_AXIMM_52_DATA_WIDTH-1:0]   M_AXIMM_52_WDATA,
    output wire [M_AXIMM_52_DATA_WIDTH/8-1:0] M_AXIMM_52_WSTRB,
    output wire                            M_AXIMM_52_WLAST,
    output wire                            M_AXIMM_52_WVALID,
    input  wire                            M_AXIMM_52_WREADY,
    input  wire [1:0]                      M_AXIMM_52_BRESP,
    input  wire                            M_AXIMM_52_BVALID,
    output wire                            M_AXIMM_52_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_52_ARADDR,
    output wire [7:0]                      M_AXIMM_52_ARLEN,
    output wire [2:0]                      M_AXIMM_52_ARSIZE,
    output wire [1:0]                      M_AXIMM_52_ARBURST,
    output wire [1:0]                      M_AXIMM_52_ARLOCK,
    output wire [3:0]                      M_AXIMM_52_ARCACHE,
    output wire [2:0]                      M_AXIMM_52_ARPROT,
    output wire [3:0]                      M_AXIMM_52_ARREGION,
    output wire [3:0]                      M_AXIMM_52_ARQOS,
    output wire                            M_AXIMM_52_ARVALID,
    input  wire                            M_AXIMM_52_ARREADY,
    input  wire [M_AXIMM_52_DATA_WIDTH-1:0]   M_AXIMM_52_RDATA,
    input  wire [1:0]                      M_AXIMM_52_RRESP,
    input  wire                            M_AXIMM_52_RLAST,
    input  wire                            M_AXIMM_52_RVALID,
    output wire                            M_AXIMM_52_RREADY,
    //AXI-MM pass-through interface 53
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_53_AWADDR,
    input wire [7:0]                      AP_AXIMM_53_AWLEN,
    input wire [2:0]                      AP_AXIMM_53_AWSIZE,
    input wire [1:0]                      AP_AXIMM_53_AWBURST,
    input wire [1:0]                      AP_AXIMM_53_AWLOCK,
    input wire [3:0]                      AP_AXIMM_53_AWCACHE,
    input wire [2:0]                      AP_AXIMM_53_AWPROT,
    input wire [3:0]                      AP_AXIMM_53_AWREGION,
    input wire [3:0]                      AP_AXIMM_53_AWQOS,
    input wire                            AP_AXIMM_53_AWVALID,
    output  wire                            AP_AXIMM_53_AWREADY,
    input wire [M_AXIMM_53_DATA_WIDTH-1:0]   AP_AXIMM_53_WDATA,
    input wire [M_AXIMM_53_DATA_WIDTH/8-1:0] AP_AXIMM_53_WSTRB,
    input wire                            AP_AXIMM_53_WLAST,
    input wire                            AP_AXIMM_53_WVALID,
    output  wire                            AP_AXIMM_53_WREADY,
    output  wire [1:0]                      AP_AXIMM_53_BRESP,
    output  wire                            AP_AXIMM_53_BVALID,
    input wire                            AP_AXIMM_53_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_53_ARADDR,
    input wire [7:0]                      AP_AXIMM_53_ARLEN,
    input wire [2:0]                      AP_AXIMM_53_ARSIZE,
    input wire [1:0]                      AP_AXIMM_53_ARBURST,
    input wire [1:0]                      AP_AXIMM_53_ARLOCK,
    input wire [3:0]                      AP_AXIMM_53_ARCACHE,
    input wire [2:0]                      AP_AXIMM_53_ARPROT,
    input wire [3:0]                      AP_AXIMM_53_ARREGION,
    input wire [3:0]                      AP_AXIMM_53_ARQOS,
    input wire                            AP_AXIMM_53_ARVALID,
    output  wire                            AP_AXIMM_53_ARREADY,
    output  wire [M_AXIMM_53_DATA_WIDTH-1:0]   AP_AXIMM_53_RDATA,
    output  wire [1:0]                      AP_AXIMM_53_RRESP,
    output  wire                            AP_AXIMM_53_RLAST,
    output  wire                            AP_AXIMM_53_RVALID,
    input  wire                            AP_AXIMM_53_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_53_AWADDR,
    output wire [7:0]                      M_AXIMM_53_AWLEN,
    output wire [2:0]                      M_AXIMM_53_AWSIZE,
    output wire [1:0]                      M_AXIMM_53_AWBURST,
    output wire [1:0]                      M_AXIMM_53_AWLOCK,
    output wire [3:0]                      M_AXIMM_53_AWCACHE,
    output wire [2:0]                      M_AXIMM_53_AWPROT,
    output wire [3:0]                      M_AXIMM_53_AWREGION,
    output wire [3:0]                      M_AXIMM_53_AWQOS,
    output wire                            M_AXIMM_53_AWVALID,
    input  wire                            M_AXIMM_53_AWREADY,
    output wire [M_AXIMM_53_DATA_WIDTH-1:0]   M_AXIMM_53_WDATA,
    output wire [M_AXIMM_53_DATA_WIDTH/8-1:0] M_AXIMM_53_WSTRB,
    output wire                            M_AXIMM_53_WLAST,
    output wire                            M_AXIMM_53_WVALID,
    input  wire                            M_AXIMM_53_WREADY,
    input  wire [1:0]                      M_AXIMM_53_BRESP,
    input  wire                            M_AXIMM_53_BVALID,
    output wire                            M_AXIMM_53_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_53_ARADDR,
    output wire [7:0]                      M_AXIMM_53_ARLEN,
    output wire [2:0]                      M_AXIMM_53_ARSIZE,
    output wire [1:0]                      M_AXIMM_53_ARBURST,
    output wire [1:0]                      M_AXIMM_53_ARLOCK,
    output wire [3:0]                      M_AXIMM_53_ARCACHE,
    output wire [2:0]                      M_AXIMM_53_ARPROT,
    output wire [3:0]                      M_AXIMM_53_ARREGION,
    output wire [3:0]                      M_AXIMM_53_ARQOS,
    output wire                            M_AXIMM_53_ARVALID,
    input  wire                            M_AXIMM_53_ARREADY,
    input  wire [M_AXIMM_53_DATA_WIDTH-1:0]   M_AXIMM_53_RDATA,
    input  wire [1:0]                      M_AXIMM_53_RRESP,
    input  wire                            M_AXIMM_53_RLAST,
    input  wire                            M_AXIMM_53_RVALID,
    output wire                            M_AXIMM_53_RREADY,
    //AXI-MM pass-through interface 54
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_54_AWADDR,
    input wire [7:0]                      AP_AXIMM_54_AWLEN,
    input wire [2:0]                      AP_AXIMM_54_AWSIZE,
    input wire [1:0]                      AP_AXIMM_54_AWBURST,
    input wire [1:0]                      AP_AXIMM_54_AWLOCK,
    input wire [3:0]                      AP_AXIMM_54_AWCACHE,
    input wire [2:0]                      AP_AXIMM_54_AWPROT,
    input wire [3:0]                      AP_AXIMM_54_AWREGION,
    input wire [3:0]                      AP_AXIMM_54_AWQOS,
    input wire                            AP_AXIMM_54_AWVALID,
    output  wire                            AP_AXIMM_54_AWREADY,
    input wire [M_AXIMM_54_DATA_WIDTH-1:0]   AP_AXIMM_54_WDATA,
    input wire [M_AXIMM_54_DATA_WIDTH/8-1:0] AP_AXIMM_54_WSTRB,
    input wire                            AP_AXIMM_54_WLAST,
    input wire                            AP_AXIMM_54_WVALID,
    output  wire                            AP_AXIMM_54_WREADY,
    output  wire [1:0]                      AP_AXIMM_54_BRESP,
    output  wire                            AP_AXIMM_54_BVALID,
    input wire                            AP_AXIMM_54_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_54_ARADDR,
    input wire [7:0]                      AP_AXIMM_54_ARLEN,
    input wire [2:0]                      AP_AXIMM_54_ARSIZE,
    input wire [1:0]                      AP_AXIMM_54_ARBURST,
    input wire [1:0]                      AP_AXIMM_54_ARLOCK,
    input wire [3:0]                      AP_AXIMM_54_ARCACHE,
    input wire [2:0]                      AP_AXIMM_54_ARPROT,
    input wire [3:0]                      AP_AXIMM_54_ARREGION,
    input wire [3:0]                      AP_AXIMM_54_ARQOS,
    input wire                            AP_AXIMM_54_ARVALID,
    output  wire                            AP_AXIMM_54_ARREADY,
    output  wire [M_AXIMM_54_DATA_WIDTH-1:0]   AP_AXIMM_54_RDATA,
    output  wire [1:0]                      AP_AXIMM_54_RRESP,
    output  wire                            AP_AXIMM_54_RLAST,
    output  wire                            AP_AXIMM_54_RVALID,
    input  wire                            AP_AXIMM_54_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_54_AWADDR,
    output wire [7:0]                      M_AXIMM_54_AWLEN,
    output wire [2:0]                      M_AXIMM_54_AWSIZE,
    output wire [1:0]                      M_AXIMM_54_AWBURST,
    output wire [1:0]                      M_AXIMM_54_AWLOCK,
    output wire [3:0]                      M_AXIMM_54_AWCACHE,
    output wire [2:0]                      M_AXIMM_54_AWPROT,
    output wire [3:0]                      M_AXIMM_54_AWREGION,
    output wire [3:0]                      M_AXIMM_54_AWQOS,
    output wire                            M_AXIMM_54_AWVALID,
    input  wire                            M_AXIMM_54_AWREADY,
    output wire [M_AXIMM_54_DATA_WIDTH-1:0]   M_AXIMM_54_WDATA,
    output wire [M_AXIMM_54_DATA_WIDTH/8-1:0] M_AXIMM_54_WSTRB,
    output wire                            M_AXIMM_54_WLAST,
    output wire                            M_AXIMM_54_WVALID,
    input  wire                            M_AXIMM_54_WREADY,
    input  wire [1:0]                      M_AXIMM_54_BRESP,
    input  wire                            M_AXIMM_54_BVALID,
    output wire                            M_AXIMM_54_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_54_ARADDR,
    output wire [7:0]                      M_AXIMM_54_ARLEN,
    output wire [2:0]                      M_AXIMM_54_ARSIZE,
    output wire [1:0]                      M_AXIMM_54_ARBURST,
    output wire [1:0]                      M_AXIMM_54_ARLOCK,
    output wire [3:0]                      M_AXIMM_54_ARCACHE,
    output wire [2:0]                      M_AXIMM_54_ARPROT,
    output wire [3:0]                      M_AXIMM_54_ARREGION,
    output wire [3:0]                      M_AXIMM_54_ARQOS,
    output wire                            M_AXIMM_54_ARVALID,
    input  wire                            M_AXIMM_54_ARREADY,
    input  wire [M_AXIMM_54_DATA_WIDTH-1:0]   M_AXIMM_54_RDATA,
    input  wire [1:0]                      M_AXIMM_54_RRESP,
    input  wire                            M_AXIMM_54_RLAST,
    input  wire                            M_AXIMM_54_RVALID,
    output wire                            M_AXIMM_54_RREADY,
    //AXI-MM pass-through interface 55
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_55_AWADDR,
    input wire [7:0]                      AP_AXIMM_55_AWLEN,
    input wire [2:0]                      AP_AXIMM_55_AWSIZE,
    input wire [1:0]                      AP_AXIMM_55_AWBURST,
    input wire [1:0]                      AP_AXIMM_55_AWLOCK,
    input wire [3:0]                      AP_AXIMM_55_AWCACHE,
    input wire [2:0]                      AP_AXIMM_55_AWPROT,
    input wire [3:0]                      AP_AXIMM_55_AWREGION,
    input wire [3:0]                      AP_AXIMM_55_AWQOS,
    input wire                            AP_AXIMM_55_AWVALID,
    output  wire                            AP_AXIMM_55_AWREADY,
    input wire [M_AXIMM_55_DATA_WIDTH-1:0]   AP_AXIMM_55_WDATA,
    input wire [M_AXIMM_55_DATA_WIDTH/8-1:0] AP_AXIMM_55_WSTRB,
    input wire                            AP_AXIMM_55_WLAST,
    input wire                            AP_AXIMM_55_WVALID,
    output  wire                            AP_AXIMM_55_WREADY,
    output  wire [1:0]                      AP_AXIMM_55_BRESP,
    output  wire                            AP_AXIMM_55_BVALID,
    input wire                            AP_AXIMM_55_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_55_ARADDR,
    input wire [7:0]                      AP_AXIMM_55_ARLEN,
    input wire [2:0]                      AP_AXIMM_55_ARSIZE,
    input wire [1:0]                      AP_AXIMM_55_ARBURST,
    input wire [1:0]                      AP_AXIMM_55_ARLOCK,
    input wire [3:0]                      AP_AXIMM_55_ARCACHE,
    input wire [2:0]                      AP_AXIMM_55_ARPROT,
    input wire [3:0]                      AP_AXIMM_55_ARREGION,
    input wire [3:0]                      AP_AXIMM_55_ARQOS,
    input wire                            AP_AXIMM_55_ARVALID,
    output  wire                            AP_AXIMM_55_ARREADY,
    output  wire [M_AXIMM_55_DATA_WIDTH-1:0]   AP_AXIMM_55_RDATA,
    output  wire [1:0]                      AP_AXIMM_55_RRESP,
    output  wire                            AP_AXIMM_55_RLAST,
    output  wire                            AP_AXIMM_55_RVALID,
    input  wire                            AP_AXIMM_55_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_55_AWADDR,
    output wire [7:0]                      M_AXIMM_55_AWLEN,
    output wire [2:0]                      M_AXIMM_55_AWSIZE,
    output wire [1:0]                      M_AXIMM_55_AWBURST,
    output wire [1:0]                      M_AXIMM_55_AWLOCK,
    output wire [3:0]                      M_AXIMM_55_AWCACHE,
    output wire [2:0]                      M_AXIMM_55_AWPROT,
    output wire [3:0]                      M_AXIMM_55_AWREGION,
    output wire [3:0]                      M_AXIMM_55_AWQOS,
    output wire                            M_AXIMM_55_AWVALID,
    input  wire                            M_AXIMM_55_AWREADY,
    output wire [M_AXIMM_55_DATA_WIDTH-1:0]   M_AXIMM_55_WDATA,
    output wire [M_AXIMM_55_DATA_WIDTH/8-1:0] M_AXIMM_55_WSTRB,
    output wire                            M_AXIMM_55_WLAST,
    output wire                            M_AXIMM_55_WVALID,
    input  wire                            M_AXIMM_55_WREADY,
    input  wire [1:0]                      M_AXIMM_55_BRESP,
    input  wire                            M_AXIMM_55_BVALID,
    output wire                            M_AXIMM_55_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_55_ARADDR,
    output wire [7:0]                      M_AXIMM_55_ARLEN,
    output wire [2:0]                      M_AXIMM_55_ARSIZE,
    output wire [1:0]                      M_AXIMM_55_ARBURST,
    output wire [1:0]                      M_AXIMM_55_ARLOCK,
    output wire [3:0]                      M_AXIMM_55_ARCACHE,
    output wire [2:0]                      M_AXIMM_55_ARPROT,
    output wire [3:0]                      M_AXIMM_55_ARREGION,
    output wire [3:0]                      M_AXIMM_55_ARQOS,
    output wire                            M_AXIMM_55_ARVALID,
    input  wire                            M_AXIMM_55_ARREADY,
    input  wire [M_AXIMM_55_DATA_WIDTH-1:0]   M_AXIMM_55_RDATA,
    input  wire [1:0]                      M_AXIMM_55_RRESP,
    input  wire                            M_AXIMM_55_RLAST,
    input  wire                            M_AXIMM_55_RVALID,
    output wire                            M_AXIMM_55_RREADY,
    //AXI-MM pass-through interface 56
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_56_AWADDR,
    input wire [7:0]                      AP_AXIMM_56_AWLEN,
    input wire [2:0]                      AP_AXIMM_56_AWSIZE,
    input wire [1:0]                      AP_AXIMM_56_AWBURST,
    input wire [1:0]                      AP_AXIMM_56_AWLOCK,
    input wire [3:0]                      AP_AXIMM_56_AWCACHE,
    input wire [2:0]                      AP_AXIMM_56_AWPROT,
    input wire [3:0]                      AP_AXIMM_56_AWREGION,
    input wire [3:0]                      AP_AXIMM_56_AWQOS,
    input wire                            AP_AXIMM_56_AWVALID,
    output  wire                            AP_AXIMM_56_AWREADY,
    input wire [M_AXIMM_56_DATA_WIDTH-1:0]   AP_AXIMM_56_WDATA,
    input wire [M_AXIMM_56_DATA_WIDTH/8-1:0] AP_AXIMM_56_WSTRB,
    input wire                            AP_AXIMM_56_WLAST,
    input wire                            AP_AXIMM_56_WVALID,
    output  wire                            AP_AXIMM_56_WREADY,
    output  wire [1:0]                      AP_AXIMM_56_BRESP,
    output  wire                            AP_AXIMM_56_BVALID,
    input wire                            AP_AXIMM_56_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_56_ARADDR,
    input wire [7:0]                      AP_AXIMM_56_ARLEN,
    input wire [2:0]                      AP_AXIMM_56_ARSIZE,
    input wire [1:0]                      AP_AXIMM_56_ARBURST,
    input wire [1:0]                      AP_AXIMM_56_ARLOCK,
    input wire [3:0]                      AP_AXIMM_56_ARCACHE,
    input wire [2:0]                      AP_AXIMM_56_ARPROT,
    input wire [3:0]                      AP_AXIMM_56_ARREGION,
    input wire [3:0]                      AP_AXIMM_56_ARQOS,
    input wire                            AP_AXIMM_56_ARVALID,
    output  wire                            AP_AXIMM_56_ARREADY,
    output  wire [M_AXIMM_56_DATA_WIDTH-1:0]   AP_AXIMM_56_RDATA,
    output  wire [1:0]                      AP_AXIMM_56_RRESP,
    output  wire                            AP_AXIMM_56_RLAST,
    output  wire                            AP_AXIMM_56_RVALID,
    input  wire                            AP_AXIMM_56_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_56_AWADDR,
    output wire [7:0]                      M_AXIMM_56_AWLEN,
    output wire [2:0]                      M_AXIMM_56_AWSIZE,
    output wire [1:0]                      M_AXIMM_56_AWBURST,
    output wire [1:0]                      M_AXIMM_56_AWLOCK,
    output wire [3:0]                      M_AXIMM_56_AWCACHE,
    output wire [2:0]                      M_AXIMM_56_AWPROT,
    output wire [3:0]                      M_AXIMM_56_AWREGION,
    output wire [3:0]                      M_AXIMM_56_AWQOS,
    output wire                            M_AXIMM_56_AWVALID,
    input  wire                            M_AXIMM_56_AWREADY,
    output wire [M_AXIMM_56_DATA_WIDTH-1:0]   M_AXIMM_56_WDATA,
    output wire [M_AXIMM_56_DATA_WIDTH/8-1:0] M_AXIMM_56_WSTRB,
    output wire                            M_AXIMM_56_WLAST,
    output wire                            M_AXIMM_56_WVALID,
    input  wire                            M_AXIMM_56_WREADY,
    input  wire [1:0]                      M_AXIMM_56_BRESP,
    input  wire                            M_AXIMM_56_BVALID,
    output wire                            M_AXIMM_56_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_56_ARADDR,
    output wire [7:0]                      M_AXIMM_56_ARLEN,
    output wire [2:0]                      M_AXIMM_56_ARSIZE,
    output wire [1:0]                      M_AXIMM_56_ARBURST,
    output wire [1:0]                      M_AXIMM_56_ARLOCK,
    output wire [3:0]                      M_AXIMM_56_ARCACHE,
    output wire [2:0]                      M_AXIMM_56_ARPROT,
    output wire [3:0]                      M_AXIMM_56_ARREGION,
    output wire [3:0]                      M_AXIMM_56_ARQOS,
    output wire                            M_AXIMM_56_ARVALID,
    input  wire                            M_AXIMM_56_ARREADY,
    input  wire [M_AXIMM_56_DATA_WIDTH-1:0]   M_AXIMM_56_RDATA,
    input  wire [1:0]                      M_AXIMM_56_RRESP,
    input  wire                            M_AXIMM_56_RLAST,
    input  wire                            M_AXIMM_56_RVALID,
    output wire                            M_AXIMM_56_RREADY,
    //AXI-MM pass-through interface 57
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_57_AWADDR,
    input wire [7:0]                      AP_AXIMM_57_AWLEN,
    input wire [2:0]                      AP_AXIMM_57_AWSIZE,
    input wire [1:0]                      AP_AXIMM_57_AWBURST,
    input wire [1:0]                      AP_AXIMM_57_AWLOCK,
    input wire [3:0]                      AP_AXIMM_57_AWCACHE,
    input wire [2:0]                      AP_AXIMM_57_AWPROT,
    input wire [3:0]                      AP_AXIMM_57_AWREGION,
    input wire [3:0]                      AP_AXIMM_57_AWQOS,
    input wire                            AP_AXIMM_57_AWVALID,
    output  wire                            AP_AXIMM_57_AWREADY,
    input wire [M_AXIMM_57_DATA_WIDTH-1:0]   AP_AXIMM_57_WDATA,
    input wire [M_AXIMM_57_DATA_WIDTH/8-1:0] AP_AXIMM_57_WSTRB,
    input wire                            AP_AXIMM_57_WLAST,
    input wire                            AP_AXIMM_57_WVALID,
    output  wire                            AP_AXIMM_57_WREADY,
    output  wire [1:0]                      AP_AXIMM_57_BRESP,
    output  wire                            AP_AXIMM_57_BVALID,
    input wire                            AP_AXIMM_57_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_57_ARADDR,
    input wire [7:0]                      AP_AXIMM_57_ARLEN,
    input wire [2:0]                      AP_AXIMM_57_ARSIZE,
    input wire [1:0]                      AP_AXIMM_57_ARBURST,
    input wire [1:0]                      AP_AXIMM_57_ARLOCK,
    input wire [3:0]                      AP_AXIMM_57_ARCACHE,
    input wire [2:0]                      AP_AXIMM_57_ARPROT,
    input wire [3:0]                      AP_AXIMM_57_ARREGION,
    input wire [3:0]                      AP_AXIMM_57_ARQOS,
    input wire                            AP_AXIMM_57_ARVALID,
    output  wire                            AP_AXIMM_57_ARREADY,
    output  wire [M_AXIMM_57_DATA_WIDTH-1:0]   AP_AXIMM_57_RDATA,
    output  wire [1:0]                      AP_AXIMM_57_RRESP,
    output  wire                            AP_AXIMM_57_RLAST,
    output  wire                            AP_AXIMM_57_RVALID,
    input  wire                            AP_AXIMM_57_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_57_AWADDR,
    output wire [7:0]                      M_AXIMM_57_AWLEN,
    output wire [2:0]                      M_AXIMM_57_AWSIZE,
    output wire [1:0]                      M_AXIMM_57_AWBURST,
    output wire [1:0]                      M_AXIMM_57_AWLOCK,
    output wire [3:0]                      M_AXIMM_57_AWCACHE,
    output wire [2:0]                      M_AXIMM_57_AWPROT,
    output wire [3:0]                      M_AXIMM_57_AWREGION,
    output wire [3:0]                      M_AXIMM_57_AWQOS,
    output wire                            M_AXIMM_57_AWVALID,
    input  wire                            M_AXIMM_57_AWREADY,
    output wire [M_AXIMM_57_DATA_WIDTH-1:0]   M_AXIMM_57_WDATA,
    output wire [M_AXIMM_57_DATA_WIDTH/8-1:0] M_AXIMM_57_WSTRB,
    output wire                            M_AXIMM_57_WLAST,
    output wire                            M_AXIMM_57_WVALID,
    input  wire                            M_AXIMM_57_WREADY,
    input  wire [1:0]                      M_AXIMM_57_BRESP,
    input  wire                            M_AXIMM_57_BVALID,
    output wire                            M_AXIMM_57_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_57_ARADDR,
    output wire [7:0]                      M_AXIMM_57_ARLEN,
    output wire [2:0]                      M_AXIMM_57_ARSIZE,
    output wire [1:0]                      M_AXIMM_57_ARBURST,
    output wire [1:0]                      M_AXIMM_57_ARLOCK,
    output wire [3:0]                      M_AXIMM_57_ARCACHE,
    output wire [2:0]                      M_AXIMM_57_ARPROT,
    output wire [3:0]                      M_AXIMM_57_ARREGION,
    output wire [3:0]                      M_AXIMM_57_ARQOS,
    output wire                            M_AXIMM_57_ARVALID,
    input  wire                            M_AXIMM_57_ARREADY,
    input  wire [M_AXIMM_57_DATA_WIDTH-1:0]   M_AXIMM_57_RDATA,
    input  wire [1:0]                      M_AXIMM_57_RRESP,
    input  wire                            M_AXIMM_57_RLAST,
    input  wire                            M_AXIMM_57_RVALID,
    output wire                            M_AXIMM_57_RREADY,
    //AXI-MM pass-through interface 58
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_58_AWADDR,
    input wire [7:0]                      AP_AXIMM_58_AWLEN,
    input wire [2:0]                      AP_AXIMM_58_AWSIZE,
    input wire [1:0]                      AP_AXIMM_58_AWBURST,
    input wire [1:0]                      AP_AXIMM_58_AWLOCK,
    input wire [3:0]                      AP_AXIMM_58_AWCACHE,
    input wire [2:0]                      AP_AXIMM_58_AWPROT,
    input wire [3:0]                      AP_AXIMM_58_AWREGION,
    input wire [3:0]                      AP_AXIMM_58_AWQOS,
    input wire                            AP_AXIMM_58_AWVALID,
    output  wire                            AP_AXIMM_58_AWREADY,
    input wire [M_AXIMM_58_DATA_WIDTH-1:0]   AP_AXIMM_58_WDATA,
    input wire [M_AXIMM_58_DATA_WIDTH/8-1:0] AP_AXIMM_58_WSTRB,
    input wire                            AP_AXIMM_58_WLAST,
    input wire                            AP_AXIMM_58_WVALID,
    output  wire                            AP_AXIMM_58_WREADY,
    output  wire [1:0]                      AP_AXIMM_58_BRESP,
    output  wire                            AP_AXIMM_58_BVALID,
    input wire                            AP_AXIMM_58_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_58_ARADDR,
    input wire [7:0]                      AP_AXIMM_58_ARLEN,
    input wire [2:0]                      AP_AXIMM_58_ARSIZE,
    input wire [1:0]                      AP_AXIMM_58_ARBURST,
    input wire [1:0]                      AP_AXIMM_58_ARLOCK,
    input wire [3:0]                      AP_AXIMM_58_ARCACHE,
    input wire [2:0]                      AP_AXIMM_58_ARPROT,
    input wire [3:0]                      AP_AXIMM_58_ARREGION,
    input wire [3:0]                      AP_AXIMM_58_ARQOS,
    input wire                            AP_AXIMM_58_ARVALID,
    output  wire                            AP_AXIMM_58_ARREADY,
    output  wire [M_AXIMM_58_DATA_WIDTH-1:0]   AP_AXIMM_58_RDATA,
    output  wire [1:0]                      AP_AXIMM_58_RRESP,
    output  wire                            AP_AXIMM_58_RLAST,
    output  wire                            AP_AXIMM_58_RVALID,
    input  wire                            AP_AXIMM_58_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_58_AWADDR,
    output wire [7:0]                      M_AXIMM_58_AWLEN,
    output wire [2:0]                      M_AXIMM_58_AWSIZE,
    output wire [1:0]                      M_AXIMM_58_AWBURST,
    output wire [1:0]                      M_AXIMM_58_AWLOCK,
    output wire [3:0]                      M_AXIMM_58_AWCACHE,
    output wire [2:0]                      M_AXIMM_58_AWPROT,
    output wire [3:0]                      M_AXIMM_58_AWREGION,
    output wire [3:0]                      M_AXIMM_58_AWQOS,
    output wire                            M_AXIMM_58_AWVALID,
    input  wire                            M_AXIMM_58_AWREADY,
    output wire [M_AXIMM_58_DATA_WIDTH-1:0]   M_AXIMM_58_WDATA,
    output wire [M_AXIMM_58_DATA_WIDTH/8-1:0] M_AXIMM_58_WSTRB,
    output wire                            M_AXIMM_58_WLAST,
    output wire                            M_AXIMM_58_WVALID,
    input  wire                            M_AXIMM_58_WREADY,
    input  wire [1:0]                      M_AXIMM_58_BRESP,
    input  wire                            M_AXIMM_58_BVALID,
    output wire                            M_AXIMM_58_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_58_ARADDR,
    output wire [7:0]                      M_AXIMM_58_ARLEN,
    output wire [2:0]                      M_AXIMM_58_ARSIZE,
    output wire [1:0]                      M_AXIMM_58_ARBURST,
    output wire [1:0]                      M_AXIMM_58_ARLOCK,
    output wire [3:0]                      M_AXIMM_58_ARCACHE,
    output wire [2:0]                      M_AXIMM_58_ARPROT,
    output wire [3:0]                      M_AXIMM_58_ARREGION,
    output wire [3:0]                      M_AXIMM_58_ARQOS,
    output wire                            M_AXIMM_58_ARVALID,
    input  wire                            M_AXIMM_58_ARREADY,
    input  wire [M_AXIMM_58_DATA_WIDTH-1:0]   M_AXIMM_58_RDATA,
    input  wire [1:0]                      M_AXIMM_58_RRESP,
    input  wire                            M_AXIMM_58_RLAST,
    input  wire                            M_AXIMM_58_RVALID,
    output wire                            M_AXIMM_58_RREADY,
    //AXI-MM pass-through interface 59
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_59_AWADDR,
    input wire [7:0]                      AP_AXIMM_59_AWLEN,
    input wire [2:0]                      AP_AXIMM_59_AWSIZE,
    input wire [1:0]                      AP_AXIMM_59_AWBURST,
    input wire [1:0]                      AP_AXIMM_59_AWLOCK,
    input wire [3:0]                      AP_AXIMM_59_AWCACHE,
    input wire [2:0]                      AP_AXIMM_59_AWPROT,
    input wire [3:0]                      AP_AXIMM_59_AWREGION,
    input wire [3:0]                      AP_AXIMM_59_AWQOS,
    input wire                            AP_AXIMM_59_AWVALID,
    output  wire                            AP_AXIMM_59_AWREADY,
    input wire [M_AXIMM_59_DATA_WIDTH-1:0]   AP_AXIMM_59_WDATA,
    input wire [M_AXIMM_59_DATA_WIDTH/8-1:0] AP_AXIMM_59_WSTRB,
    input wire                            AP_AXIMM_59_WLAST,
    input wire                            AP_AXIMM_59_WVALID,
    output  wire                            AP_AXIMM_59_WREADY,
    output  wire [1:0]                      AP_AXIMM_59_BRESP,
    output  wire                            AP_AXIMM_59_BVALID,
    input wire                            AP_AXIMM_59_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_59_ARADDR,
    input wire [7:0]                      AP_AXIMM_59_ARLEN,
    input wire [2:0]                      AP_AXIMM_59_ARSIZE,
    input wire [1:0]                      AP_AXIMM_59_ARBURST,
    input wire [1:0]                      AP_AXIMM_59_ARLOCK,
    input wire [3:0]                      AP_AXIMM_59_ARCACHE,
    input wire [2:0]                      AP_AXIMM_59_ARPROT,
    input wire [3:0]                      AP_AXIMM_59_ARREGION,
    input wire [3:0]                      AP_AXIMM_59_ARQOS,
    input wire                            AP_AXIMM_59_ARVALID,
    output  wire                            AP_AXIMM_59_ARREADY,
    output  wire [M_AXIMM_59_DATA_WIDTH-1:0]   AP_AXIMM_59_RDATA,
    output  wire [1:0]                      AP_AXIMM_59_RRESP,
    output  wire                            AP_AXIMM_59_RLAST,
    output  wire                            AP_AXIMM_59_RVALID,
    input  wire                            AP_AXIMM_59_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_59_AWADDR,
    output wire [7:0]                      M_AXIMM_59_AWLEN,
    output wire [2:0]                      M_AXIMM_59_AWSIZE,
    output wire [1:0]                      M_AXIMM_59_AWBURST,
    output wire [1:0]                      M_AXIMM_59_AWLOCK,
    output wire [3:0]                      M_AXIMM_59_AWCACHE,
    output wire [2:0]                      M_AXIMM_59_AWPROT,
    output wire [3:0]                      M_AXIMM_59_AWREGION,
    output wire [3:0]                      M_AXIMM_59_AWQOS,
    output wire                            M_AXIMM_59_AWVALID,
    input  wire                            M_AXIMM_59_AWREADY,
    output wire [M_AXIMM_59_DATA_WIDTH-1:0]   M_AXIMM_59_WDATA,
    output wire [M_AXIMM_59_DATA_WIDTH/8-1:0] M_AXIMM_59_WSTRB,
    output wire                            M_AXIMM_59_WLAST,
    output wire                            M_AXIMM_59_WVALID,
    input  wire                            M_AXIMM_59_WREADY,
    input  wire [1:0]                      M_AXIMM_59_BRESP,
    input  wire                            M_AXIMM_59_BVALID,
    output wire                            M_AXIMM_59_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_59_ARADDR,
    output wire [7:0]                      M_AXIMM_59_ARLEN,
    output wire [2:0]                      M_AXIMM_59_ARSIZE,
    output wire [1:0]                      M_AXIMM_59_ARBURST,
    output wire [1:0]                      M_AXIMM_59_ARLOCK,
    output wire [3:0]                      M_AXIMM_59_ARCACHE,
    output wire [2:0]                      M_AXIMM_59_ARPROT,
    output wire [3:0]                      M_AXIMM_59_ARREGION,
    output wire [3:0]                      M_AXIMM_59_ARQOS,
    output wire                            M_AXIMM_59_ARVALID,
    input  wire                            M_AXIMM_59_ARREADY,
    input  wire [M_AXIMM_59_DATA_WIDTH-1:0]   M_AXIMM_59_RDATA,
    input  wire [1:0]                      M_AXIMM_59_RRESP,
    input  wire                            M_AXIMM_59_RLAST,
    input  wire                            M_AXIMM_59_RVALID,
    output wire                            M_AXIMM_59_RREADY,
    //AXI-MM pass-through interface 60
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_60_AWADDR,
    input wire [7:0]                      AP_AXIMM_60_AWLEN,
    input wire [2:0]                      AP_AXIMM_60_AWSIZE,
    input wire [1:0]                      AP_AXIMM_60_AWBURST,
    input wire [1:0]                      AP_AXIMM_60_AWLOCK,
    input wire [3:0]                      AP_AXIMM_60_AWCACHE,
    input wire [2:0]                      AP_AXIMM_60_AWPROT,
    input wire [3:0]                      AP_AXIMM_60_AWREGION,
    input wire [3:0]                      AP_AXIMM_60_AWQOS,
    input wire                            AP_AXIMM_60_AWVALID,
    output  wire                            AP_AXIMM_60_AWREADY,
    input wire [M_AXIMM_60_DATA_WIDTH-1:0]   AP_AXIMM_60_WDATA,
    input wire [M_AXIMM_60_DATA_WIDTH/8-1:0] AP_AXIMM_60_WSTRB,
    input wire                            AP_AXIMM_60_WLAST,
    input wire                            AP_AXIMM_60_WVALID,
    output  wire                            AP_AXIMM_60_WREADY,
    output  wire [1:0]                      AP_AXIMM_60_BRESP,
    output  wire                            AP_AXIMM_60_BVALID,
    input wire                            AP_AXIMM_60_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_60_ARADDR,
    input wire [7:0]                      AP_AXIMM_60_ARLEN,
    input wire [2:0]                      AP_AXIMM_60_ARSIZE,
    input wire [1:0]                      AP_AXIMM_60_ARBURST,
    input wire [1:0]                      AP_AXIMM_60_ARLOCK,
    input wire [3:0]                      AP_AXIMM_60_ARCACHE,
    input wire [2:0]                      AP_AXIMM_60_ARPROT,
    input wire [3:0]                      AP_AXIMM_60_ARREGION,
    input wire [3:0]                      AP_AXIMM_60_ARQOS,
    input wire                            AP_AXIMM_60_ARVALID,
    output  wire                            AP_AXIMM_60_ARREADY,
    output  wire [M_AXIMM_60_DATA_WIDTH-1:0]   AP_AXIMM_60_RDATA,
    output  wire [1:0]                      AP_AXIMM_60_RRESP,
    output  wire                            AP_AXIMM_60_RLAST,
    output  wire                            AP_AXIMM_60_RVALID,
    input  wire                            AP_AXIMM_60_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_60_AWADDR,
    output wire [7:0]                      M_AXIMM_60_AWLEN,
    output wire [2:0]                      M_AXIMM_60_AWSIZE,
    output wire [1:0]                      M_AXIMM_60_AWBURST,
    output wire [1:0]                      M_AXIMM_60_AWLOCK,
    output wire [3:0]                      M_AXIMM_60_AWCACHE,
    output wire [2:0]                      M_AXIMM_60_AWPROT,
    output wire [3:0]                      M_AXIMM_60_AWREGION,
    output wire [3:0]                      M_AXIMM_60_AWQOS,
    output wire                            M_AXIMM_60_AWVALID,
    input  wire                            M_AXIMM_60_AWREADY,
    output wire [M_AXIMM_60_DATA_WIDTH-1:0]   M_AXIMM_60_WDATA,
    output wire [M_AXIMM_60_DATA_WIDTH/8-1:0] M_AXIMM_60_WSTRB,
    output wire                            M_AXIMM_60_WLAST,
    output wire                            M_AXIMM_60_WVALID,
    input  wire                            M_AXIMM_60_WREADY,
    input  wire [1:0]                      M_AXIMM_60_BRESP,
    input  wire                            M_AXIMM_60_BVALID,
    output wire                            M_AXIMM_60_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_60_ARADDR,
    output wire [7:0]                      M_AXIMM_60_ARLEN,
    output wire [2:0]                      M_AXIMM_60_ARSIZE,
    output wire [1:0]                      M_AXIMM_60_ARBURST,
    output wire [1:0]                      M_AXIMM_60_ARLOCK,
    output wire [3:0]                      M_AXIMM_60_ARCACHE,
    output wire [2:0]                      M_AXIMM_60_ARPROT,
    output wire [3:0]                      M_AXIMM_60_ARREGION,
    output wire [3:0]                      M_AXIMM_60_ARQOS,
    output wire                            M_AXIMM_60_ARVALID,
    input  wire                            M_AXIMM_60_ARREADY,
    input  wire [M_AXIMM_60_DATA_WIDTH-1:0]   M_AXIMM_60_RDATA,
    input  wire [1:0]                      M_AXIMM_60_RRESP,
    input  wire                            M_AXIMM_60_RLAST,
    input  wire                            M_AXIMM_60_RVALID,
    output wire                            M_AXIMM_60_RREADY,
    //AXI-MM pass-through interface 61
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_61_AWADDR,
    input wire [7:0]                      AP_AXIMM_61_AWLEN,
    input wire [2:0]                      AP_AXIMM_61_AWSIZE,
    input wire [1:0]                      AP_AXIMM_61_AWBURST,
    input wire [1:0]                      AP_AXIMM_61_AWLOCK,
    input wire [3:0]                      AP_AXIMM_61_AWCACHE,
    input wire [2:0]                      AP_AXIMM_61_AWPROT,
    input wire [3:0]                      AP_AXIMM_61_AWREGION,
    input wire [3:0]                      AP_AXIMM_61_AWQOS,
    input wire                            AP_AXIMM_61_AWVALID,
    output  wire                            AP_AXIMM_61_AWREADY,
    input wire [M_AXIMM_61_DATA_WIDTH-1:0]   AP_AXIMM_61_WDATA,
    input wire [M_AXIMM_61_DATA_WIDTH/8-1:0] AP_AXIMM_61_WSTRB,
    input wire                            AP_AXIMM_61_WLAST,
    input wire                            AP_AXIMM_61_WVALID,
    output  wire                            AP_AXIMM_61_WREADY,
    output  wire [1:0]                      AP_AXIMM_61_BRESP,
    output  wire                            AP_AXIMM_61_BVALID,
    input wire                            AP_AXIMM_61_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_61_ARADDR,
    input wire [7:0]                      AP_AXIMM_61_ARLEN,
    input wire [2:0]                      AP_AXIMM_61_ARSIZE,
    input wire [1:0]                      AP_AXIMM_61_ARBURST,
    input wire [1:0]                      AP_AXIMM_61_ARLOCK,
    input wire [3:0]                      AP_AXIMM_61_ARCACHE,
    input wire [2:0]                      AP_AXIMM_61_ARPROT,
    input wire [3:0]                      AP_AXIMM_61_ARREGION,
    input wire [3:0]                      AP_AXIMM_61_ARQOS,
    input wire                            AP_AXIMM_61_ARVALID,
    output  wire                            AP_AXIMM_61_ARREADY,
    output  wire [M_AXIMM_61_DATA_WIDTH-1:0]   AP_AXIMM_61_RDATA,
    output  wire [1:0]                      AP_AXIMM_61_RRESP,
    output  wire                            AP_AXIMM_61_RLAST,
    output  wire                            AP_AXIMM_61_RVALID,
    input  wire                            AP_AXIMM_61_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_61_AWADDR,
    output wire [7:0]                      M_AXIMM_61_AWLEN,
    output wire [2:0]                      M_AXIMM_61_AWSIZE,
    output wire [1:0]                      M_AXIMM_61_AWBURST,
    output wire [1:0]                      M_AXIMM_61_AWLOCK,
    output wire [3:0]                      M_AXIMM_61_AWCACHE,
    output wire [2:0]                      M_AXIMM_61_AWPROT,
    output wire [3:0]                      M_AXIMM_61_AWREGION,
    output wire [3:0]                      M_AXIMM_61_AWQOS,
    output wire                            M_AXIMM_61_AWVALID,
    input  wire                            M_AXIMM_61_AWREADY,
    output wire [M_AXIMM_61_DATA_WIDTH-1:0]   M_AXIMM_61_WDATA,
    output wire [M_AXIMM_61_DATA_WIDTH/8-1:0] M_AXIMM_61_WSTRB,
    output wire                            M_AXIMM_61_WLAST,
    output wire                            M_AXIMM_61_WVALID,
    input  wire                            M_AXIMM_61_WREADY,
    input  wire [1:0]                      M_AXIMM_61_BRESP,
    input  wire                            M_AXIMM_61_BVALID,
    output wire                            M_AXIMM_61_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_61_ARADDR,
    output wire [7:0]                      M_AXIMM_61_ARLEN,
    output wire [2:0]                      M_AXIMM_61_ARSIZE,
    output wire [1:0]                      M_AXIMM_61_ARBURST,
    output wire [1:0]                      M_AXIMM_61_ARLOCK,
    output wire [3:0]                      M_AXIMM_61_ARCACHE,
    output wire [2:0]                      M_AXIMM_61_ARPROT,
    output wire [3:0]                      M_AXIMM_61_ARREGION,
    output wire [3:0]                      M_AXIMM_61_ARQOS,
    output wire                            M_AXIMM_61_ARVALID,
    input  wire                            M_AXIMM_61_ARREADY,
    input  wire [M_AXIMM_61_DATA_WIDTH-1:0]   M_AXIMM_61_RDATA,
    input  wire [1:0]                      M_AXIMM_61_RRESP,
    input  wire                            M_AXIMM_61_RLAST,
    input  wire                            M_AXIMM_61_RVALID,
    output wire                            M_AXIMM_61_RREADY,
    //AXI-MM pass-through interface 62
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_62_AWADDR,
    input wire [7:0]                      AP_AXIMM_62_AWLEN,
    input wire [2:0]                      AP_AXIMM_62_AWSIZE,
    input wire [1:0]                      AP_AXIMM_62_AWBURST,
    input wire [1:0]                      AP_AXIMM_62_AWLOCK,
    input wire [3:0]                      AP_AXIMM_62_AWCACHE,
    input wire [2:0]                      AP_AXIMM_62_AWPROT,
    input wire [3:0]                      AP_AXIMM_62_AWREGION,
    input wire [3:0]                      AP_AXIMM_62_AWQOS,
    input wire                            AP_AXIMM_62_AWVALID,
    output  wire                            AP_AXIMM_62_AWREADY,
    input wire [M_AXIMM_62_DATA_WIDTH-1:0]   AP_AXIMM_62_WDATA,
    input wire [M_AXIMM_62_DATA_WIDTH/8-1:0] AP_AXIMM_62_WSTRB,
    input wire                            AP_AXIMM_62_WLAST,
    input wire                            AP_AXIMM_62_WVALID,
    output  wire                            AP_AXIMM_62_WREADY,
    output  wire [1:0]                      AP_AXIMM_62_BRESP,
    output  wire                            AP_AXIMM_62_BVALID,
    input wire                            AP_AXIMM_62_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_62_ARADDR,
    input wire [7:0]                      AP_AXIMM_62_ARLEN,
    input wire [2:0]                      AP_AXIMM_62_ARSIZE,
    input wire [1:0]                      AP_AXIMM_62_ARBURST,
    input wire [1:0]                      AP_AXIMM_62_ARLOCK,
    input wire [3:0]                      AP_AXIMM_62_ARCACHE,
    input wire [2:0]                      AP_AXIMM_62_ARPROT,
    input wire [3:0]                      AP_AXIMM_62_ARREGION,
    input wire [3:0]                      AP_AXIMM_62_ARQOS,
    input wire                            AP_AXIMM_62_ARVALID,
    output  wire                            AP_AXIMM_62_ARREADY,
    output  wire [M_AXIMM_62_DATA_WIDTH-1:0]   AP_AXIMM_62_RDATA,
    output  wire [1:0]                      AP_AXIMM_62_RRESP,
    output  wire                            AP_AXIMM_62_RLAST,
    output  wire                            AP_AXIMM_62_RVALID,
    input  wire                            AP_AXIMM_62_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_62_AWADDR,
    output wire [7:0]                      M_AXIMM_62_AWLEN,
    output wire [2:0]                      M_AXIMM_62_AWSIZE,
    output wire [1:0]                      M_AXIMM_62_AWBURST,
    output wire [1:0]                      M_AXIMM_62_AWLOCK,
    output wire [3:0]                      M_AXIMM_62_AWCACHE,
    output wire [2:0]                      M_AXIMM_62_AWPROT,
    output wire [3:0]                      M_AXIMM_62_AWREGION,
    output wire [3:0]                      M_AXIMM_62_AWQOS,
    output wire                            M_AXIMM_62_AWVALID,
    input  wire                            M_AXIMM_62_AWREADY,
    output wire [M_AXIMM_62_DATA_WIDTH-1:0]   M_AXIMM_62_WDATA,
    output wire [M_AXIMM_62_DATA_WIDTH/8-1:0] M_AXIMM_62_WSTRB,
    output wire                            M_AXIMM_62_WLAST,
    output wire                            M_AXIMM_62_WVALID,
    input  wire                            M_AXIMM_62_WREADY,
    input  wire [1:0]                      M_AXIMM_62_BRESP,
    input  wire                            M_AXIMM_62_BVALID,
    output wire                            M_AXIMM_62_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_62_ARADDR,
    output wire [7:0]                      M_AXIMM_62_ARLEN,
    output wire [2:0]                      M_AXIMM_62_ARSIZE,
    output wire [1:0]                      M_AXIMM_62_ARBURST,
    output wire [1:0]                      M_AXIMM_62_ARLOCK,
    output wire [3:0]                      M_AXIMM_62_ARCACHE,
    output wire [2:0]                      M_AXIMM_62_ARPROT,
    output wire [3:0]                      M_AXIMM_62_ARREGION,
    output wire [3:0]                      M_AXIMM_62_ARQOS,
    output wire                            M_AXIMM_62_ARVALID,
    input  wire                            M_AXIMM_62_ARREADY,
    input  wire [M_AXIMM_62_DATA_WIDTH-1:0]   M_AXIMM_62_RDATA,
    input  wire [1:0]                      M_AXIMM_62_RRESP,
    input  wire                            M_AXIMM_62_RLAST,
    input  wire                            M_AXIMM_62_RVALID,
    output wire                            M_AXIMM_62_RREADY,
    //AXI-MM pass-through interface 63
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_63_AWADDR,
    input wire [7:0]                      AP_AXIMM_63_AWLEN,
    input wire [2:0]                      AP_AXIMM_63_AWSIZE,
    input wire [1:0]                      AP_AXIMM_63_AWBURST,
    input wire [1:0]                      AP_AXIMM_63_AWLOCK,
    input wire [3:0]                      AP_AXIMM_63_AWCACHE,
    input wire [2:0]                      AP_AXIMM_63_AWPROT,
    input wire [3:0]                      AP_AXIMM_63_AWREGION,
    input wire [3:0]                      AP_AXIMM_63_AWQOS,
    input wire                            AP_AXIMM_63_AWVALID,
    output  wire                            AP_AXIMM_63_AWREADY,
    input wire [M_AXIMM_63_DATA_WIDTH-1:0]   AP_AXIMM_63_WDATA,
    input wire [M_AXIMM_63_DATA_WIDTH/8-1:0] AP_AXIMM_63_WSTRB,
    input wire                            AP_AXIMM_63_WLAST,
    input wire                            AP_AXIMM_63_WVALID,
    output  wire                            AP_AXIMM_63_WREADY,
    output  wire [1:0]                      AP_AXIMM_63_BRESP,
    output  wire                            AP_AXIMM_63_BVALID,
    input wire                            AP_AXIMM_63_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_63_ARADDR,
    input wire [7:0]                      AP_AXIMM_63_ARLEN,
    input wire [2:0]                      AP_AXIMM_63_ARSIZE,
    input wire [1:0]                      AP_AXIMM_63_ARBURST,
    input wire [1:0]                      AP_AXIMM_63_ARLOCK,
    input wire [3:0]                      AP_AXIMM_63_ARCACHE,
    input wire [2:0]                      AP_AXIMM_63_ARPROT,
    input wire [3:0]                      AP_AXIMM_63_ARREGION,
    input wire [3:0]                      AP_AXIMM_63_ARQOS,
    input wire                            AP_AXIMM_63_ARVALID,
    output  wire                            AP_AXIMM_63_ARREADY,
    output  wire [M_AXIMM_63_DATA_WIDTH-1:0]   AP_AXIMM_63_RDATA,
    output  wire [1:0]                      AP_AXIMM_63_RRESP,
    output  wire                            AP_AXIMM_63_RLAST,
    output  wire                            AP_AXIMM_63_RVALID,
    input  wire                            AP_AXIMM_63_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_63_AWADDR,
    output wire [7:0]                      M_AXIMM_63_AWLEN,
    output wire [2:0]                      M_AXIMM_63_AWSIZE,
    output wire [1:0]                      M_AXIMM_63_AWBURST,
    output wire [1:0]                      M_AXIMM_63_AWLOCK,
    output wire [3:0]                      M_AXIMM_63_AWCACHE,
    output wire [2:0]                      M_AXIMM_63_AWPROT,
    output wire [3:0]                      M_AXIMM_63_AWREGION,
    output wire [3:0]                      M_AXIMM_63_AWQOS,
    output wire                            M_AXIMM_63_AWVALID,
    input  wire                            M_AXIMM_63_AWREADY,
    output wire [M_AXIMM_63_DATA_WIDTH-1:0]   M_AXIMM_63_WDATA,
    output wire [M_AXIMM_63_DATA_WIDTH/8-1:0] M_AXIMM_63_WSTRB,
    output wire                            M_AXIMM_63_WLAST,
    output wire                            M_AXIMM_63_WVALID,
    input  wire                            M_AXIMM_63_WREADY,
    input  wire [1:0]                      M_AXIMM_63_BRESP,
    input  wire                            M_AXIMM_63_BVALID,
    output wire                            M_AXIMM_63_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_63_ARADDR,
    output wire [7:0]                      M_AXIMM_63_ARLEN,
    output wire [2:0]                      M_AXIMM_63_ARSIZE,
    output wire [1:0]                      M_AXIMM_63_ARBURST,
    output wire [1:0]                      M_AXIMM_63_ARLOCK,
    output wire [3:0]                      M_AXIMM_63_ARCACHE,
    output wire [2:0]                      M_AXIMM_63_ARPROT,
    output wire [3:0]                      M_AXIMM_63_ARREGION,
    output wire [3:0]                      M_AXIMM_63_ARQOS,
    output wire                            M_AXIMM_63_ARVALID,
    input  wire                            M_AXIMM_63_ARREADY,
    input  wire [M_AXIMM_63_DATA_WIDTH-1:0]   M_AXIMM_63_RDATA,
    input  wire [1:0]                      M_AXIMM_63_RRESP,
    input  wire                            M_AXIMM_63_RLAST,
    input  wire                            M_AXIMM_63_RVALID,
    output wire                            M_AXIMM_63_RREADY,
    //AXI-MM pass-through interface 64
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_64_AWADDR,
    input wire [7:0]                      AP_AXIMM_64_AWLEN,
    input wire [2:0]                      AP_AXIMM_64_AWSIZE,
    input wire [1:0]                      AP_AXIMM_64_AWBURST,
    input wire [1:0]                      AP_AXIMM_64_AWLOCK,
    input wire [3:0]                      AP_AXIMM_64_AWCACHE,
    input wire [2:0]                      AP_AXIMM_64_AWPROT,
    input wire [3:0]                      AP_AXIMM_64_AWREGION,
    input wire [3:0]                      AP_AXIMM_64_AWQOS,
    input wire                            AP_AXIMM_64_AWVALID,
    output  wire                            AP_AXIMM_64_AWREADY,
    input wire [M_AXIMM_64_DATA_WIDTH-1:0]   AP_AXIMM_64_WDATA,
    input wire [M_AXIMM_64_DATA_WIDTH/8-1:0] AP_AXIMM_64_WSTRB,
    input wire                            AP_AXIMM_64_WLAST,
    input wire                            AP_AXIMM_64_WVALID,
    output  wire                            AP_AXIMM_64_WREADY,
    output  wire [1:0]                      AP_AXIMM_64_BRESP,
    output  wire                            AP_AXIMM_64_BVALID,
    input wire                            AP_AXIMM_64_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_64_ARADDR,
    input wire [7:0]                      AP_AXIMM_64_ARLEN,
    input wire [2:0]                      AP_AXIMM_64_ARSIZE,
    input wire [1:0]                      AP_AXIMM_64_ARBURST,
    input wire [1:0]                      AP_AXIMM_64_ARLOCK,
    input wire [3:0]                      AP_AXIMM_64_ARCACHE,
    input wire [2:0]                      AP_AXIMM_64_ARPROT,
    input wire [3:0]                      AP_AXIMM_64_ARREGION,
    input wire [3:0]                      AP_AXIMM_64_ARQOS,
    input wire                            AP_AXIMM_64_ARVALID,
    output  wire                            AP_AXIMM_64_ARREADY,
    output  wire [M_AXIMM_64_DATA_WIDTH-1:0]   AP_AXIMM_64_RDATA,
    output  wire [1:0]                      AP_AXIMM_64_RRESP,
    output  wire                            AP_AXIMM_64_RLAST,
    output  wire                            AP_AXIMM_64_RVALID,
    input  wire                            AP_AXIMM_64_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_64_AWADDR,
    output wire [7:0]                      M_AXIMM_64_AWLEN,
    output wire [2:0]                      M_AXIMM_64_AWSIZE,
    output wire [1:0]                      M_AXIMM_64_AWBURST,
    output wire [1:0]                      M_AXIMM_64_AWLOCK,
    output wire [3:0]                      M_AXIMM_64_AWCACHE,
    output wire [2:0]                      M_AXIMM_64_AWPROT,
    output wire [3:0]                      M_AXIMM_64_AWREGION,
    output wire [3:0]                      M_AXIMM_64_AWQOS,
    output wire                            M_AXIMM_64_AWVALID,
    input  wire                            M_AXIMM_64_AWREADY,
    output wire [M_AXIMM_64_DATA_WIDTH-1:0]   M_AXIMM_64_WDATA,
    output wire [M_AXIMM_64_DATA_WIDTH/8-1:0] M_AXIMM_64_WSTRB,
    output wire                            M_AXIMM_64_WLAST,
    output wire                            M_AXIMM_64_WVALID,
    input  wire                            M_AXIMM_64_WREADY,
    input  wire [1:0]                      M_AXIMM_64_BRESP,
    input  wire                            M_AXIMM_64_BVALID,
    output wire                            M_AXIMM_64_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_64_ARADDR,
    output wire [7:0]                      M_AXIMM_64_ARLEN,
    output wire [2:0]                      M_AXIMM_64_ARSIZE,
    output wire [1:0]                      M_AXIMM_64_ARBURST,
    output wire [1:0]                      M_AXIMM_64_ARLOCK,
    output wire [3:0]                      M_AXIMM_64_ARCACHE,
    output wire [2:0]                      M_AXIMM_64_ARPROT,
    output wire [3:0]                      M_AXIMM_64_ARREGION,
    output wire [3:0]                      M_AXIMM_64_ARQOS,
    output wire                            M_AXIMM_64_ARVALID,
    input  wire                            M_AXIMM_64_ARREADY,
    input  wire [M_AXIMM_64_DATA_WIDTH-1:0]   M_AXIMM_64_RDATA,
    input  wire [1:0]                      M_AXIMM_64_RRESP,
    input  wire                            M_AXIMM_64_RLAST,
    input  wire                            M_AXIMM_64_RVALID,
    output wire                            M_AXIMM_64_RREADY,
    //AXI-MM pass-through interface 65
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_65_AWADDR,
    input wire [7:0]                      AP_AXIMM_65_AWLEN,
    input wire [2:0]                      AP_AXIMM_65_AWSIZE,
    input wire [1:0]                      AP_AXIMM_65_AWBURST,
    input wire [1:0]                      AP_AXIMM_65_AWLOCK,
    input wire [3:0]                      AP_AXIMM_65_AWCACHE,
    input wire [2:0]                      AP_AXIMM_65_AWPROT,
    input wire [3:0]                      AP_AXIMM_65_AWREGION,
    input wire [3:0]                      AP_AXIMM_65_AWQOS,
    input wire                            AP_AXIMM_65_AWVALID,
    output  wire                            AP_AXIMM_65_AWREADY,
    input wire [M_AXIMM_65_DATA_WIDTH-1:0]   AP_AXIMM_65_WDATA,
    input wire [M_AXIMM_65_DATA_WIDTH/8-1:0] AP_AXIMM_65_WSTRB,
    input wire                            AP_AXIMM_65_WLAST,
    input wire                            AP_AXIMM_65_WVALID,
    output  wire                            AP_AXIMM_65_WREADY,
    output  wire [1:0]                      AP_AXIMM_65_BRESP,
    output  wire                            AP_AXIMM_65_BVALID,
    input wire                            AP_AXIMM_65_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_65_ARADDR,
    input wire [7:0]                      AP_AXIMM_65_ARLEN,
    input wire [2:0]                      AP_AXIMM_65_ARSIZE,
    input wire [1:0]                      AP_AXIMM_65_ARBURST,
    input wire [1:0]                      AP_AXIMM_65_ARLOCK,
    input wire [3:0]                      AP_AXIMM_65_ARCACHE,
    input wire [2:0]                      AP_AXIMM_65_ARPROT,
    input wire [3:0]                      AP_AXIMM_65_ARREGION,
    input wire [3:0]                      AP_AXIMM_65_ARQOS,
    input wire                            AP_AXIMM_65_ARVALID,
    output  wire                            AP_AXIMM_65_ARREADY,
    output  wire [M_AXIMM_65_DATA_WIDTH-1:0]   AP_AXIMM_65_RDATA,
    output  wire [1:0]                      AP_AXIMM_65_RRESP,
    output  wire                            AP_AXIMM_65_RLAST,
    output  wire                            AP_AXIMM_65_RVALID,
    input  wire                            AP_AXIMM_65_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_65_AWADDR,
    output wire [7:0]                      M_AXIMM_65_AWLEN,
    output wire [2:0]                      M_AXIMM_65_AWSIZE,
    output wire [1:0]                      M_AXIMM_65_AWBURST,
    output wire [1:0]                      M_AXIMM_65_AWLOCK,
    output wire [3:0]                      M_AXIMM_65_AWCACHE,
    output wire [2:0]                      M_AXIMM_65_AWPROT,
    output wire [3:0]                      M_AXIMM_65_AWREGION,
    output wire [3:0]                      M_AXIMM_65_AWQOS,
    output wire                            M_AXIMM_65_AWVALID,
    input  wire                            M_AXIMM_65_AWREADY,
    output wire [M_AXIMM_65_DATA_WIDTH-1:0]   M_AXIMM_65_WDATA,
    output wire [M_AXIMM_65_DATA_WIDTH/8-1:0] M_AXIMM_65_WSTRB,
    output wire                            M_AXIMM_65_WLAST,
    output wire                            M_AXIMM_65_WVALID,
    input  wire                            M_AXIMM_65_WREADY,
    input  wire [1:0]                      M_AXIMM_65_BRESP,
    input  wire                            M_AXIMM_65_BVALID,
    output wire                            M_AXIMM_65_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_65_ARADDR,
    output wire [7:0]                      M_AXIMM_65_ARLEN,
    output wire [2:0]                      M_AXIMM_65_ARSIZE,
    output wire [1:0]                      M_AXIMM_65_ARBURST,
    output wire [1:0]                      M_AXIMM_65_ARLOCK,
    output wire [3:0]                      M_AXIMM_65_ARCACHE,
    output wire [2:0]                      M_AXIMM_65_ARPROT,
    output wire [3:0]                      M_AXIMM_65_ARREGION,
    output wire [3:0]                      M_AXIMM_65_ARQOS,
    output wire                            M_AXIMM_65_ARVALID,
    input  wire                            M_AXIMM_65_ARREADY,
    input  wire [M_AXIMM_65_DATA_WIDTH-1:0]   M_AXIMM_65_RDATA,
    input  wire [1:0]                      M_AXIMM_65_RRESP,
    input  wire                            M_AXIMM_65_RLAST,
    input  wire                            M_AXIMM_65_RVALID,
    output wire                            M_AXIMM_65_RREADY,
    //AXI-MM pass-through interface 66
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_66_AWADDR,
    input wire [7:0]                      AP_AXIMM_66_AWLEN,
    input wire [2:0]                      AP_AXIMM_66_AWSIZE,
    input wire [1:0]                      AP_AXIMM_66_AWBURST,
    input wire [1:0]                      AP_AXIMM_66_AWLOCK,
    input wire [3:0]                      AP_AXIMM_66_AWCACHE,
    input wire [2:0]                      AP_AXIMM_66_AWPROT,
    input wire [3:0]                      AP_AXIMM_66_AWREGION,
    input wire [3:0]                      AP_AXIMM_66_AWQOS,
    input wire                            AP_AXIMM_66_AWVALID,
    output  wire                            AP_AXIMM_66_AWREADY,
    input wire [M_AXIMM_66_DATA_WIDTH-1:0]   AP_AXIMM_66_WDATA,
    input wire [M_AXIMM_66_DATA_WIDTH/8-1:0] AP_AXIMM_66_WSTRB,
    input wire                            AP_AXIMM_66_WLAST,
    input wire                            AP_AXIMM_66_WVALID,
    output  wire                            AP_AXIMM_66_WREADY,
    output  wire [1:0]                      AP_AXIMM_66_BRESP,
    output  wire                            AP_AXIMM_66_BVALID,
    input wire                            AP_AXIMM_66_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_66_ARADDR,
    input wire [7:0]                      AP_AXIMM_66_ARLEN,
    input wire [2:0]                      AP_AXIMM_66_ARSIZE,
    input wire [1:0]                      AP_AXIMM_66_ARBURST,
    input wire [1:0]                      AP_AXIMM_66_ARLOCK,
    input wire [3:0]                      AP_AXIMM_66_ARCACHE,
    input wire [2:0]                      AP_AXIMM_66_ARPROT,
    input wire [3:0]                      AP_AXIMM_66_ARREGION,
    input wire [3:0]                      AP_AXIMM_66_ARQOS,
    input wire                            AP_AXIMM_66_ARVALID,
    output  wire                            AP_AXIMM_66_ARREADY,
    output  wire [M_AXIMM_66_DATA_WIDTH-1:0]   AP_AXIMM_66_RDATA,
    output  wire [1:0]                      AP_AXIMM_66_RRESP,
    output  wire                            AP_AXIMM_66_RLAST,
    output  wire                            AP_AXIMM_66_RVALID,
    input  wire                            AP_AXIMM_66_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_66_AWADDR,
    output wire [7:0]                      M_AXIMM_66_AWLEN,
    output wire [2:0]                      M_AXIMM_66_AWSIZE,
    output wire [1:0]                      M_AXIMM_66_AWBURST,
    output wire [1:0]                      M_AXIMM_66_AWLOCK,
    output wire [3:0]                      M_AXIMM_66_AWCACHE,
    output wire [2:0]                      M_AXIMM_66_AWPROT,
    output wire [3:0]                      M_AXIMM_66_AWREGION,
    output wire [3:0]                      M_AXIMM_66_AWQOS,
    output wire                            M_AXIMM_66_AWVALID,
    input  wire                            M_AXIMM_66_AWREADY,
    output wire [M_AXIMM_66_DATA_WIDTH-1:0]   M_AXIMM_66_WDATA,
    output wire [M_AXIMM_66_DATA_WIDTH/8-1:0] M_AXIMM_66_WSTRB,
    output wire                            M_AXIMM_66_WLAST,
    output wire                            M_AXIMM_66_WVALID,
    input  wire                            M_AXIMM_66_WREADY,
    input  wire [1:0]                      M_AXIMM_66_BRESP,
    input  wire                            M_AXIMM_66_BVALID,
    output wire                            M_AXIMM_66_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_66_ARADDR,
    output wire [7:0]                      M_AXIMM_66_ARLEN,
    output wire [2:0]                      M_AXIMM_66_ARSIZE,
    output wire [1:0]                      M_AXIMM_66_ARBURST,
    output wire [1:0]                      M_AXIMM_66_ARLOCK,
    output wire [3:0]                      M_AXIMM_66_ARCACHE,
    output wire [2:0]                      M_AXIMM_66_ARPROT,
    output wire [3:0]                      M_AXIMM_66_ARREGION,
    output wire [3:0]                      M_AXIMM_66_ARQOS,
    output wire                            M_AXIMM_66_ARVALID,
    input  wire                            M_AXIMM_66_ARREADY,
    input  wire [M_AXIMM_66_DATA_WIDTH-1:0]   M_AXIMM_66_RDATA,
    input  wire [1:0]                      M_AXIMM_66_RRESP,
    input  wire                            M_AXIMM_66_RLAST,
    input  wire                            M_AXIMM_66_RVALID,
    output wire                            M_AXIMM_66_RREADY,
    //AXI-MM pass-through interface 67
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_67_AWADDR,
    input wire [7:0]                      AP_AXIMM_67_AWLEN,
    input wire [2:0]                      AP_AXIMM_67_AWSIZE,
    input wire [1:0]                      AP_AXIMM_67_AWBURST,
    input wire [1:0]                      AP_AXIMM_67_AWLOCK,
    input wire [3:0]                      AP_AXIMM_67_AWCACHE,
    input wire [2:0]                      AP_AXIMM_67_AWPROT,
    input wire [3:0]                      AP_AXIMM_67_AWREGION,
    input wire [3:0]                      AP_AXIMM_67_AWQOS,
    input wire                            AP_AXIMM_67_AWVALID,
    output  wire                            AP_AXIMM_67_AWREADY,
    input wire [M_AXIMM_67_DATA_WIDTH-1:0]   AP_AXIMM_67_WDATA,
    input wire [M_AXIMM_67_DATA_WIDTH/8-1:0] AP_AXIMM_67_WSTRB,
    input wire                            AP_AXIMM_67_WLAST,
    input wire                            AP_AXIMM_67_WVALID,
    output  wire                            AP_AXIMM_67_WREADY,
    output  wire [1:0]                      AP_AXIMM_67_BRESP,
    output  wire                            AP_AXIMM_67_BVALID,
    input wire                            AP_AXIMM_67_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_67_ARADDR,
    input wire [7:0]                      AP_AXIMM_67_ARLEN,
    input wire [2:0]                      AP_AXIMM_67_ARSIZE,
    input wire [1:0]                      AP_AXIMM_67_ARBURST,
    input wire [1:0]                      AP_AXIMM_67_ARLOCK,
    input wire [3:0]                      AP_AXIMM_67_ARCACHE,
    input wire [2:0]                      AP_AXIMM_67_ARPROT,
    input wire [3:0]                      AP_AXIMM_67_ARREGION,
    input wire [3:0]                      AP_AXIMM_67_ARQOS,
    input wire                            AP_AXIMM_67_ARVALID,
    output  wire                            AP_AXIMM_67_ARREADY,
    output  wire [M_AXIMM_67_DATA_WIDTH-1:0]   AP_AXIMM_67_RDATA,
    output  wire [1:0]                      AP_AXIMM_67_RRESP,
    output  wire                            AP_AXIMM_67_RLAST,
    output  wire                            AP_AXIMM_67_RVALID,
    input  wire                            AP_AXIMM_67_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_67_AWADDR,
    output wire [7:0]                      M_AXIMM_67_AWLEN,
    output wire [2:0]                      M_AXIMM_67_AWSIZE,
    output wire [1:0]                      M_AXIMM_67_AWBURST,
    output wire [1:0]                      M_AXIMM_67_AWLOCK,
    output wire [3:0]                      M_AXIMM_67_AWCACHE,
    output wire [2:0]                      M_AXIMM_67_AWPROT,
    output wire [3:0]                      M_AXIMM_67_AWREGION,
    output wire [3:0]                      M_AXIMM_67_AWQOS,
    output wire                            M_AXIMM_67_AWVALID,
    input  wire                            M_AXIMM_67_AWREADY,
    output wire [M_AXIMM_67_DATA_WIDTH-1:0]   M_AXIMM_67_WDATA,
    output wire [M_AXIMM_67_DATA_WIDTH/8-1:0] M_AXIMM_67_WSTRB,
    output wire                            M_AXIMM_67_WLAST,
    output wire                            M_AXIMM_67_WVALID,
    input  wire                            M_AXIMM_67_WREADY,
    input  wire [1:0]                      M_AXIMM_67_BRESP,
    input  wire                            M_AXIMM_67_BVALID,
    output wire                            M_AXIMM_67_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_67_ARADDR,
    output wire [7:0]                      M_AXIMM_67_ARLEN,
    output wire [2:0]                      M_AXIMM_67_ARSIZE,
    output wire [1:0]                      M_AXIMM_67_ARBURST,
    output wire [1:0]                      M_AXIMM_67_ARLOCK,
    output wire [3:0]                      M_AXIMM_67_ARCACHE,
    output wire [2:0]                      M_AXIMM_67_ARPROT,
    output wire [3:0]                      M_AXIMM_67_ARREGION,
    output wire [3:0]                      M_AXIMM_67_ARQOS,
    output wire                            M_AXIMM_67_ARVALID,
    input  wire                            M_AXIMM_67_ARREADY,
    input  wire [M_AXIMM_67_DATA_WIDTH-1:0]   M_AXIMM_67_RDATA,
    input  wire [1:0]                      M_AXIMM_67_RRESP,
    input  wire                            M_AXIMM_67_RLAST,
    input  wire                            M_AXIMM_67_RVALID,
    output wire                            M_AXIMM_67_RREADY,
    //AXI-MM pass-through interface 68
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_68_AWADDR,
    input wire [7:0]                      AP_AXIMM_68_AWLEN,
    input wire [2:0]                      AP_AXIMM_68_AWSIZE,
    input wire [1:0]                      AP_AXIMM_68_AWBURST,
    input wire [1:0]                      AP_AXIMM_68_AWLOCK,
    input wire [3:0]                      AP_AXIMM_68_AWCACHE,
    input wire [2:0]                      AP_AXIMM_68_AWPROT,
    input wire [3:0]                      AP_AXIMM_68_AWREGION,
    input wire [3:0]                      AP_AXIMM_68_AWQOS,
    input wire                            AP_AXIMM_68_AWVALID,
    output  wire                            AP_AXIMM_68_AWREADY,
    input wire [M_AXIMM_68_DATA_WIDTH-1:0]   AP_AXIMM_68_WDATA,
    input wire [M_AXIMM_68_DATA_WIDTH/8-1:0] AP_AXIMM_68_WSTRB,
    input wire                            AP_AXIMM_68_WLAST,
    input wire                            AP_AXIMM_68_WVALID,
    output  wire                            AP_AXIMM_68_WREADY,
    output  wire [1:0]                      AP_AXIMM_68_BRESP,
    output  wire                            AP_AXIMM_68_BVALID,
    input wire                            AP_AXIMM_68_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_68_ARADDR,
    input wire [7:0]                      AP_AXIMM_68_ARLEN,
    input wire [2:0]                      AP_AXIMM_68_ARSIZE,
    input wire [1:0]                      AP_AXIMM_68_ARBURST,
    input wire [1:0]                      AP_AXIMM_68_ARLOCK,
    input wire [3:0]                      AP_AXIMM_68_ARCACHE,
    input wire [2:0]                      AP_AXIMM_68_ARPROT,
    input wire [3:0]                      AP_AXIMM_68_ARREGION,
    input wire [3:0]                      AP_AXIMM_68_ARQOS,
    input wire                            AP_AXIMM_68_ARVALID,
    output  wire                            AP_AXIMM_68_ARREADY,
    output  wire [M_AXIMM_68_DATA_WIDTH-1:0]   AP_AXIMM_68_RDATA,
    output  wire [1:0]                      AP_AXIMM_68_RRESP,
    output  wire                            AP_AXIMM_68_RLAST,
    output  wire                            AP_AXIMM_68_RVALID,
    input  wire                            AP_AXIMM_68_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_68_AWADDR,
    output wire [7:0]                      M_AXIMM_68_AWLEN,
    output wire [2:0]                      M_AXIMM_68_AWSIZE,
    output wire [1:0]                      M_AXIMM_68_AWBURST,
    output wire [1:0]                      M_AXIMM_68_AWLOCK,
    output wire [3:0]                      M_AXIMM_68_AWCACHE,
    output wire [2:0]                      M_AXIMM_68_AWPROT,
    output wire [3:0]                      M_AXIMM_68_AWREGION,
    output wire [3:0]                      M_AXIMM_68_AWQOS,
    output wire                            M_AXIMM_68_AWVALID,
    input  wire                            M_AXIMM_68_AWREADY,
    output wire [M_AXIMM_68_DATA_WIDTH-1:0]   M_AXIMM_68_WDATA,
    output wire [M_AXIMM_68_DATA_WIDTH/8-1:0] M_AXIMM_68_WSTRB,
    output wire                            M_AXIMM_68_WLAST,
    output wire                            M_AXIMM_68_WVALID,
    input  wire                            M_AXIMM_68_WREADY,
    input  wire [1:0]                      M_AXIMM_68_BRESP,
    input  wire                            M_AXIMM_68_BVALID,
    output wire                            M_AXIMM_68_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_68_ARADDR,
    output wire [7:0]                      M_AXIMM_68_ARLEN,
    output wire [2:0]                      M_AXIMM_68_ARSIZE,
    output wire [1:0]                      M_AXIMM_68_ARBURST,
    output wire [1:0]                      M_AXIMM_68_ARLOCK,
    output wire [3:0]                      M_AXIMM_68_ARCACHE,
    output wire [2:0]                      M_AXIMM_68_ARPROT,
    output wire [3:0]                      M_AXIMM_68_ARREGION,
    output wire [3:0]                      M_AXIMM_68_ARQOS,
    output wire                            M_AXIMM_68_ARVALID,
    input  wire                            M_AXIMM_68_ARREADY,
    input  wire [M_AXIMM_68_DATA_WIDTH-1:0]   M_AXIMM_68_RDATA,
    input  wire [1:0]                      M_AXIMM_68_RRESP,
    input  wire                            M_AXIMM_68_RLAST,
    input  wire                            M_AXIMM_68_RVALID,
    output wire                            M_AXIMM_68_RREADY,
    //AXI-MM pass-through interface 69
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_69_AWADDR,
    input wire [7:0]                      AP_AXIMM_69_AWLEN,
    input wire [2:0]                      AP_AXIMM_69_AWSIZE,
    input wire [1:0]                      AP_AXIMM_69_AWBURST,
    input wire [1:0]                      AP_AXIMM_69_AWLOCK,
    input wire [3:0]                      AP_AXIMM_69_AWCACHE,
    input wire [2:0]                      AP_AXIMM_69_AWPROT,
    input wire [3:0]                      AP_AXIMM_69_AWREGION,
    input wire [3:0]                      AP_AXIMM_69_AWQOS,
    input wire                            AP_AXIMM_69_AWVALID,
    output  wire                            AP_AXIMM_69_AWREADY,
    input wire [M_AXIMM_69_DATA_WIDTH-1:0]   AP_AXIMM_69_WDATA,
    input wire [M_AXIMM_69_DATA_WIDTH/8-1:0] AP_AXIMM_69_WSTRB,
    input wire                            AP_AXIMM_69_WLAST,
    input wire                            AP_AXIMM_69_WVALID,
    output  wire                            AP_AXIMM_69_WREADY,
    output  wire [1:0]                      AP_AXIMM_69_BRESP,
    output  wire                            AP_AXIMM_69_BVALID,
    input wire                            AP_AXIMM_69_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_69_ARADDR,
    input wire [7:0]                      AP_AXIMM_69_ARLEN,
    input wire [2:0]                      AP_AXIMM_69_ARSIZE,
    input wire [1:0]                      AP_AXIMM_69_ARBURST,
    input wire [1:0]                      AP_AXIMM_69_ARLOCK,
    input wire [3:0]                      AP_AXIMM_69_ARCACHE,
    input wire [2:0]                      AP_AXIMM_69_ARPROT,
    input wire [3:0]                      AP_AXIMM_69_ARREGION,
    input wire [3:0]                      AP_AXIMM_69_ARQOS,
    input wire                            AP_AXIMM_69_ARVALID,
    output  wire                            AP_AXIMM_69_ARREADY,
    output  wire [M_AXIMM_69_DATA_WIDTH-1:0]   AP_AXIMM_69_RDATA,
    output  wire [1:0]                      AP_AXIMM_69_RRESP,
    output  wire                            AP_AXIMM_69_RLAST,
    output  wire                            AP_AXIMM_69_RVALID,
    input  wire                            AP_AXIMM_69_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_69_AWADDR,
    output wire [7:0]                      M_AXIMM_69_AWLEN,
    output wire [2:0]                      M_AXIMM_69_AWSIZE,
    output wire [1:0]                      M_AXIMM_69_AWBURST,
    output wire [1:0]                      M_AXIMM_69_AWLOCK,
    output wire [3:0]                      M_AXIMM_69_AWCACHE,
    output wire [2:0]                      M_AXIMM_69_AWPROT,
    output wire [3:0]                      M_AXIMM_69_AWREGION,
    output wire [3:0]                      M_AXIMM_69_AWQOS,
    output wire                            M_AXIMM_69_AWVALID,
    input  wire                            M_AXIMM_69_AWREADY,
    output wire [M_AXIMM_69_DATA_WIDTH-1:0]   M_AXIMM_69_WDATA,
    output wire [M_AXIMM_69_DATA_WIDTH/8-1:0] M_AXIMM_69_WSTRB,
    output wire                            M_AXIMM_69_WLAST,
    output wire                            M_AXIMM_69_WVALID,
    input  wire                            M_AXIMM_69_WREADY,
    input  wire [1:0]                      M_AXIMM_69_BRESP,
    input  wire                            M_AXIMM_69_BVALID,
    output wire                            M_AXIMM_69_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_69_ARADDR,
    output wire [7:0]                      M_AXIMM_69_ARLEN,
    output wire [2:0]                      M_AXIMM_69_ARSIZE,
    output wire [1:0]                      M_AXIMM_69_ARBURST,
    output wire [1:0]                      M_AXIMM_69_ARLOCK,
    output wire [3:0]                      M_AXIMM_69_ARCACHE,
    output wire [2:0]                      M_AXIMM_69_ARPROT,
    output wire [3:0]                      M_AXIMM_69_ARREGION,
    output wire [3:0]                      M_AXIMM_69_ARQOS,
    output wire                            M_AXIMM_69_ARVALID,
    input  wire                            M_AXIMM_69_ARREADY,
    input  wire [M_AXIMM_69_DATA_WIDTH-1:0]   M_AXIMM_69_RDATA,
    input  wire [1:0]                      M_AXIMM_69_RRESP,
    input  wire                            M_AXIMM_69_RLAST,
    input  wire                            M_AXIMM_69_RVALID,
    output wire                            M_AXIMM_69_RREADY,
    //AXI-MM pass-through interface 70
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_70_AWADDR,
    input wire [7:0]                      AP_AXIMM_70_AWLEN,
    input wire [2:0]                      AP_AXIMM_70_AWSIZE,
    input wire [1:0]                      AP_AXIMM_70_AWBURST,
    input wire [1:0]                      AP_AXIMM_70_AWLOCK,
    input wire [3:0]                      AP_AXIMM_70_AWCACHE,
    input wire [2:0]                      AP_AXIMM_70_AWPROT,
    input wire [3:0]                      AP_AXIMM_70_AWREGION,
    input wire [3:0]                      AP_AXIMM_70_AWQOS,
    input wire                            AP_AXIMM_70_AWVALID,
    output  wire                            AP_AXIMM_70_AWREADY,
    input wire [M_AXIMM_70_DATA_WIDTH-1:0]   AP_AXIMM_70_WDATA,
    input wire [M_AXIMM_70_DATA_WIDTH/8-1:0] AP_AXIMM_70_WSTRB,
    input wire                            AP_AXIMM_70_WLAST,
    input wire                            AP_AXIMM_70_WVALID,
    output  wire                            AP_AXIMM_70_WREADY,
    output  wire [1:0]                      AP_AXIMM_70_BRESP,
    output  wire                            AP_AXIMM_70_BVALID,
    input wire                            AP_AXIMM_70_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_70_ARADDR,
    input wire [7:0]                      AP_AXIMM_70_ARLEN,
    input wire [2:0]                      AP_AXIMM_70_ARSIZE,
    input wire [1:0]                      AP_AXIMM_70_ARBURST,
    input wire [1:0]                      AP_AXIMM_70_ARLOCK,
    input wire [3:0]                      AP_AXIMM_70_ARCACHE,
    input wire [2:0]                      AP_AXIMM_70_ARPROT,
    input wire [3:0]                      AP_AXIMM_70_ARREGION,
    input wire [3:0]                      AP_AXIMM_70_ARQOS,
    input wire                            AP_AXIMM_70_ARVALID,
    output  wire                            AP_AXIMM_70_ARREADY,
    output  wire [M_AXIMM_70_DATA_WIDTH-1:0]   AP_AXIMM_70_RDATA,
    output  wire [1:0]                      AP_AXIMM_70_RRESP,
    output  wire                            AP_AXIMM_70_RLAST,
    output  wire                            AP_AXIMM_70_RVALID,
    input  wire                            AP_AXIMM_70_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_70_AWADDR,
    output wire [7:0]                      M_AXIMM_70_AWLEN,
    output wire [2:0]                      M_AXIMM_70_AWSIZE,
    output wire [1:0]                      M_AXIMM_70_AWBURST,
    output wire [1:0]                      M_AXIMM_70_AWLOCK,
    output wire [3:0]                      M_AXIMM_70_AWCACHE,
    output wire [2:0]                      M_AXIMM_70_AWPROT,
    output wire [3:0]                      M_AXIMM_70_AWREGION,
    output wire [3:0]                      M_AXIMM_70_AWQOS,
    output wire                            M_AXIMM_70_AWVALID,
    input  wire                            M_AXIMM_70_AWREADY,
    output wire [M_AXIMM_70_DATA_WIDTH-1:0]   M_AXIMM_70_WDATA,
    output wire [M_AXIMM_70_DATA_WIDTH/8-1:0] M_AXIMM_70_WSTRB,
    output wire                            M_AXIMM_70_WLAST,
    output wire                            M_AXIMM_70_WVALID,
    input  wire                            M_AXIMM_70_WREADY,
    input  wire [1:0]                      M_AXIMM_70_BRESP,
    input  wire                            M_AXIMM_70_BVALID,
    output wire                            M_AXIMM_70_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_70_ARADDR,
    output wire [7:0]                      M_AXIMM_70_ARLEN,
    output wire [2:0]                      M_AXIMM_70_ARSIZE,
    output wire [1:0]                      M_AXIMM_70_ARBURST,
    output wire [1:0]                      M_AXIMM_70_ARLOCK,
    output wire [3:0]                      M_AXIMM_70_ARCACHE,
    output wire [2:0]                      M_AXIMM_70_ARPROT,
    output wire [3:0]                      M_AXIMM_70_ARREGION,
    output wire [3:0]                      M_AXIMM_70_ARQOS,
    output wire                            M_AXIMM_70_ARVALID,
    input  wire                            M_AXIMM_70_ARREADY,
    input  wire [M_AXIMM_70_DATA_WIDTH-1:0]   M_AXIMM_70_RDATA,
    input  wire [1:0]                      M_AXIMM_70_RRESP,
    input  wire                            M_AXIMM_70_RLAST,
    input  wire                            M_AXIMM_70_RVALID,
    output wire                            M_AXIMM_70_RREADY,
    //AXI-MM pass-through interface 71
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_71_AWADDR,
    input wire [7:0]                      AP_AXIMM_71_AWLEN,
    input wire [2:0]                      AP_AXIMM_71_AWSIZE,
    input wire [1:0]                      AP_AXIMM_71_AWBURST,
    input wire [1:0]                      AP_AXIMM_71_AWLOCK,
    input wire [3:0]                      AP_AXIMM_71_AWCACHE,
    input wire [2:0]                      AP_AXIMM_71_AWPROT,
    input wire [3:0]                      AP_AXIMM_71_AWREGION,
    input wire [3:0]                      AP_AXIMM_71_AWQOS,
    input wire                            AP_AXIMM_71_AWVALID,
    output  wire                            AP_AXIMM_71_AWREADY,
    input wire [M_AXIMM_71_DATA_WIDTH-1:0]   AP_AXIMM_71_WDATA,
    input wire [M_AXIMM_71_DATA_WIDTH/8-1:0] AP_AXIMM_71_WSTRB,
    input wire                            AP_AXIMM_71_WLAST,
    input wire                            AP_AXIMM_71_WVALID,
    output  wire                            AP_AXIMM_71_WREADY,
    output  wire [1:0]                      AP_AXIMM_71_BRESP,
    output  wire                            AP_AXIMM_71_BVALID,
    input wire                            AP_AXIMM_71_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_71_ARADDR,
    input wire [7:0]                      AP_AXIMM_71_ARLEN,
    input wire [2:0]                      AP_AXIMM_71_ARSIZE,
    input wire [1:0]                      AP_AXIMM_71_ARBURST,
    input wire [1:0]                      AP_AXIMM_71_ARLOCK,
    input wire [3:0]                      AP_AXIMM_71_ARCACHE,
    input wire [2:0]                      AP_AXIMM_71_ARPROT,
    input wire [3:0]                      AP_AXIMM_71_ARREGION,
    input wire [3:0]                      AP_AXIMM_71_ARQOS,
    input wire                            AP_AXIMM_71_ARVALID,
    output  wire                            AP_AXIMM_71_ARREADY,
    output  wire [M_AXIMM_71_DATA_WIDTH-1:0]   AP_AXIMM_71_RDATA,
    output  wire [1:0]                      AP_AXIMM_71_RRESP,
    output  wire                            AP_AXIMM_71_RLAST,
    output  wire                            AP_AXIMM_71_RVALID,
    input  wire                            AP_AXIMM_71_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_71_AWADDR,
    output wire [7:0]                      M_AXIMM_71_AWLEN,
    output wire [2:0]                      M_AXIMM_71_AWSIZE,
    output wire [1:0]                      M_AXIMM_71_AWBURST,
    output wire [1:0]                      M_AXIMM_71_AWLOCK,
    output wire [3:0]                      M_AXIMM_71_AWCACHE,
    output wire [2:0]                      M_AXIMM_71_AWPROT,
    output wire [3:0]                      M_AXIMM_71_AWREGION,
    output wire [3:0]                      M_AXIMM_71_AWQOS,
    output wire                            M_AXIMM_71_AWVALID,
    input  wire                            M_AXIMM_71_AWREADY,
    output wire [M_AXIMM_71_DATA_WIDTH-1:0]   M_AXIMM_71_WDATA,
    output wire [M_AXIMM_71_DATA_WIDTH/8-1:0] M_AXIMM_71_WSTRB,
    output wire                            M_AXIMM_71_WLAST,
    output wire                            M_AXIMM_71_WVALID,
    input  wire                            M_AXIMM_71_WREADY,
    input  wire [1:0]                      M_AXIMM_71_BRESP,
    input  wire                            M_AXIMM_71_BVALID,
    output wire                            M_AXIMM_71_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_71_ARADDR,
    output wire [7:0]                      M_AXIMM_71_ARLEN,
    output wire [2:0]                      M_AXIMM_71_ARSIZE,
    output wire [1:0]                      M_AXIMM_71_ARBURST,
    output wire [1:0]                      M_AXIMM_71_ARLOCK,
    output wire [3:0]                      M_AXIMM_71_ARCACHE,
    output wire [2:0]                      M_AXIMM_71_ARPROT,
    output wire [3:0]                      M_AXIMM_71_ARREGION,
    output wire [3:0]                      M_AXIMM_71_ARQOS,
    output wire                            M_AXIMM_71_ARVALID,
    input  wire                            M_AXIMM_71_ARREADY,
    input  wire [M_AXIMM_71_DATA_WIDTH-1:0]   M_AXIMM_71_RDATA,
    input  wire [1:0]                      M_AXIMM_71_RRESP,
    input  wire                            M_AXIMM_71_RLAST,
    input  wire                            M_AXIMM_71_RVALID,
    output wire                            M_AXIMM_71_RREADY,
    //AXI-MM pass-through interface 72
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_72_AWADDR,
    input wire [7:0]                      AP_AXIMM_72_AWLEN,
    input wire [2:0]                      AP_AXIMM_72_AWSIZE,
    input wire [1:0]                      AP_AXIMM_72_AWBURST,
    input wire [1:0]                      AP_AXIMM_72_AWLOCK,
    input wire [3:0]                      AP_AXIMM_72_AWCACHE,
    input wire [2:0]                      AP_AXIMM_72_AWPROT,
    input wire [3:0]                      AP_AXIMM_72_AWREGION,
    input wire [3:0]                      AP_AXIMM_72_AWQOS,
    input wire                            AP_AXIMM_72_AWVALID,
    output  wire                            AP_AXIMM_72_AWREADY,
    input wire [M_AXIMM_72_DATA_WIDTH-1:0]   AP_AXIMM_72_WDATA,
    input wire [M_AXIMM_72_DATA_WIDTH/8-1:0] AP_AXIMM_72_WSTRB,
    input wire                            AP_AXIMM_72_WLAST,
    input wire                            AP_AXIMM_72_WVALID,
    output  wire                            AP_AXIMM_72_WREADY,
    output  wire [1:0]                      AP_AXIMM_72_BRESP,
    output  wire                            AP_AXIMM_72_BVALID,
    input wire                            AP_AXIMM_72_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_72_ARADDR,
    input wire [7:0]                      AP_AXIMM_72_ARLEN,
    input wire [2:0]                      AP_AXIMM_72_ARSIZE,
    input wire [1:0]                      AP_AXIMM_72_ARBURST,
    input wire [1:0]                      AP_AXIMM_72_ARLOCK,
    input wire [3:0]                      AP_AXIMM_72_ARCACHE,
    input wire [2:0]                      AP_AXIMM_72_ARPROT,
    input wire [3:0]                      AP_AXIMM_72_ARREGION,
    input wire [3:0]                      AP_AXIMM_72_ARQOS,
    input wire                            AP_AXIMM_72_ARVALID,
    output  wire                            AP_AXIMM_72_ARREADY,
    output  wire [M_AXIMM_72_DATA_WIDTH-1:0]   AP_AXIMM_72_RDATA,
    output  wire [1:0]                      AP_AXIMM_72_RRESP,
    output  wire                            AP_AXIMM_72_RLAST,
    output  wire                            AP_AXIMM_72_RVALID,
    input  wire                            AP_AXIMM_72_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_72_AWADDR,
    output wire [7:0]                      M_AXIMM_72_AWLEN,
    output wire [2:0]                      M_AXIMM_72_AWSIZE,
    output wire [1:0]                      M_AXIMM_72_AWBURST,
    output wire [1:0]                      M_AXIMM_72_AWLOCK,
    output wire [3:0]                      M_AXIMM_72_AWCACHE,
    output wire [2:0]                      M_AXIMM_72_AWPROT,
    output wire [3:0]                      M_AXIMM_72_AWREGION,
    output wire [3:0]                      M_AXIMM_72_AWQOS,
    output wire                            M_AXIMM_72_AWVALID,
    input  wire                            M_AXIMM_72_AWREADY,
    output wire [M_AXIMM_72_DATA_WIDTH-1:0]   M_AXIMM_72_WDATA,
    output wire [M_AXIMM_72_DATA_WIDTH/8-1:0] M_AXIMM_72_WSTRB,
    output wire                            M_AXIMM_72_WLAST,
    output wire                            M_AXIMM_72_WVALID,
    input  wire                            M_AXIMM_72_WREADY,
    input  wire [1:0]                      M_AXIMM_72_BRESP,
    input  wire                            M_AXIMM_72_BVALID,
    output wire                            M_AXIMM_72_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_72_ARADDR,
    output wire [7:0]                      M_AXIMM_72_ARLEN,
    output wire [2:0]                      M_AXIMM_72_ARSIZE,
    output wire [1:0]                      M_AXIMM_72_ARBURST,
    output wire [1:0]                      M_AXIMM_72_ARLOCK,
    output wire [3:0]                      M_AXIMM_72_ARCACHE,
    output wire [2:0]                      M_AXIMM_72_ARPROT,
    output wire [3:0]                      M_AXIMM_72_ARREGION,
    output wire [3:0]                      M_AXIMM_72_ARQOS,
    output wire                            M_AXIMM_72_ARVALID,
    input  wire                            M_AXIMM_72_ARREADY,
    input  wire [M_AXIMM_72_DATA_WIDTH-1:0]   M_AXIMM_72_RDATA,
    input  wire [1:0]                      M_AXIMM_72_RRESP,
    input  wire                            M_AXIMM_72_RLAST,
    input  wire                            M_AXIMM_72_RVALID,
    output wire                            M_AXIMM_72_RREADY,
    //AXI-MM pass-through interface 73
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_73_AWADDR,
    input wire [7:0]                      AP_AXIMM_73_AWLEN,
    input wire [2:0]                      AP_AXIMM_73_AWSIZE,
    input wire [1:0]                      AP_AXIMM_73_AWBURST,
    input wire [1:0]                      AP_AXIMM_73_AWLOCK,
    input wire [3:0]                      AP_AXIMM_73_AWCACHE,
    input wire [2:0]                      AP_AXIMM_73_AWPROT,
    input wire [3:0]                      AP_AXIMM_73_AWREGION,
    input wire [3:0]                      AP_AXIMM_73_AWQOS,
    input wire                            AP_AXIMM_73_AWVALID,
    output  wire                            AP_AXIMM_73_AWREADY,
    input wire [M_AXIMM_73_DATA_WIDTH-1:0]   AP_AXIMM_73_WDATA,
    input wire [M_AXIMM_73_DATA_WIDTH/8-1:0] AP_AXIMM_73_WSTRB,
    input wire                            AP_AXIMM_73_WLAST,
    input wire                            AP_AXIMM_73_WVALID,
    output  wire                            AP_AXIMM_73_WREADY,
    output  wire [1:0]                      AP_AXIMM_73_BRESP,
    output  wire                            AP_AXIMM_73_BVALID,
    input wire                            AP_AXIMM_73_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_73_ARADDR,
    input wire [7:0]                      AP_AXIMM_73_ARLEN,
    input wire [2:0]                      AP_AXIMM_73_ARSIZE,
    input wire [1:0]                      AP_AXIMM_73_ARBURST,
    input wire [1:0]                      AP_AXIMM_73_ARLOCK,
    input wire [3:0]                      AP_AXIMM_73_ARCACHE,
    input wire [2:0]                      AP_AXIMM_73_ARPROT,
    input wire [3:0]                      AP_AXIMM_73_ARREGION,
    input wire [3:0]                      AP_AXIMM_73_ARQOS,
    input wire                            AP_AXIMM_73_ARVALID,
    output  wire                            AP_AXIMM_73_ARREADY,
    output  wire [M_AXIMM_73_DATA_WIDTH-1:0]   AP_AXIMM_73_RDATA,
    output  wire [1:0]                      AP_AXIMM_73_RRESP,
    output  wire                            AP_AXIMM_73_RLAST,
    output  wire                            AP_AXIMM_73_RVALID,
    input  wire                            AP_AXIMM_73_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_73_AWADDR,
    output wire [7:0]                      M_AXIMM_73_AWLEN,
    output wire [2:0]                      M_AXIMM_73_AWSIZE,
    output wire [1:0]                      M_AXIMM_73_AWBURST,
    output wire [1:0]                      M_AXIMM_73_AWLOCK,
    output wire [3:0]                      M_AXIMM_73_AWCACHE,
    output wire [2:0]                      M_AXIMM_73_AWPROT,
    output wire [3:0]                      M_AXIMM_73_AWREGION,
    output wire [3:0]                      M_AXIMM_73_AWQOS,
    output wire                            M_AXIMM_73_AWVALID,
    input  wire                            M_AXIMM_73_AWREADY,
    output wire [M_AXIMM_73_DATA_WIDTH-1:0]   M_AXIMM_73_WDATA,
    output wire [M_AXIMM_73_DATA_WIDTH/8-1:0] M_AXIMM_73_WSTRB,
    output wire                            M_AXIMM_73_WLAST,
    output wire                            M_AXIMM_73_WVALID,
    input  wire                            M_AXIMM_73_WREADY,
    input  wire [1:0]                      M_AXIMM_73_BRESP,
    input  wire                            M_AXIMM_73_BVALID,
    output wire                            M_AXIMM_73_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_73_ARADDR,
    output wire [7:0]                      M_AXIMM_73_ARLEN,
    output wire [2:0]                      M_AXIMM_73_ARSIZE,
    output wire [1:0]                      M_AXIMM_73_ARBURST,
    output wire [1:0]                      M_AXIMM_73_ARLOCK,
    output wire [3:0]                      M_AXIMM_73_ARCACHE,
    output wire [2:0]                      M_AXIMM_73_ARPROT,
    output wire [3:0]                      M_AXIMM_73_ARREGION,
    output wire [3:0]                      M_AXIMM_73_ARQOS,
    output wire                            M_AXIMM_73_ARVALID,
    input  wire                            M_AXIMM_73_ARREADY,
    input  wire [M_AXIMM_73_DATA_WIDTH-1:0]   M_AXIMM_73_RDATA,
    input  wire [1:0]                      M_AXIMM_73_RRESP,
    input  wire                            M_AXIMM_73_RLAST,
    input  wire                            M_AXIMM_73_RVALID,
    output wire                            M_AXIMM_73_RREADY,
    //AXI-MM pass-through interface 74
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_74_AWADDR,
    input wire [7:0]                      AP_AXIMM_74_AWLEN,
    input wire [2:0]                      AP_AXIMM_74_AWSIZE,
    input wire [1:0]                      AP_AXIMM_74_AWBURST,
    input wire [1:0]                      AP_AXIMM_74_AWLOCK,
    input wire [3:0]                      AP_AXIMM_74_AWCACHE,
    input wire [2:0]                      AP_AXIMM_74_AWPROT,
    input wire [3:0]                      AP_AXIMM_74_AWREGION,
    input wire [3:0]                      AP_AXIMM_74_AWQOS,
    input wire                            AP_AXIMM_74_AWVALID,
    output  wire                            AP_AXIMM_74_AWREADY,
    input wire [M_AXIMM_74_DATA_WIDTH-1:0]   AP_AXIMM_74_WDATA,
    input wire [M_AXIMM_74_DATA_WIDTH/8-1:0] AP_AXIMM_74_WSTRB,
    input wire                            AP_AXIMM_74_WLAST,
    input wire                            AP_AXIMM_74_WVALID,
    output  wire                            AP_AXIMM_74_WREADY,
    output  wire [1:0]                      AP_AXIMM_74_BRESP,
    output  wire                            AP_AXIMM_74_BVALID,
    input wire                            AP_AXIMM_74_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_74_ARADDR,
    input wire [7:0]                      AP_AXIMM_74_ARLEN,
    input wire [2:0]                      AP_AXIMM_74_ARSIZE,
    input wire [1:0]                      AP_AXIMM_74_ARBURST,
    input wire [1:0]                      AP_AXIMM_74_ARLOCK,
    input wire [3:0]                      AP_AXIMM_74_ARCACHE,
    input wire [2:0]                      AP_AXIMM_74_ARPROT,
    input wire [3:0]                      AP_AXIMM_74_ARREGION,
    input wire [3:0]                      AP_AXIMM_74_ARQOS,
    input wire                            AP_AXIMM_74_ARVALID,
    output  wire                            AP_AXIMM_74_ARREADY,
    output  wire [M_AXIMM_74_DATA_WIDTH-1:0]   AP_AXIMM_74_RDATA,
    output  wire [1:0]                      AP_AXIMM_74_RRESP,
    output  wire                            AP_AXIMM_74_RLAST,
    output  wire                            AP_AXIMM_74_RVALID,
    input  wire                            AP_AXIMM_74_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_74_AWADDR,
    output wire [7:0]                      M_AXIMM_74_AWLEN,
    output wire [2:0]                      M_AXIMM_74_AWSIZE,
    output wire [1:0]                      M_AXIMM_74_AWBURST,
    output wire [1:0]                      M_AXIMM_74_AWLOCK,
    output wire [3:0]                      M_AXIMM_74_AWCACHE,
    output wire [2:0]                      M_AXIMM_74_AWPROT,
    output wire [3:0]                      M_AXIMM_74_AWREGION,
    output wire [3:0]                      M_AXIMM_74_AWQOS,
    output wire                            M_AXIMM_74_AWVALID,
    input  wire                            M_AXIMM_74_AWREADY,
    output wire [M_AXIMM_74_DATA_WIDTH-1:0]   M_AXIMM_74_WDATA,
    output wire [M_AXIMM_74_DATA_WIDTH/8-1:0] M_AXIMM_74_WSTRB,
    output wire                            M_AXIMM_74_WLAST,
    output wire                            M_AXIMM_74_WVALID,
    input  wire                            M_AXIMM_74_WREADY,
    input  wire [1:0]                      M_AXIMM_74_BRESP,
    input  wire                            M_AXIMM_74_BVALID,
    output wire                            M_AXIMM_74_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_74_ARADDR,
    output wire [7:0]                      M_AXIMM_74_ARLEN,
    output wire [2:0]                      M_AXIMM_74_ARSIZE,
    output wire [1:0]                      M_AXIMM_74_ARBURST,
    output wire [1:0]                      M_AXIMM_74_ARLOCK,
    output wire [3:0]                      M_AXIMM_74_ARCACHE,
    output wire [2:0]                      M_AXIMM_74_ARPROT,
    output wire [3:0]                      M_AXIMM_74_ARREGION,
    output wire [3:0]                      M_AXIMM_74_ARQOS,
    output wire                            M_AXIMM_74_ARVALID,
    input  wire                            M_AXIMM_74_ARREADY,
    input  wire [M_AXIMM_74_DATA_WIDTH-1:0]   M_AXIMM_74_RDATA,
    input  wire [1:0]                      M_AXIMM_74_RRESP,
    input  wire                            M_AXIMM_74_RLAST,
    input  wire                            M_AXIMM_74_RVALID,
    output wire                            M_AXIMM_74_RREADY,
    //AXI-MM pass-through interface 75
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_75_AWADDR,
    input wire [7:0]                      AP_AXIMM_75_AWLEN,
    input wire [2:0]                      AP_AXIMM_75_AWSIZE,
    input wire [1:0]                      AP_AXIMM_75_AWBURST,
    input wire [1:0]                      AP_AXIMM_75_AWLOCK,
    input wire [3:0]                      AP_AXIMM_75_AWCACHE,
    input wire [2:0]                      AP_AXIMM_75_AWPROT,
    input wire [3:0]                      AP_AXIMM_75_AWREGION,
    input wire [3:0]                      AP_AXIMM_75_AWQOS,
    input wire                            AP_AXIMM_75_AWVALID,
    output  wire                            AP_AXIMM_75_AWREADY,
    input wire [M_AXIMM_75_DATA_WIDTH-1:0]   AP_AXIMM_75_WDATA,
    input wire [M_AXIMM_75_DATA_WIDTH/8-1:0] AP_AXIMM_75_WSTRB,
    input wire                            AP_AXIMM_75_WLAST,
    input wire                            AP_AXIMM_75_WVALID,
    output  wire                            AP_AXIMM_75_WREADY,
    output  wire [1:0]                      AP_AXIMM_75_BRESP,
    output  wire                            AP_AXIMM_75_BVALID,
    input wire                            AP_AXIMM_75_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_75_ARADDR,
    input wire [7:0]                      AP_AXIMM_75_ARLEN,
    input wire [2:0]                      AP_AXIMM_75_ARSIZE,
    input wire [1:0]                      AP_AXIMM_75_ARBURST,
    input wire [1:0]                      AP_AXIMM_75_ARLOCK,
    input wire [3:0]                      AP_AXIMM_75_ARCACHE,
    input wire [2:0]                      AP_AXIMM_75_ARPROT,
    input wire [3:0]                      AP_AXIMM_75_ARREGION,
    input wire [3:0]                      AP_AXIMM_75_ARQOS,
    input wire                            AP_AXIMM_75_ARVALID,
    output  wire                            AP_AXIMM_75_ARREADY,
    output  wire [M_AXIMM_75_DATA_WIDTH-1:0]   AP_AXIMM_75_RDATA,
    output  wire [1:0]                      AP_AXIMM_75_RRESP,
    output  wire                            AP_AXIMM_75_RLAST,
    output  wire                            AP_AXIMM_75_RVALID,
    input  wire                            AP_AXIMM_75_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_75_AWADDR,
    output wire [7:0]                      M_AXIMM_75_AWLEN,
    output wire [2:0]                      M_AXIMM_75_AWSIZE,
    output wire [1:0]                      M_AXIMM_75_AWBURST,
    output wire [1:0]                      M_AXIMM_75_AWLOCK,
    output wire [3:0]                      M_AXIMM_75_AWCACHE,
    output wire [2:0]                      M_AXIMM_75_AWPROT,
    output wire [3:0]                      M_AXIMM_75_AWREGION,
    output wire [3:0]                      M_AXIMM_75_AWQOS,
    output wire                            M_AXIMM_75_AWVALID,
    input  wire                            M_AXIMM_75_AWREADY,
    output wire [M_AXIMM_75_DATA_WIDTH-1:0]   M_AXIMM_75_WDATA,
    output wire [M_AXIMM_75_DATA_WIDTH/8-1:0] M_AXIMM_75_WSTRB,
    output wire                            M_AXIMM_75_WLAST,
    output wire                            M_AXIMM_75_WVALID,
    input  wire                            M_AXIMM_75_WREADY,
    input  wire [1:0]                      M_AXIMM_75_BRESP,
    input  wire                            M_AXIMM_75_BVALID,
    output wire                            M_AXIMM_75_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_75_ARADDR,
    output wire [7:0]                      M_AXIMM_75_ARLEN,
    output wire [2:0]                      M_AXIMM_75_ARSIZE,
    output wire [1:0]                      M_AXIMM_75_ARBURST,
    output wire [1:0]                      M_AXIMM_75_ARLOCK,
    output wire [3:0]                      M_AXIMM_75_ARCACHE,
    output wire [2:0]                      M_AXIMM_75_ARPROT,
    output wire [3:0]                      M_AXIMM_75_ARREGION,
    output wire [3:0]                      M_AXIMM_75_ARQOS,
    output wire                            M_AXIMM_75_ARVALID,
    input  wire                            M_AXIMM_75_ARREADY,
    input  wire [M_AXIMM_75_DATA_WIDTH-1:0]   M_AXIMM_75_RDATA,
    input  wire [1:0]                      M_AXIMM_75_RRESP,
    input  wire                            M_AXIMM_75_RLAST,
    input  wire                            M_AXIMM_75_RVALID,
    output wire                            M_AXIMM_75_RREADY,
    //AXI-MM pass-through interface 76
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_76_AWADDR,
    input wire [7:0]                      AP_AXIMM_76_AWLEN,
    input wire [2:0]                      AP_AXIMM_76_AWSIZE,
    input wire [1:0]                      AP_AXIMM_76_AWBURST,
    input wire [1:0]                      AP_AXIMM_76_AWLOCK,
    input wire [3:0]                      AP_AXIMM_76_AWCACHE,
    input wire [2:0]                      AP_AXIMM_76_AWPROT,
    input wire [3:0]                      AP_AXIMM_76_AWREGION,
    input wire [3:0]                      AP_AXIMM_76_AWQOS,
    input wire                            AP_AXIMM_76_AWVALID,
    output  wire                            AP_AXIMM_76_AWREADY,
    input wire [M_AXIMM_76_DATA_WIDTH-1:0]   AP_AXIMM_76_WDATA,
    input wire [M_AXIMM_76_DATA_WIDTH/8-1:0] AP_AXIMM_76_WSTRB,
    input wire                            AP_AXIMM_76_WLAST,
    input wire                            AP_AXIMM_76_WVALID,
    output  wire                            AP_AXIMM_76_WREADY,
    output  wire [1:0]                      AP_AXIMM_76_BRESP,
    output  wire                            AP_AXIMM_76_BVALID,
    input wire                            AP_AXIMM_76_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_76_ARADDR,
    input wire [7:0]                      AP_AXIMM_76_ARLEN,
    input wire [2:0]                      AP_AXIMM_76_ARSIZE,
    input wire [1:0]                      AP_AXIMM_76_ARBURST,
    input wire [1:0]                      AP_AXIMM_76_ARLOCK,
    input wire [3:0]                      AP_AXIMM_76_ARCACHE,
    input wire [2:0]                      AP_AXIMM_76_ARPROT,
    input wire [3:0]                      AP_AXIMM_76_ARREGION,
    input wire [3:0]                      AP_AXIMM_76_ARQOS,
    input wire                            AP_AXIMM_76_ARVALID,
    output  wire                            AP_AXIMM_76_ARREADY,
    output  wire [M_AXIMM_76_DATA_WIDTH-1:0]   AP_AXIMM_76_RDATA,
    output  wire [1:0]                      AP_AXIMM_76_RRESP,
    output  wire                            AP_AXIMM_76_RLAST,
    output  wire                            AP_AXIMM_76_RVALID,
    input  wire                            AP_AXIMM_76_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_76_AWADDR,
    output wire [7:0]                      M_AXIMM_76_AWLEN,
    output wire [2:0]                      M_AXIMM_76_AWSIZE,
    output wire [1:0]                      M_AXIMM_76_AWBURST,
    output wire [1:0]                      M_AXIMM_76_AWLOCK,
    output wire [3:0]                      M_AXIMM_76_AWCACHE,
    output wire [2:0]                      M_AXIMM_76_AWPROT,
    output wire [3:0]                      M_AXIMM_76_AWREGION,
    output wire [3:0]                      M_AXIMM_76_AWQOS,
    output wire                            M_AXIMM_76_AWVALID,
    input  wire                            M_AXIMM_76_AWREADY,
    output wire [M_AXIMM_76_DATA_WIDTH-1:0]   M_AXIMM_76_WDATA,
    output wire [M_AXIMM_76_DATA_WIDTH/8-1:0] M_AXIMM_76_WSTRB,
    output wire                            M_AXIMM_76_WLAST,
    output wire                            M_AXIMM_76_WVALID,
    input  wire                            M_AXIMM_76_WREADY,
    input  wire [1:0]                      M_AXIMM_76_BRESP,
    input  wire                            M_AXIMM_76_BVALID,
    output wire                            M_AXIMM_76_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_76_ARADDR,
    output wire [7:0]                      M_AXIMM_76_ARLEN,
    output wire [2:0]                      M_AXIMM_76_ARSIZE,
    output wire [1:0]                      M_AXIMM_76_ARBURST,
    output wire [1:0]                      M_AXIMM_76_ARLOCK,
    output wire [3:0]                      M_AXIMM_76_ARCACHE,
    output wire [2:0]                      M_AXIMM_76_ARPROT,
    output wire [3:0]                      M_AXIMM_76_ARREGION,
    output wire [3:0]                      M_AXIMM_76_ARQOS,
    output wire                            M_AXIMM_76_ARVALID,
    input  wire                            M_AXIMM_76_ARREADY,
    input  wire [M_AXIMM_76_DATA_WIDTH-1:0]   M_AXIMM_76_RDATA,
    input  wire [1:0]                      M_AXIMM_76_RRESP,
    input  wire                            M_AXIMM_76_RLAST,
    input  wire                            M_AXIMM_76_RVALID,
    output wire                            M_AXIMM_76_RREADY,
    //AXI-MM pass-through interface 77
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_77_AWADDR,
    input wire [7:0]                      AP_AXIMM_77_AWLEN,
    input wire [2:0]                      AP_AXIMM_77_AWSIZE,
    input wire [1:0]                      AP_AXIMM_77_AWBURST,
    input wire [1:0]                      AP_AXIMM_77_AWLOCK,
    input wire [3:0]                      AP_AXIMM_77_AWCACHE,
    input wire [2:0]                      AP_AXIMM_77_AWPROT,
    input wire [3:0]                      AP_AXIMM_77_AWREGION,
    input wire [3:0]                      AP_AXIMM_77_AWQOS,
    input wire                            AP_AXIMM_77_AWVALID,
    output  wire                            AP_AXIMM_77_AWREADY,
    input wire [M_AXIMM_77_DATA_WIDTH-1:0]   AP_AXIMM_77_WDATA,
    input wire [M_AXIMM_77_DATA_WIDTH/8-1:0] AP_AXIMM_77_WSTRB,
    input wire                            AP_AXIMM_77_WLAST,
    input wire                            AP_AXIMM_77_WVALID,
    output  wire                            AP_AXIMM_77_WREADY,
    output  wire [1:0]                      AP_AXIMM_77_BRESP,
    output  wire                            AP_AXIMM_77_BVALID,
    input wire                            AP_AXIMM_77_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_77_ARADDR,
    input wire [7:0]                      AP_AXIMM_77_ARLEN,
    input wire [2:0]                      AP_AXIMM_77_ARSIZE,
    input wire [1:0]                      AP_AXIMM_77_ARBURST,
    input wire [1:0]                      AP_AXIMM_77_ARLOCK,
    input wire [3:0]                      AP_AXIMM_77_ARCACHE,
    input wire [2:0]                      AP_AXIMM_77_ARPROT,
    input wire [3:0]                      AP_AXIMM_77_ARREGION,
    input wire [3:0]                      AP_AXIMM_77_ARQOS,
    input wire                            AP_AXIMM_77_ARVALID,
    output  wire                            AP_AXIMM_77_ARREADY,
    output  wire [M_AXIMM_77_DATA_WIDTH-1:0]   AP_AXIMM_77_RDATA,
    output  wire [1:0]                      AP_AXIMM_77_RRESP,
    output  wire                            AP_AXIMM_77_RLAST,
    output  wire                            AP_AXIMM_77_RVALID,
    input  wire                            AP_AXIMM_77_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_77_AWADDR,
    output wire [7:0]                      M_AXIMM_77_AWLEN,
    output wire [2:0]                      M_AXIMM_77_AWSIZE,
    output wire [1:0]                      M_AXIMM_77_AWBURST,
    output wire [1:0]                      M_AXIMM_77_AWLOCK,
    output wire [3:0]                      M_AXIMM_77_AWCACHE,
    output wire [2:0]                      M_AXIMM_77_AWPROT,
    output wire [3:0]                      M_AXIMM_77_AWREGION,
    output wire [3:0]                      M_AXIMM_77_AWQOS,
    output wire                            M_AXIMM_77_AWVALID,
    input  wire                            M_AXIMM_77_AWREADY,
    output wire [M_AXIMM_77_DATA_WIDTH-1:0]   M_AXIMM_77_WDATA,
    output wire [M_AXIMM_77_DATA_WIDTH/8-1:0] M_AXIMM_77_WSTRB,
    output wire                            M_AXIMM_77_WLAST,
    output wire                            M_AXIMM_77_WVALID,
    input  wire                            M_AXIMM_77_WREADY,
    input  wire [1:0]                      M_AXIMM_77_BRESP,
    input  wire                            M_AXIMM_77_BVALID,
    output wire                            M_AXIMM_77_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_77_ARADDR,
    output wire [7:0]                      M_AXIMM_77_ARLEN,
    output wire [2:0]                      M_AXIMM_77_ARSIZE,
    output wire [1:0]                      M_AXIMM_77_ARBURST,
    output wire [1:0]                      M_AXIMM_77_ARLOCK,
    output wire [3:0]                      M_AXIMM_77_ARCACHE,
    output wire [2:0]                      M_AXIMM_77_ARPROT,
    output wire [3:0]                      M_AXIMM_77_ARREGION,
    output wire [3:0]                      M_AXIMM_77_ARQOS,
    output wire                            M_AXIMM_77_ARVALID,
    input  wire                            M_AXIMM_77_ARREADY,
    input  wire [M_AXIMM_77_DATA_WIDTH-1:0]   M_AXIMM_77_RDATA,
    input  wire [1:0]                      M_AXIMM_77_RRESP,
    input  wire                            M_AXIMM_77_RLAST,
    input  wire                            M_AXIMM_77_RVALID,
    output wire                            M_AXIMM_77_RREADY,
    //AXI-MM pass-through interface 78
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_78_AWADDR,
    input wire [7:0]                      AP_AXIMM_78_AWLEN,
    input wire [2:0]                      AP_AXIMM_78_AWSIZE,
    input wire [1:0]                      AP_AXIMM_78_AWBURST,
    input wire [1:0]                      AP_AXIMM_78_AWLOCK,
    input wire [3:0]                      AP_AXIMM_78_AWCACHE,
    input wire [2:0]                      AP_AXIMM_78_AWPROT,
    input wire [3:0]                      AP_AXIMM_78_AWREGION,
    input wire [3:0]                      AP_AXIMM_78_AWQOS,
    input wire                            AP_AXIMM_78_AWVALID,
    output  wire                            AP_AXIMM_78_AWREADY,
    input wire [M_AXIMM_78_DATA_WIDTH-1:0]   AP_AXIMM_78_WDATA,
    input wire [M_AXIMM_78_DATA_WIDTH/8-1:0] AP_AXIMM_78_WSTRB,
    input wire                            AP_AXIMM_78_WLAST,
    input wire                            AP_AXIMM_78_WVALID,
    output  wire                            AP_AXIMM_78_WREADY,
    output  wire [1:0]                      AP_AXIMM_78_BRESP,
    output  wire                            AP_AXIMM_78_BVALID,
    input wire                            AP_AXIMM_78_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_78_ARADDR,
    input wire [7:0]                      AP_AXIMM_78_ARLEN,
    input wire [2:0]                      AP_AXIMM_78_ARSIZE,
    input wire [1:0]                      AP_AXIMM_78_ARBURST,
    input wire [1:0]                      AP_AXIMM_78_ARLOCK,
    input wire [3:0]                      AP_AXIMM_78_ARCACHE,
    input wire [2:0]                      AP_AXIMM_78_ARPROT,
    input wire [3:0]                      AP_AXIMM_78_ARREGION,
    input wire [3:0]                      AP_AXIMM_78_ARQOS,
    input wire                            AP_AXIMM_78_ARVALID,
    output  wire                            AP_AXIMM_78_ARREADY,
    output  wire [M_AXIMM_78_DATA_WIDTH-1:0]   AP_AXIMM_78_RDATA,
    output  wire [1:0]                      AP_AXIMM_78_RRESP,
    output  wire                            AP_AXIMM_78_RLAST,
    output  wire                            AP_AXIMM_78_RVALID,
    input  wire                            AP_AXIMM_78_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_78_AWADDR,
    output wire [7:0]                      M_AXIMM_78_AWLEN,
    output wire [2:0]                      M_AXIMM_78_AWSIZE,
    output wire [1:0]                      M_AXIMM_78_AWBURST,
    output wire [1:0]                      M_AXIMM_78_AWLOCK,
    output wire [3:0]                      M_AXIMM_78_AWCACHE,
    output wire [2:0]                      M_AXIMM_78_AWPROT,
    output wire [3:0]                      M_AXIMM_78_AWREGION,
    output wire [3:0]                      M_AXIMM_78_AWQOS,
    output wire                            M_AXIMM_78_AWVALID,
    input  wire                            M_AXIMM_78_AWREADY,
    output wire [M_AXIMM_78_DATA_WIDTH-1:0]   M_AXIMM_78_WDATA,
    output wire [M_AXIMM_78_DATA_WIDTH/8-1:0] M_AXIMM_78_WSTRB,
    output wire                            M_AXIMM_78_WLAST,
    output wire                            M_AXIMM_78_WVALID,
    input  wire                            M_AXIMM_78_WREADY,
    input  wire [1:0]                      M_AXIMM_78_BRESP,
    input  wire                            M_AXIMM_78_BVALID,
    output wire                            M_AXIMM_78_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_78_ARADDR,
    output wire [7:0]                      M_AXIMM_78_ARLEN,
    output wire [2:0]                      M_AXIMM_78_ARSIZE,
    output wire [1:0]                      M_AXIMM_78_ARBURST,
    output wire [1:0]                      M_AXIMM_78_ARLOCK,
    output wire [3:0]                      M_AXIMM_78_ARCACHE,
    output wire [2:0]                      M_AXIMM_78_ARPROT,
    output wire [3:0]                      M_AXIMM_78_ARREGION,
    output wire [3:0]                      M_AXIMM_78_ARQOS,
    output wire                            M_AXIMM_78_ARVALID,
    input  wire                            M_AXIMM_78_ARREADY,
    input  wire [M_AXIMM_78_DATA_WIDTH-1:0]   M_AXIMM_78_RDATA,
    input  wire [1:0]                      M_AXIMM_78_RRESP,
    input  wire                            M_AXIMM_78_RLAST,
    input  wire                            M_AXIMM_78_RVALID,
    output wire                            M_AXIMM_78_RREADY,
    //AXI-MM pass-through interface 79
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_79_AWADDR,
    input wire [7:0]                      AP_AXIMM_79_AWLEN,
    input wire [2:0]                      AP_AXIMM_79_AWSIZE,
    input wire [1:0]                      AP_AXIMM_79_AWBURST,
    input wire [1:0]                      AP_AXIMM_79_AWLOCK,
    input wire [3:0]                      AP_AXIMM_79_AWCACHE,
    input wire [2:0]                      AP_AXIMM_79_AWPROT,
    input wire [3:0]                      AP_AXIMM_79_AWREGION,
    input wire [3:0]                      AP_AXIMM_79_AWQOS,
    input wire                            AP_AXIMM_79_AWVALID,
    output  wire                            AP_AXIMM_79_AWREADY,
    input wire [M_AXIMM_79_DATA_WIDTH-1:0]   AP_AXIMM_79_WDATA,
    input wire [M_AXIMM_79_DATA_WIDTH/8-1:0] AP_AXIMM_79_WSTRB,
    input wire                            AP_AXIMM_79_WLAST,
    input wire                            AP_AXIMM_79_WVALID,
    output  wire                            AP_AXIMM_79_WREADY,
    output  wire [1:0]                      AP_AXIMM_79_BRESP,
    output  wire                            AP_AXIMM_79_BVALID,
    input wire                            AP_AXIMM_79_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_79_ARADDR,
    input wire [7:0]                      AP_AXIMM_79_ARLEN,
    input wire [2:0]                      AP_AXIMM_79_ARSIZE,
    input wire [1:0]                      AP_AXIMM_79_ARBURST,
    input wire [1:0]                      AP_AXIMM_79_ARLOCK,
    input wire [3:0]                      AP_AXIMM_79_ARCACHE,
    input wire [2:0]                      AP_AXIMM_79_ARPROT,
    input wire [3:0]                      AP_AXIMM_79_ARREGION,
    input wire [3:0]                      AP_AXIMM_79_ARQOS,
    input wire                            AP_AXIMM_79_ARVALID,
    output  wire                            AP_AXIMM_79_ARREADY,
    output  wire [M_AXIMM_79_DATA_WIDTH-1:0]   AP_AXIMM_79_RDATA,
    output  wire [1:0]                      AP_AXIMM_79_RRESP,
    output  wire                            AP_AXIMM_79_RLAST,
    output  wire                            AP_AXIMM_79_RVALID,
    input  wire                            AP_AXIMM_79_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_79_AWADDR,
    output wire [7:0]                      M_AXIMM_79_AWLEN,
    output wire [2:0]                      M_AXIMM_79_AWSIZE,
    output wire [1:0]                      M_AXIMM_79_AWBURST,
    output wire [1:0]                      M_AXIMM_79_AWLOCK,
    output wire [3:0]                      M_AXIMM_79_AWCACHE,
    output wire [2:0]                      M_AXIMM_79_AWPROT,
    output wire [3:0]                      M_AXIMM_79_AWREGION,
    output wire [3:0]                      M_AXIMM_79_AWQOS,
    output wire                            M_AXIMM_79_AWVALID,
    input  wire                            M_AXIMM_79_AWREADY,
    output wire [M_AXIMM_79_DATA_WIDTH-1:0]   M_AXIMM_79_WDATA,
    output wire [M_AXIMM_79_DATA_WIDTH/8-1:0] M_AXIMM_79_WSTRB,
    output wire                            M_AXIMM_79_WLAST,
    output wire                            M_AXIMM_79_WVALID,
    input  wire                            M_AXIMM_79_WREADY,
    input  wire [1:0]                      M_AXIMM_79_BRESP,
    input  wire                            M_AXIMM_79_BVALID,
    output wire                            M_AXIMM_79_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_79_ARADDR,
    output wire [7:0]                      M_AXIMM_79_ARLEN,
    output wire [2:0]                      M_AXIMM_79_ARSIZE,
    output wire [1:0]                      M_AXIMM_79_ARBURST,
    output wire [1:0]                      M_AXIMM_79_ARLOCK,
    output wire [3:0]                      M_AXIMM_79_ARCACHE,
    output wire [2:0]                      M_AXIMM_79_ARPROT,
    output wire [3:0]                      M_AXIMM_79_ARREGION,
    output wire [3:0]                      M_AXIMM_79_ARQOS,
    output wire                            M_AXIMM_79_ARVALID,
    input  wire                            M_AXIMM_79_ARREADY,
    input  wire [M_AXIMM_79_DATA_WIDTH-1:0]   M_AXIMM_79_RDATA,
    input  wire [1:0]                      M_AXIMM_79_RRESP,
    input  wire                            M_AXIMM_79_RLAST,
    input  wire                            M_AXIMM_79_RVALID,
    output wire                            M_AXIMM_79_RREADY,
    //AXI-MM pass-through interface 80
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_80_AWADDR,
    input wire [7:0]                      AP_AXIMM_80_AWLEN,
    input wire [2:0]                      AP_AXIMM_80_AWSIZE,
    input wire [1:0]                      AP_AXIMM_80_AWBURST,
    input wire [1:0]                      AP_AXIMM_80_AWLOCK,
    input wire [3:0]                      AP_AXIMM_80_AWCACHE,
    input wire [2:0]                      AP_AXIMM_80_AWPROT,
    input wire [3:0]                      AP_AXIMM_80_AWREGION,
    input wire [3:0]                      AP_AXIMM_80_AWQOS,
    input wire                            AP_AXIMM_80_AWVALID,
    output  wire                            AP_AXIMM_80_AWREADY,
    input wire [M_AXIMM_80_DATA_WIDTH-1:0]   AP_AXIMM_80_WDATA,
    input wire [M_AXIMM_80_DATA_WIDTH/8-1:0] AP_AXIMM_80_WSTRB,
    input wire                            AP_AXIMM_80_WLAST,
    input wire                            AP_AXIMM_80_WVALID,
    output  wire                            AP_AXIMM_80_WREADY,
    output  wire [1:0]                      AP_AXIMM_80_BRESP,
    output  wire                            AP_AXIMM_80_BVALID,
    input wire                            AP_AXIMM_80_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_80_ARADDR,
    input wire [7:0]                      AP_AXIMM_80_ARLEN,
    input wire [2:0]                      AP_AXIMM_80_ARSIZE,
    input wire [1:0]                      AP_AXIMM_80_ARBURST,
    input wire [1:0]                      AP_AXIMM_80_ARLOCK,
    input wire [3:0]                      AP_AXIMM_80_ARCACHE,
    input wire [2:0]                      AP_AXIMM_80_ARPROT,
    input wire [3:0]                      AP_AXIMM_80_ARREGION,
    input wire [3:0]                      AP_AXIMM_80_ARQOS,
    input wire                            AP_AXIMM_80_ARVALID,
    output  wire                            AP_AXIMM_80_ARREADY,
    output  wire [M_AXIMM_80_DATA_WIDTH-1:0]   AP_AXIMM_80_RDATA,
    output  wire [1:0]                      AP_AXIMM_80_RRESP,
    output  wire                            AP_AXIMM_80_RLAST,
    output  wire                            AP_AXIMM_80_RVALID,
    input  wire                            AP_AXIMM_80_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_80_AWADDR,
    output wire [7:0]                      M_AXIMM_80_AWLEN,
    output wire [2:0]                      M_AXIMM_80_AWSIZE,
    output wire [1:0]                      M_AXIMM_80_AWBURST,
    output wire [1:0]                      M_AXIMM_80_AWLOCK,
    output wire [3:0]                      M_AXIMM_80_AWCACHE,
    output wire [2:0]                      M_AXIMM_80_AWPROT,
    output wire [3:0]                      M_AXIMM_80_AWREGION,
    output wire [3:0]                      M_AXIMM_80_AWQOS,
    output wire                            M_AXIMM_80_AWVALID,
    input  wire                            M_AXIMM_80_AWREADY,
    output wire [M_AXIMM_80_DATA_WIDTH-1:0]   M_AXIMM_80_WDATA,
    output wire [M_AXIMM_80_DATA_WIDTH/8-1:0] M_AXIMM_80_WSTRB,
    output wire                            M_AXIMM_80_WLAST,
    output wire                            M_AXIMM_80_WVALID,
    input  wire                            M_AXIMM_80_WREADY,
    input  wire [1:0]                      M_AXIMM_80_BRESP,
    input  wire                            M_AXIMM_80_BVALID,
    output wire                            M_AXIMM_80_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_80_ARADDR,
    output wire [7:0]                      M_AXIMM_80_ARLEN,
    output wire [2:0]                      M_AXIMM_80_ARSIZE,
    output wire [1:0]                      M_AXIMM_80_ARBURST,
    output wire [1:0]                      M_AXIMM_80_ARLOCK,
    output wire [3:0]                      M_AXIMM_80_ARCACHE,
    output wire [2:0]                      M_AXIMM_80_ARPROT,
    output wire [3:0]                      M_AXIMM_80_ARREGION,
    output wire [3:0]                      M_AXIMM_80_ARQOS,
    output wire                            M_AXIMM_80_ARVALID,
    input  wire                            M_AXIMM_80_ARREADY,
    input  wire [M_AXIMM_80_DATA_WIDTH-1:0]   M_AXIMM_80_RDATA,
    input  wire [1:0]                      M_AXIMM_80_RRESP,
    input  wire                            M_AXIMM_80_RLAST,
    input  wire                            M_AXIMM_80_RVALID,
    output wire                            M_AXIMM_80_RREADY,
    //AXI-MM pass-through interface 81
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_81_AWADDR,
    input wire [7:0]                      AP_AXIMM_81_AWLEN,
    input wire [2:0]                      AP_AXIMM_81_AWSIZE,
    input wire [1:0]                      AP_AXIMM_81_AWBURST,
    input wire [1:0]                      AP_AXIMM_81_AWLOCK,
    input wire [3:0]                      AP_AXIMM_81_AWCACHE,
    input wire [2:0]                      AP_AXIMM_81_AWPROT,
    input wire [3:0]                      AP_AXIMM_81_AWREGION,
    input wire [3:0]                      AP_AXIMM_81_AWQOS,
    input wire                            AP_AXIMM_81_AWVALID,
    output  wire                            AP_AXIMM_81_AWREADY,
    input wire [M_AXIMM_81_DATA_WIDTH-1:0]   AP_AXIMM_81_WDATA,
    input wire [M_AXIMM_81_DATA_WIDTH/8-1:0] AP_AXIMM_81_WSTRB,
    input wire                            AP_AXIMM_81_WLAST,
    input wire                            AP_AXIMM_81_WVALID,
    output  wire                            AP_AXIMM_81_WREADY,
    output  wire [1:0]                      AP_AXIMM_81_BRESP,
    output  wire                            AP_AXIMM_81_BVALID,
    input wire                            AP_AXIMM_81_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_81_ARADDR,
    input wire [7:0]                      AP_AXIMM_81_ARLEN,
    input wire [2:0]                      AP_AXIMM_81_ARSIZE,
    input wire [1:0]                      AP_AXIMM_81_ARBURST,
    input wire [1:0]                      AP_AXIMM_81_ARLOCK,
    input wire [3:0]                      AP_AXIMM_81_ARCACHE,
    input wire [2:0]                      AP_AXIMM_81_ARPROT,
    input wire [3:0]                      AP_AXIMM_81_ARREGION,
    input wire [3:0]                      AP_AXIMM_81_ARQOS,
    input wire                            AP_AXIMM_81_ARVALID,
    output  wire                            AP_AXIMM_81_ARREADY,
    output  wire [M_AXIMM_81_DATA_WIDTH-1:0]   AP_AXIMM_81_RDATA,
    output  wire [1:0]                      AP_AXIMM_81_RRESP,
    output  wire                            AP_AXIMM_81_RLAST,
    output  wire                            AP_AXIMM_81_RVALID,
    input  wire                            AP_AXIMM_81_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_81_AWADDR,
    output wire [7:0]                      M_AXIMM_81_AWLEN,
    output wire [2:0]                      M_AXIMM_81_AWSIZE,
    output wire [1:0]                      M_AXIMM_81_AWBURST,
    output wire [1:0]                      M_AXIMM_81_AWLOCK,
    output wire [3:0]                      M_AXIMM_81_AWCACHE,
    output wire [2:0]                      M_AXIMM_81_AWPROT,
    output wire [3:0]                      M_AXIMM_81_AWREGION,
    output wire [3:0]                      M_AXIMM_81_AWQOS,
    output wire                            M_AXIMM_81_AWVALID,
    input  wire                            M_AXIMM_81_AWREADY,
    output wire [M_AXIMM_81_DATA_WIDTH-1:0]   M_AXIMM_81_WDATA,
    output wire [M_AXIMM_81_DATA_WIDTH/8-1:0] M_AXIMM_81_WSTRB,
    output wire                            M_AXIMM_81_WLAST,
    output wire                            M_AXIMM_81_WVALID,
    input  wire                            M_AXIMM_81_WREADY,
    input  wire [1:0]                      M_AXIMM_81_BRESP,
    input  wire                            M_AXIMM_81_BVALID,
    output wire                            M_AXIMM_81_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_81_ARADDR,
    output wire [7:0]                      M_AXIMM_81_ARLEN,
    output wire [2:0]                      M_AXIMM_81_ARSIZE,
    output wire [1:0]                      M_AXIMM_81_ARBURST,
    output wire [1:0]                      M_AXIMM_81_ARLOCK,
    output wire [3:0]                      M_AXIMM_81_ARCACHE,
    output wire [2:0]                      M_AXIMM_81_ARPROT,
    output wire [3:0]                      M_AXIMM_81_ARREGION,
    output wire [3:0]                      M_AXIMM_81_ARQOS,
    output wire                            M_AXIMM_81_ARVALID,
    input  wire                            M_AXIMM_81_ARREADY,
    input  wire [M_AXIMM_81_DATA_WIDTH-1:0]   M_AXIMM_81_RDATA,
    input  wire [1:0]                      M_AXIMM_81_RRESP,
    input  wire                            M_AXIMM_81_RLAST,
    input  wire                            M_AXIMM_81_RVALID,
    output wire                            M_AXIMM_81_RREADY,
    //AXI-MM pass-through interface 82
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_82_AWADDR,
    input wire [7:0]                      AP_AXIMM_82_AWLEN,
    input wire [2:0]                      AP_AXIMM_82_AWSIZE,
    input wire [1:0]                      AP_AXIMM_82_AWBURST,
    input wire [1:0]                      AP_AXIMM_82_AWLOCK,
    input wire [3:0]                      AP_AXIMM_82_AWCACHE,
    input wire [2:0]                      AP_AXIMM_82_AWPROT,
    input wire [3:0]                      AP_AXIMM_82_AWREGION,
    input wire [3:0]                      AP_AXIMM_82_AWQOS,
    input wire                            AP_AXIMM_82_AWVALID,
    output  wire                            AP_AXIMM_82_AWREADY,
    input wire [M_AXIMM_82_DATA_WIDTH-1:0]   AP_AXIMM_82_WDATA,
    input wire [M_AXIMM_82_DATA_WIDTH/8-1:0] AP_AXIMM_82_WSTRB,
    input wire                            AP_AXIMM_82_WLAST,
    input wire                            AP_AXIMM_82_WVALID,
    output  wire                            AP_AXIMM_82_WREADY,
    output  wire [1:0]                      AP_AXIMM_82_BRESP,
    output  wire                            AP_AXIMM_82_BVALID,
    input wire                            AP_AXIMM_82_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_82_ARADDR,
    input wire [7:0]                      AP_AXIMM_82_ARLEN,
    input wire [2:0]                      AP_AXIMM_82_ARSIZE,
    input wire [1:0]                      AP_AXIMM_82_ARBURST,
    input wire [1:0]                      AP_AXIMM_82_ARLOCK,
    input wire [3:0]                      AP_AXIMM_82_ARCACHE,
    input wire [2:0]                      AP_AXIMM_82_ARPROT,
    input wire [3:0]                      AP_AXIMM_82_ARREGION,
    input wire [3:0]                      AP_AXIMM_82_ARQOS,
    input wire                            AP_AXIMM_82_ARVALID,
    output  wire                            AP_AXIMM_82_ARREADY,
    output  wire [M_AXIMM_82_DATA_WIDTH-1:0]   AP_AXIMM_82_RDATA,
    output  wire [1:0]                      AP_AXIMM_82_RRESP,
    output  wire                            AP_AXIMM_82_RLAST,
    output  wire                            AP_AXIMM_82_RVALID,
    input  wire                            AP_AXIMM_82_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_82_AWADDR,
    output wire [7:0]                      M_AXIMM_82_AWLEN,
    output wire [2:0]                      M_AXIMM_82_AWSIZE,
    output wire [1:0]                      M_AXIMM_82_AWBURST,
    output wire [1:0]                      M_AXIMM_82_AWLOCK,
    output wire [3:0]                      M_AXIMM_82_AWCACHE,
    output wire [2:0]                      M_AXIMM_82_AWPROT,
    output wire [3:0]                      M_AXIMM_82_AWREGION,
    output wire [3:0]                      M_AXIMM_82_AWQOS,
    output wire                            M_AXIMM_82_AWVALID,
    input  wire                            M_AXIMM_82_AWREADY,
    output wire [M_AXIMM_82_DATA_WIDTH-1:0]   M_AXIMM_82_WDATA,
    output wire [M_AXIMM_82_DATA_WIDTH/8-1:0] M_AXIMM_82_WSTRB,
    output wire                            M_AXIMM_82_WLAST,
    output wire                            M_AXIMM_82_WVALID,
    input  wire                            M_AXIMM_82_WREADY,
    input  wire [1:0]                      M_AXIMM_82_BRESP,
    input  wire                            M_AXIMM_82_BVALID,
    output wire                            M_AXIMM_82_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_82_ARADDR,
    output wire [7:0]                      M_AXIMM_82_ARLEN,
    output wire [2:0]                      M_AXIMM_82_ARSIZE,
    output wire [1:0]                      M_AXIMM_82_ARBURST,
    output wire [1:0]                      M_AXIMM_82_ARLOCK,
    output wire [3:0]                      M_AXIMM_82_ARCACHE,
    output wire [2:0]                      M_AXIMM_82_ARPROT,
    output wire [3:0]                      M_AXIMM_82_ARREGION,
    output wire [3:0]                      M_AXIMM_82_ARQOS,
    output wire                            M_AXIMM_82_ARVALID,
    input  wire                            M_AXIMM_82_ARREADY,
    input  wire [M_AXIMM_82_DATA_WIDTH-1:0]   M_AXIMM_82_RDATA,
    input  wire [1:0]                      M_AXIMM_82_RRESP,
    input  wire                            M_AXIMM_82_RLAST,
    input  wire                            M_AXIMM_82_RVALID,
    output wire                            M_AXIMM_82_RREADY,
    //AXI-MM pass-through interface 83
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_83_AWADDR,
    input wire [7:0]                      AP_AXIMM_83_AWLEN,
    input wire [2:0]                      AP_AXIMM_83_AWSIZE,
    input wire [1:0]                      AP_AXIMM_83_AWBURST,
    input wire [1:0]                      AP_AXIMM_83_AWLOCK,
    input wire [3:0]                      AP_AXIMM_83_AWCACHE,
    input wire [2:0]                      AP_AXIMM_83_AWPROT,
    input wire [3:0]                      AP_AXIMM_83_AWREGION,
    input wire [3:0]                      AP_AXIMM_83_AWQOS,
    input wire                            AP_AXIMM_83_AWVALID,
    output  wire                            AP_AXIMM_83_AWREADY,
    input wire [M_AXIMM_83_DATA_WIDTH-1:0]   AP_AXIMM_83_WDATA,
    input wire [M_AXIMM_83_DATA_WIDTH/8-1:0] AP_AXIMM_83_WSTRB,
    input wire                            AP_AXIMM_83_WLAST,
    input wire                            AP_AXIMM_83_WVALID,
    output  wire                            AP_AXIMM_83_WREADY,
    output  wire [1:0]                      AP_AXIMM_83_BRESP,
    output  wire                            AP_AXIMM_83_BVALID,
    input wire                            AP_AXIMM_83_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_83_ARADDR,
    input wire [7:0]                      AP_AXIMM_83_ARLEN,
    input wire [2:0]                      AP_AXIMM_83_ARSIZE,
    input wire [1:0]                      AP_AXIMM_83_ARBURST,
    input wire [1:0]                      AP_AXIMM_83_ARLOCK,
    input wire [3:0]                      AP_AXIMM_83_ARCACHE,
    input wire [2:0]                      AP_AXIMM_83_ARPROT,
    input wire [3:0]                      AP_AXIMM_83_ARREGION,
    input wire [3:0]                      AP_AXIMM_83_ARQOS,
    input wire                            AP_AXIMM_83_ARVALID,
    output  wire                            AP_AXIMM_83_ARREADY,
    output  wire [M_AXIMM_83_DATA_WIDTH-1:0]   AP_AXIMM_83_RDATA,
    output  wire [1:0]                      AP_AXIMM_83_RRESP,
    output  wire                            AP_AXIMM_83_RLAST,
    output  wire                            AP_AXIMM_83_RVALID,
    input  wire                            AP_AXIMM_83_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_83_AWADDR,
    output wire [7:0]                      M_AXIMM_83_AWLEN,
    output wire [2:0]                      M_AXIMM_83_AWSIZE,
    output wire [1:0]                      M_AXIMM_83_AWBURST,
    output wire [1:0]                      M_AXIMM_83_AWLOCK,
    output wire [3:0]                      M_AXIMM_83_AWCACHE,
    output wire [2:0]                      M_AXIMM_83_AWPROT,
    output wire [3:0]                      M_AXIMM_83_AWREGION,
    output wire [3:0]                      M_AXIMM_83_AWQOS,
    output wire                            M_AXIMM_83_AWVALID,
    input  wire                            M_AXIMM_83_AWREADY,
    output wire [M_AXIMM_83_DATA_WIDTH-1:0]   M_AXIMM_83_WDATA,
    output wire [M_AXIMM_83_DATA_WIDTH/8-1:0] M_AXIMM_83_WSTRB,
    output wire                            M_AXIMM_83_WLAST,
    output wire                            M_AXIMM_83_WVALID,
    input  wire                            M_AXIMM_83_WREADY,
    input  wire [1:0]                      M_AXIMM_83_BRESP,
    input  wire                            M_AXIMM_83_BVALID,
    output wire                            M_AXIMM_83_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_83_ARADDR,
    output wire [7:0]                      M_AXIMM_83_ARLEN,
    output wire [2:0]                      M_AXIMM_83_ARSIZE,
    output wire [1:0]                      M_AXIMM_83_ARBURST,
    output wire [1:0]                      M_AXIMM_83_ARLOCK,
    output wire [3:0]                      M_AXIMM_83_ARCACHE,
    output wire [2:0]                      M_AXIMM_83_ARPROT,
    output wire [3:0]                      M_AXIMM_83_ARREGION,
    output wire [3:0]                      M_AXIMM_83_ARQOS,
    output wire                            M_AXIMM_83_ARVALID,
    input  wire                            M_AXIMM_83_ARREADY,
    input  wire [M_AXIMM_83_DATA_WIDTH-1:0]   M_AXIMM_83_RDATA,
    input  wire [1:0]                      M_AXIMM_83_RRESP,
    input  wire                            M_AXIMM_83_RLAST,
    input  wire                            M_AXIMM_83_RVALID,
    output wire                            M_AXIMM_83_RREADY,
    //AXI-MM pass-through interface 84
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_84_AWADDR,
    input wire [7:0]                      AP_AXIMM_84_AWLEN,
    input wire [2:0]                      AP_AXIMM_84_AWSIZE,
    input wire [1:0]                      AP_AXIMM_84_AWBURST,
    input wire [1:0]                      AP_AXIMM_84_AWLOCK,
    input wire [3:0]                      AP_AXIMM_84_AWCACHE,
    input wire [2:0]                      AP_AXIMM_84_AWPROT,
    input wire [3:0]                      AP_AXIMM_84_AWREGION,
    input wire [3:0]                      AP_AXIMM_84_AWQOS,
    input wire                            AP_AXIMM_84_AWVALID,
    output  wire                            AP_AXIMM_84_AWREADY,
    input wire [M_AXIMM_84_DATA_WIDTH-1:0]   AP_AXIMM_84_WDATA,
    input wire [M_AXIMM_84_DATA_WIDTH/8-1:0] AP_AXIMM_84_WSTRB,
    input wire                            AP_AXIMM_84_WLAST,
    input wire                            AP_AXIMM_84_WVALID,
    output  wire                            AP_AXIMM_84_WREADY,
    output  wire [1:0]                      AP_AXIMM_84_BRESP,
    output  wire                            AP_AXIMM_84_BVALID,
    input wire                            AP_AXIMM_84_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_84_ARADDR,
    input wire [7:0]                      AP_AXIMM_84_ARLEN,
    input wire [2:0]                      AP_AXIMM_84_ARSIZE,
    input wire [1:0]                      AP_AXIMM_84_ARBURST,
    input wire [1:0]                      AP_AXIMM_84_ARLOCK,
    input wire [3:0]                      AP_AXIMM_84_ARCACHE,
    input wire [2:0]                      AP_AXIMM_84_ARPROT,
    input wire [3:0]                      AP_AXIMM_84_ARREGION,
    input wire [3:0]                      AP_AXIMM_84_ARQOS,
    input wire                            AP_AXIMM_84_ARVALID,
    output  wire                            AP_AXIMM_84_ARREADY,
    output  wire [M_AXIMM_84_DATA_WIDTH-1:0]   AP_AXIMM_84_RDATA,
    output  wire [1:0]                      AP_AXIMM_84_RRESP,
    output  wire                            AP_AXIMM_84_RLAST,
    output  wire                            AP_AXIMM_84_RVALID,
    input  wire                            AP_AXIMM_84_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_84_AWADDR,
    output wire [7:0]                      M_AXIMM_84_AWLEN,
    output wire [2:0]                      M_AXIMM_84_AWSIZE,
    output wire [1:0]                      M_AXIMM_84_AWBURST,
    output wire [1:0]                      M_AXIMM_84_AWLOCK,
    output wire [3:0]                      M_AXIMM_84_AWCACHE,
    output wire [2:0]                      M_AXIMM_84_AWPROT,
    output wire [3:0]                      M_AXIMM_84_AWREGION,
    output wire [3:0]                      M_AXIMM_84_AWQOS,
    output wire                            M_AXIMM_84_AWVALID,
    input  wire                            M_AXIMM_84_AWREADY,
    output wire [M_AXIMM_84_DATA_WIDTH-1:0]   M_AXIMM_84_WDATA,
    output wire [M_AXIMM_84_DATA_WIDTH/8-1:0] M_AXIMM_84_WSTRB,
    output wire                            M_AXIMM_84_WLAST,
    output wire                            M_AXIMM_84_WVALID,
    input  wire                            M_AXIMM_84_WREADY,
    input  wire [1:0]                      M_AXIMM_84_BRESP,
    input  wire                            M_AXIMM_84_BVALID,
    output wire                            M_AXIMM_84_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_84_ARADDR,
    output wire [7:0]                      M_AXIMM_84_ARLEN,
    output wire [2:0]                      M_AXIMM_84_ARSIZE,
    output wire [1:0]                      M_AXIMM_84_ARBURST,
    output wire [1:0]                      M_AXIMM_84_ARLOCK,
    output wire [3:0]                      M_AXIMM_84_ARCACHE,
    output wire [2:0]                      M_AXIMM_84_ARPROT,
    output wire [3:0]                      M_AXIMM_84_ARREGION,
    output wire [3:0]                      M_AXIMM_84_ARQOS,
    output wire                            M_AXIMM_84_ARVALID,
    input  wire                            M_AXIMM_84_ARREADY,
    input  wire [M_AXIMM_84_DATA_WIDTH-1:0]   M_AXIMM_84_RDATA,
    input  wire [1:0]                      M_AXIMM_84_RRESP,
    input  wire                            M_AXIMM_84_RLAST,
    input  wire                            M_AXIMM_84_RVALID,
    output wire                            M_AXIMM_84_RREADY,
    //AXI-MM pass-through interface 85
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_85_AWADDR,
    input wire [7:0]                      AP_AXIMM_85_AWLEN,
    input wire [2:0]                      AP_AXIMM_85_AWSIZE,
    input wire [1:0]                      AP_AXIMM_85_AWBURST,
    input wire [1:0]                      AP_AXIMM_85_AWLOCK,
    input wire [3:0]                      AP_AXIMM_85_AWCACHE,
    input wire [2:0]                      AP_AXIMM_85_AWPROT,
    input wire [3:0]                      AP_AXIMM_85_AWREGION,
    input wire [3:0]                      AP_AXIMM_85_AWQOS,
    input wire                            AP_AXIMM_85_AWVALID,
    output  wire                            AP_AXIMM_85_AWREADY,
    input wire [M_AXIMM_85_DATA_WIDTH-1:0]   AP_AXIMM_85_WDATA,
    input wire [M_AXIMM_85_DATA_WIDTH/8-1:0] AP_AXIMM_85_WSTRB,
    input wire                            AP_AXIMM_85_WLAST,
    input wire                            AP_AXIMM_85_WVALID,
    output  wire                            AP_AXIMM_85_WREADY,
    output  wire [1:0]                      AP_AXIMM_85_BRESP,
    output  wire                            AP_AXIMM_85_BVALID,
    input wire                            AP_AXIMM_85_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_85_ARADDR,
    input wire [7:0]                      AP_AXIMM_85_ARLEN,
    input wire [2:0]                      AP_AXIMM_85_ARSIZE,
    input wire [1:0]                      AP_AXIMM_85_ARBURST,
    input wire [1:0]                      AP_AXIMM_85_ARLOCK,
    input wire [3:0]                      AP_AXIMM_85_ARCACHE,
    input wire [2:0]                      AP_AXIMM_85_ARPROT,
    input wire [3:0]                      AP_AXIMM_85_ARREGION,
    input wire [3:0]                      AP_AXIMM_85_ARQOS,
    input wire                            AP_AXIMM_85_ARVALID,
    output  wire                            AP_AXIMM_85_ARREADY,
    output  wire [M_AXIMM_85_DATA_WIDTH-1:0]   AP_AXIMM_85_RDATA,
    output  wire [1:0]                      AP_AXIMM_85_RRESP,
    output  wire                            AP_AXIMM_85_RLAST,
    output  wire                            AP_AXIMM_85_RVALID,
    input  wire                            AP_AXIMM_85_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_85_AWADDR,
    output wire [7:0]                      M_AXIMM_85_AWLEN,
    output wire [2:0]                      M_AXIMM_85_AWSIZE,
    output wire [1:0]                      M_AXIMM_85_AWBURST,
    output wire [1:0]                      M_AXIMM_85_AWLOCK,
    output wire [3:0]                      M_AXIMM_85_AWCACHE,
    output wire [2:0]                      M_AXIMM_85_AWPROT,
    output wire [3:0]                      M_AXIMM_85_AWREGION,
    output wire [3:0]                      M_AXIMM_85_AWQOS,
    output wire                            M_AXIMM_85_AWVALID,
    input  wire                            M_AXIMM_85_AWREADY,
    output wire [M_AXIMM_85_DATA_WIDTH-1:0]   M_AXIMM_85_WDATA,
    output wire [M_AXIMM_85_DATA_WIDTH/8-1:0] M_AXIMM_85_WSTRB,
    output wire                            M_AXIMM_85_WLAST,
    output wire                            M_AXIMM_85_WVALID,
    input  wire                            M_AXIMM_85_WREADY,
    input  wire [1:0]                      M_AXIMM_85_BRESP,
    input  wire                            M_AXIMM_85_BVALID,
    output wire                            M_AXIMM_85_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_85_ARADDR,
    output wire [7:0]                      M_AXIMM_85_ARLEN,
    output wire [2:0]                      M_AXIMM_85_ARSIZE,
    output wire [1:0]                      M_AXIMM_85_ARBURST,
    output wire [1:0]                      M_AXIMM_85_ARLOCK,
    output wire [3:0]                      M_AXIMM_85_ARCACHE,
    output wire [2:0]                      M_AXIMM_85_ARPROT,
    output wire [3:0]                      M_AXIMM_85_ARREGION,
    output wire [3:0]                      M_AXIMM_85_ARQOS,
    output wire                            M_AXIMM_85_ARVALID,
    input  wire                            M_AXIMM_85_ARREADY,
    input  wire [M_AXIMM_85_DATA_WIDTH-1:0]   M_AXIMM_85_RDATA,
    input  wire [1:0]                      M_AXIMM_85_RRESP,
    input  wire                            M_AXIMM_85_RLAST,
    input  wire                            M_AXIMM_85_RVALID,
    output wire                            M_AXIMM_85_RREADY,
    //AXI-MM pass-through interface 86
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_86_AWADDR,
    input wire [7:0]                      AP_AXIMM_86_AWLEN,
    input wire [2:0]                      AP_AXIMM_86_AWSIZE,
    input wire [1:0]                      AP_AXIMM_86_AWBURST,
    input wire [1:0]                      AP_AXIMM_86_AWLOCK,
    input wire [3:0]                      AP_AXIMM_86_AWCACHE,
    input wire [2:0]                      AP_AXIMM_86_AWPROT,
    input wire [3:0]                      AP_AXIMM_86_AWREGION,
    input wire [3:0]                      AP_AXIMM_86_AWQOS,
    input wire                            AP_AXIMM_86_AWVALID,
    output  wire                            AP_AXIMM_86_AWREADY,
    input wire [M_AXIMM_86_DATA_WIDTH-1:0]   AP_AXIMM_86_WDATA,
    input wire [M_AXIMM_86_DATA_WIDTH/8-1:0] AP_AXIMM_86_WSTRB,
    input wire                            AP_AXIMM_86_WLAST,
    input wire                            AP_AXIMM_86_WVALID,
    output  wire                            AP_AXIMM_86_WREADY,
    output  wire [1:0]                      AP_AXIMM_86_BRESP,
    output  wire                            AP_AXIMM_86_BVALID,
    input wire                            AP_AXIMM_86_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_86_ARADDR,
    input wire [7:0]                      AP_AXIMM_86_ARLEN,
    input wire [2:0]                      AP_AXIMM_86_ARSIZE,
    input wire [1:0]                      AP_AXIMM_86_ARBURST,
    input wire [1:0]                      AP_AXIMM_86_ARLOCK,
    input wire [3:0]                      AP_AXIMM_86_ARCACHE,
    input wire [2:0]                      AP_AXIMM_86_ARPROT,
    input wire [3:0]                      AP_AXIMM_86_ARREGION,
    input wire [3:0]                      AP_AXIMM_86_ARQOS,
    input wire                            AP_AXIMM_86_ARVALID,
    output  wire                            AP_AXIMM_86_ARREADY,
    output  wire [M_AXIMM_86_DATA_WIDTH-1:0]   AP_AXIMM_86_RDATA,
    output  wire [1:0]                      AP_AXIMM_86_RRESP,
    output  wire                            AP_AXIMM_86_RLAST,
    output  wire                            AP_AXIMM_86_RVALID,
    input  wire                            AP_AXIMM_86_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_86_AWADDR,
    output wire [7:0]                      M_AXIMM_86_AWLEN,
    output wire [2:0]                      M_AXIMM_86_AWSIZE,
    output wire [1:0]                      M_AXIMM_86_AWBURST,
    output wire [1:0]                      M_AXIMM_86_AWLOCK,
    output wire [3:0]                      M_AXIMM_86_AWCACHE,
    output wire [2:0]                      M_AXIMM_86_AWPROT,
    output wire [3:0]                      M_AXIMM_86_AWREGION,
    output wire [3:0]                      M_AXIMM_86_AWQOS,
    output wire                            M_AXIMM_86_AWVALID,
    input  wire                            M_AXIMM_86_AWREADY,
    output wire [M_AXIMM_86_DATA_WIDTH-1:0]   M_AXIMM_86_WDATA,
    output wire [M_AXIMM_86_DATA_WIDTH/8-1:0] M_AXIMM_86_WSTRB,
    output wire                            M_AXIMM_86_WLAST,
    output wire                            M_AXIMM_86_WVALID,
    input  wire                            M_AXIMM_86_WREADY,
    input  wire [1:0]                      M_AXIMM_86_BRESP,
    input  wire                            M_AXIMM_86_BVALID,
    output wire                            M_AXIMM_86_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_86_ARADDR,
    output wire [7:0]                      M_AXIMM_86_ARLEN,
    output wire [2:0]                      M_AXIMM_86_ARSIZE,
    output wire [1:0]                      M_AXIMM_86_ARBURST,
    output wire [1:0]                      M_AXIMM_86_ARLOCK,
    output wire [3:0]                      M_AXIMM_86_ARCACHE,
    output wire [2:0]                      M_AXIMM_86_ARPROT,
    output wire [3:0]                      M_AXIMM_86_ARREGION,
    output wire [3:0]                      M_AXIMM_86_ARQOS,
    output wire                            M_AXIMM_86_ARVALID,
    input  wire                            M_AXIMM_86_ARREADY,
    input  wire [M_AXIMM_86_DATA_WIDTH-1:0]   M_AXIMM_86_RDATA,
    input  wire [1:0]                      M_AXIMM_86_RRESP,
    input  wire                            M_AXIMM_86_RLAST,
    input  wire                            M_AXIMM_86_RVALID,
    output wire                            M_AXIMM_86_RREADY,
    //AXI-MM pass-through interface 87
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_87_AWADDR,
    input wire [7:0]                      AP_AXIMM_87_AWLEN,
    input wire [2:0]                      AP_AXIMM_87_AWSIZE,
    input wire [1:0]                      AP_AXIMM_87_AWBURST,
    input wire [1:0]                      AP_AXIMM_87_AWLOCK,
    input wire [3:0]                      AP_AXIMM_87_AWCACHE,
    input wire [2:0]                      AP_AXIMM_87_AWPROT,
    input wire [3:0]                      AP_AXIMM_87_AWREGION,
    input wire [3:0]                      AP_AXIMM_87_AWQOS,
    input wire                            AP_AXIMM_87_AWVALID,
    output  wire                            AP_AXIMM_87_AWREADY,
    input wire [M_AXIMM_87_DATA_WIDTH-1:0]   AP_AXIMM_87_WDATA,
    input wire [M_AXIMM_87_DATA_WIDTH/8-1:0] AP_AXIMM_87_WSTRB,
    input wire                            AP_AXIMM_87_WLAST,
    input wire                            AP_AXIMM_87_WVALID,
    output  wire                            AP_AXIMM_87_WREADY,
    output  wire [1:0]                      AP_AXIMM_87_BRESP,
    output  wire                            AP_AXIMM_87_BVALID,
    input wire                            AP_AXIMM_87_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_87_ARADDR,
    input wire [7:0]                      AP_AXIMM_87_ARLEN,
    input wire [2:0]                      AP_AXIMM_87_ARSIZE,
    input wire [1:0]                      AP_AXIMM_87_ARBURST,
    input wire [1:0]                      AP_AXIMM_87_ARLOCK,
    input wire [3:0]                      AP_AXIMM_87_ARCACHE,
    input wire [2:0]                      AP_AXIMM_87_ARPROT,
    input wire [3:0]                      AP_AXIMM_87_ARREGION,
    input wire [3:0]                      AP_AXIMM_87_ARQOS,
    input wire                            AP_AXIMM_87_ARVALID,
    output  wire                            AP_AXIMM_87_ARREADY,
    output  wire [M_AXIMM_87_DATA_WIDTH-1:0]   AP_AXIMM_87_RDATA,
    output  wire [1:0]                      AP_AXIMM_87_RRESP,
    output  wire                            AP_AXIMM_87_RLAST,
    output  wire                            AP_AXIMM_87_RVALID,
    input  wire                            AP_AXIMM_87_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_87_AWADDR,
    output wire [7:0]                      M_AXIMM_87_AWLEN,
    output wire [2:0]                      M_AXIMM_87_AWSIZE,
    output wire [1:0]                      M_AXIMM_87_AWBURST,
    output wire [1:0]                      M_AXIMM_87_AWLOCK,
    output wire [3:0]                      M_AXIMM_87_AWCACHE,
    output wire [2:0]                      M_AXIMM_87_AWPROT,
    output wire [3:0]                      M_AXIMM_87_AWREGION,
    output wire [3:0]                      M_AXIMM_87_AWQOS,
    output wire                            M_AXIMM_87_AWVALID,
    input  wire                            M_AXIMM_87_AWREADY,
    output wire [M_AXIMM_87_DATA_WIDTH-1:0]   M_AXIMM_87_WDATA,
    output wire [M_AXIMM_87_DATA_WIDTH/8-1:0] M_AXIMM_87_WSTRB,
    output wire                            M_AXIMM_87_WLAST,
    output wire                            M_AXIMM_87_WVALID,
    input  wire                            M_AXIMM_87_WREADY,
    input  wire [1:0]                      M_AXIMM_87_BRESP,
    input  wire                            M_AXIMM_87_BVALID,
    output wire                            M_AXIMM_87_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_87_ARADDR,
    output wire [7:0]                      M_AXIMM_87_ARLEN,
    output wire [2:0]                      M_AXIMM_87_ARSIZE,
    output wire [1:0]                      M_AXIMM_87_ARBURST,
    output wire [1:0]                      M_AXIMM_87_ARLOCK,
    output wire [3:0]                      M_AXIMM_87_ARCACHE,
    output wire [2:0]                      M_AXIMM_87_ARPROT,
    output wire [3:0]                      M_AXIMM_87_ARREGION,
    output wire [3:0]                      M_AXIMM_87_ARQOS,
    output wire                            M_AXIMM_87_ARVALID,
    input  wire                            M_AXIMM_87_ARREADY,
    input  wire [M_AXIMM_87_DATA_WIDTH-1:0]   M_AXIMM_87_RDATA,
    input  wire [1:0]                      M_AXIMM_87_RRESP,
    input  wire                            M_AXIMM_87_RLAST,
    input  wire                            M_AXIMM_87_RVALID,
    output wire                            M_AXIMM_87_RREADY,
    //AXI-MM pass-through interface 88
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_88_AWADDR,
    input wire [7:0]                      AP_AXIMM_88_AWLEN,
    input wire [2:0]                      AP_AXIMM_88_AWSIZE,
    input wire [1:0]                      AP_AXIMM_88_AWBURST,
    input wire [1:0]                      AP_AXIMM_88_AWLOCK,
    input wire [3:0]                      AP_AXIMM_88_AWCACHE,
    input wire [2:0]                      AP_AXIMM_88_AWPROT,
    input wire [3:0]                      AP_AXIMM_88_AWREGION,
    input wire [3:0]                      AP_AXIMM_88_AWQOS,
    input wire                            AP_AXIMM_88_AWVALID,
    output  wire                            AP_AXIMM_88_AWREADY,
    input wire [M_AXIMM_88_DATA_WIDTH-1:0]   AP_AXIMM_88_WDATA,
    input wire [M_AXIMM_88_DATA_WIDTH/8-1:0] AP_AXIMM_88_WSTRB,
    input wire                            AP_AXIMM_88_WLAST,
    input wire                            AP_AXIMM_88_WVALID,
    output  wire                            AP_AXIMM_88_WREADY,
    output  wire [1:0]                      AP_AXIMM_88_BRESP,
    output  wire                            AP_AXIMM_88_BVALID,
    input wire                            AP_AXIMM_88_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_88_ARADDR,
    input wire [7:0]                      AP_AXIMM_88_ARLEN,
    input wire [2:0]                      AP_AXIMM_88_ARSIZE,
    input wire [1:0]                      AP_AXIMM_88_ARBURST,
    input wire [1:0]                      AP_AXIMM_88_ARLOCK,
    input wire [3:0]                      AP_AXIMM_88_ARCACHE,
    input wire [2:0]                      AP_AXIMM_88_ARPROT,
    input wire [3:0]                      AP_AXIMM_88_ARREGION,
    input wire [3:0]                      AP_AXIMM_88_ARQOS,
    input wire                            AP_AXIMM_88_ARVALID,
    output  wire                            AP_AXIMM_88_ARREADY,
    output  wire [M_AXIMM_88_DATA_WIDTH-1:0]   AP_AXIMM_88_RDATA,
    output  wire [1:0]                      AP_AXIMM_88_RRESP,
    output  wire                            AP_AXIMM_88_RLAST,
    output  wire                            AP_AXIMM_88_RVALID,
    input  wire                            AP_AXIMM_88_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_88_AWADDR,
    output wire [7:0]                      M_AXIMM_88_AWLEN,
    output wire [2:0]                      M_AXIMM_88_AWSIZE,
    output wire [1:0]                      M_AXIMM_88_AWBURST,
    output wire [1:0]                      M_AXIMM_88_AWLOCK,
    output wire [3:0]                      M_AXIMM_88_AWCACHE,
    output wire [2:0]                      M_AXIMM_88_AWPROT,
    output wire [3:0]                      M_AXIMM_88_AWREGION,
    output wire [3:0]                      M_AXIMM_88_AWQOS,
    output wire                            M_AXIMM_88_AWVALID,
    input  wire                            M_AXIMM_88_AWREADY,
    output wire [M_AXIMM_88_DATA_WIDTH-1:0]   M_AXIMM_88_WDATA,
    output wire [M_AXIMM_88_DATA_WIDTH/8-1:0] M_AXIMM_88_WSTRB,
    output wire                            M_AXIMM_88_WLAST,
    output wire                            M_AXIMM_88_WVALID,
    input  wire                            M_AXIMM_88_WREADY,
    input  wire [1:0]                      M_AXIMM_88_BRESP,
    input  wire                            M_AXIMM_88_BVALID,
    output wire                            M_AXIMM_88_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_88_ARADDR,
    output wire [7:0]                      M_AXIMM_88_ARLEN,
    output wire [2:0]                      M_AXIMM_88_ARSIZE,
    output wire [1:0]                      M_AXIMM_88_ARBURST,
    output wire [1:0]                      M_AXIMM_88_ARLOCK,
    output wire [3:0]                      M_AXIMM_88_ARCACHE,
    output wire [2:0]                      M_AXIMM_88_ARPROT,
    output wire [3:0]                      M_AXIMM_88_ARREGION,
    output wire [3:0]                      M_AXIMM_88_ARQOS,
    output wire                            M_AXIMM_88_ARVALID,
    input  wire                            M_AXIMM_88_ARREADY,
    input  wire [M_AXIMM_88_DATA_WIDTH-1:0]   M_AXIMM_88_RDATA,
    input  wire [1:0]                      M_AXIMM_88_RRESP,
    input  wire                            M_AXIMM_88_RLAST,
    input  wire                            M_AXIMM_88_RVALID,
    output wire                            M_AXIMM_88_RREADY,
    //AXI-MM pass-through interface 89
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_89_AWADDR,
    input wire [7:0]                      AP_AXIMM_89_AWLEN,
    input wire [2:0]                      AP_AXIMM_89_AWSIZE,
    input wire [1:0]                      AP_AXIMM_89_AWBURST,
    input wire [1:0]                      AP_AXIMM_89_AWLOCK,
    input wire [3:0]                      AP_AXIMM_89_AWCACHE,
    input wire [2:0]                      AP_AXIMM_89_AWPROT,
    input wire [3:0]                      AP_AXIMM_89_AWREGION,
    input wire [3:0]                      AP_AXIMM_89_AWQOS,
    input wire                            AP_AXIMM_89_AWVALID,
    output  wire                            AP_AXIMM_89_AWREADY,
    input wire [M_AXIMM_89_DATA_WIDTH-1:0]   AP_AXIMM_89_WDATA,
    input wire [M_AXIMM_89_DATA_WIDTH/8-1:0] AP_AXIMM_89_WSTRB,
    input wire                            AP_AXIMM_89_WLAST,
    input wire                            AP_AXIMM_89_WVALID,
    output  wire                            AP_AXIMM_89_WREADY,
    output  wire [1:0]                      AP_AXIMM_89_BRESP,
    output  wire                            AP_AXIMM_89_BVALID,
    input wire                            AP_AXIMM_89_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_89_ARADDR,
    input wire [7:0]                      AP_AXIMM_89_ARLEN,
    input wire [2:0]                      AP_AXIMM_89_ARSIZE,
    input wire [1:0]                      AP_AXIMM_89_ARBURST,
    input wire [1:0]                      AP_AXIMM_89_ARLOCK,
    input wire [3:0]                      AP_AXIMM_89_ARCACHE,
    input wire [2:0]                      AP_AXIMM_89_ARPROT,
    input wire [3:0]                      AP_AXIMM_89_ARREGION,
    input wire [3:0]                      AP_AXIMM_89_ARQOS,
    input wire                            AP_AXIMM_89_ARVALID,
    output  wire                            AP_AXIMM_89_ARREADY,
    output  wire [M_AXIMM_89_DATA_WIDTH-1:0]   AP_AXIMM_89_RDATA,
    output  wire [1:0]                      AP_AXIMM_89_RRESP,
    output  wire                            AP_AXIMM_89_RLAST,
    output  wire                            AP_AXIMM_89_RVALID,
    input  wire                            AP_AXIMM_89_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_89_AWADDR,
    output wire [7:0]                      M_AXIMM_89_AWLEN,
    output wire [2:0]                      M_AXIMM_89_AWSIZE,
    output wire [1:0]                      M_AXIMM_89_AWBURST,
    output wire [1:0]                      M_AXIMM_89_AWLOCK,
    output wire [3:0]                      M_AXIMM_89_AWCACHE,
    output wire [2:0]                      M_AXIMM_89_AWPROT,
    output wire [3:0]                      M_AXIMM_89_AWREGION,
    output wire [3:0]                      M_AXIMM_89_AWQOS,
    output wire                            M_AXIMM_89_AWVALID,
    input  wire                            M_AXIMM_89_AWREADY,
    output wire [M_AXIMM_89_DATA_WIDTH-1:0]   M_AXIMM_89_WDATA,
    output wire [M_AXIMM_89_DATA_WIDTH/8-1:0] M_AXIMM_89_WSTRB,
    output wire                            M_AXIMM_89_WLAST,
    output wire                            M_AXIMM_89_WVALID,
    input  wire                            M_AXIMM_89_WREADY,
    input  wire [1:0]                      M_AXIMM_89_BRESP,
    input  wire                            M_AXIMM_89_BVALID,
    output wire                            M_AXIMM_89_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_89_ARADDR,
    output wire [7:0]                      M_AXIMM_89_ARLEN,
    output wire [2:0]                      M_AXIMM_89_ARSIZE,
    output wire [1:0]                      M_AXIMM_89_ARBURST,
    output wire [1:0]                      M_AXIMM_89_ARLOCK,
    output wire [3:0]                      M_AXIMM_89_ARCACHE,
    output wire [2:0]                      M_AXIMM_89_ARPROT,
    output wire [3:0]                      M_AXIMM_89_ARREGION,
    output wire [3:0]                      M_AXIMM_89_ARQOS,
    output wire                            M_AXIMM_89_ARVALID,
    input  wire                            M_AXIMM_89_ARREADY,
    input  wire [M_AXIMM_89_DATA_WIDTH-1:0]   M_AXIMM_89_RDATA,
    input  wire [1:0]                      M_AXIMM_89_RRESP,
    input  wire                            M_AXIMM_89_RLAST,
    input  wire                            M_AXIMM_89_RVALID,
    output wire                            M_AXIMM_89_RREADY,
    //AXI-MM pass-through interface 90
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_90_AWADDR,
    input wire [7:0]                      AP_AXIMM_90_AWLEN,
    input wire [2:0]                      AP_AXIMM_90_AWSIZE,
    input wire [1:0]                      AP_AXIMM_90_AWBURST,
    input wire [1:0]                      AP_AXIMM_90_AWLOCK,
    input wire [3:0]                      AP_AXIMM_90_AWCACHE,
    input wire [2:0]                      AP_AXIMM_90_AWPROT,
    input wire [3:0]                      AP_AXIMM_90_AWREGION,
    input wire [3:0]                      AP_AXIMM_90_AWQOS,
    input wire                            AP_AXIMM_90_AWVALID,
    output  wire                            AP_AXIMM_90_AWREADY,
    input wire [M_AXIMM_90_DATA_WIDTH-1:0]   AP_AXIMM_90_WDATA,
    input wire [M_AXIMM_90_DATA_WIDTH/8-1:0] AP_AXIMM_90_WSTRB,
    input wire                            AP_AXIMM_90_WLAST,
    input wire                            AP_AXIMM_90_WVALID,
    output  wire                            AP_AXIMM_90_WREADY,
    output  wire [1:0]                      AP_AXIMM_90_BRESP,
    output  wire                            AP_AXIMM_90_BVALID,
    input wire                            AP_AXIMM_90_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_90_ARADDR,
    input wire [7:0]                      AP_AXIMM_90_ARLEN,
    input wire [2:0]                      AP_AXIMM_90_ARSIZE,
    input wire [1:0]                      AP_AXIMM_90_ARBURST,
    input wire [1:0]                      AP_AXIMM_90_ARLOCK,
    input wire [3:0]                      AP_AXIMM_90_ARCACHE,
    input wire [2:0]                      AP_AXIMM_90_ARPROT,
    input wire [3:0]                      AP_AXIMM_90_ARREGION,
    input wire [3:0]                      AP_AXIMM_90_ARQOS,
    input wire                            AP_AXIMM_90_ARVALID,
    output  wire                            AP_AXIMM_90_ARREADY,
    output  wire [M_AXIMM_90_DATA_WIDTH-1:0]   AP_AXIMM_90_RDATA,
    output  wire [1:0]                      AP_AXIMM_90_RRESP,
    output  wire                            AP_AXIMM_90_RLAST,
    output  wire                            AP_AXIMM_90_RVALID,
    input  wire                            AP_AXIMM_90_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_90_AWADDR,
    output wire [7:0]                      M_AXIMM_90_AWLEN,
    output wire [2:0]                      M_AXIMM_90_AWSIZE,
    output wire [1:0]                      M_AXIMM_90_AWBURST,
    output wire [1:0]                      M_AXIMM_90_AWLOCK,
    output wire [3:0]                      M_AXIMM_90_AWCACHE,
    output wire [2:0]                      M_AXIMM_90_AWPROT,
    output wire [3:0]                      M_AXIMM_90_AWREGION,
    output wire [3:0]                      M_AXIMM_90_AWQOS,
    output wire                            M_AXIMM_90_AWVALID,
    input  wire                            M_AXIMM_90_AWREADY,
    output wire [M_AXIMM_90_DATA_WIDTH-1:0]   M_AXIMM_90_WDATA,
    output wire [M_AXIMM_90_DATA_WIDTH/8-1:0] M_AXIMM_90_WSTRB,
    output wire                            M_AXIMM_90_WLAST,
    output wire                            M_AXIMM_90_WVALID,
    input  wire                            M_AXIMM_90_WREADY,
    input  wire [1:0]                      M_AXIMM_90_BRESP,
    input  wire                            M_AXIMM_90_BVALID,
    output wire                            M_AXIMM_90_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_90_ARADDR,
    output wire [7:0]                      M_AXIMM_90_ARLEN,
    output wire [2:0]                      M_AXIMM_90_ARSIZE,
    output wire [1:0]                      M_AXIMM_90_ARBURST,
    output wire [1:0]                      M_AXIMM_90_ARLOCK,
    output wire [3:0]                      M_AXIMM_90_ARCACHE,
    output wire [2:0]                      M_AXIMM_90_ARPROT,
    output wire [3:0]                      M_AXIMM_90_ARREGION,
    output wire [3:0]                      M_AXIMM_90_ARQOS,
    output wire                            M_AXIMM_90_ARVALID,
    input  wire                            M_AXIMM_90_ARREADY,
    input  wire [M_AXIMM_90_DATA_WIDTH-1:0]   M_AXIMM_90_RDATA,
    input  wire [1:0]                      M_AXIMM_90_RRESP,
    input  wire                            M_AXIMM_90_RLAST,
    input  wire                            M_AXIMM_90_RVALID,
    output wire                            M_AXIMM_90_RREADY,
    //AXI-MM pass-through interface 91
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_91_AWADDR,
    input wire [7:0]                      AP_AXIMM_91_AWLEN,
    input wire [2:0]                      AP_AXIMM_91_AWSIZE,
    input wire [1:0]                      AP_AXIMM_91_AWBURST,
    input wire [1:0]                      AP_AXIMM_91_AWLOCK,
    input wire [3:0]                      AP_AXIMM_91_AWCACHE,
    input wire [2:0]                      AP_AXIMM_91_AWPROT,
    input wire [3:0]                      AP_AXIMM_91_AWREGION,
    input wire [3:0]                      AP_AXIMM_91_AWQOS,
    input wire                            AP_AXIMM_91_AWVALID,
    output  wire                            AP_AXIMM_91_AWREADY,
    input wire [M_AXIMM_91_DATA_WIDTH-1:0]   AP_AXIMM_91_WDATA,
    input wire [M_AXIMM_91_DATA_WIDTH/8-1:0] AP_AXIMM_91_WSTRB,
    input wire                            AP_AXIMM_91_WLAST,
    input wire                            AP_AXIMM_91_WVALID,
    output  wire                            AP_AXIMM_91_WREADY,
    output  wire [1:0]                      AP_AXIMM_91_BRESP,
    output  wire                            AP_AXIMM_91_BVALID,
    input wire                            AP_AXIMM_91_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_91_ARADDR,
    input wire [7:0]                      AP_AXIMM_91_ARLEN,
    input wire [2:0]                      AP_AXIMM_91_ARSIZE,
    input wire [1:0]                      AP_AXIMM_91_ARBURST,
    input wire [1:0]                      AP_AXIMM_91_ARLOCK,
    input wire [3:0]                      AP_AXIMM_91_ARCACHE,
    input wire [2:0]                      AP_AXIMM_91_ARPROT,
    input wire [3:0]                      AP_AXIMM_91_ARREGION,
    input wire [3:0]                      AP_AXIMM_91_ARQOS,
    input wire                            AP_AXIMM_91_ARVALID,
    output  wire                            AP_AXIMM_91_ARREADY,
    output  wire [M_AXIMM_91_DATA_WIDTH-1:0]   AP_AXIMM_91_RDATA,
    output  wire [1:0]                      AP_AXIMM_91_RRESP,
    output  wire                            AP_AXIMM_91_RLAST,
    output  wire                            AP_AXIMM_91_RVALID,
    input  wire                            AP_AXIMM_91_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_91_AWADDR,
    output wire [7:0]                      M_AXIMM_91_AWLEN,
    output wire [2:0]                      M_AXIMM_91_AWSIZE,
    output wire [1:0]                      M_AXIMM_91_AWBURST,
    output wire [1:0]                      M_AXIMM_91_AWLOCK,
    output wire [3:0]                      M_AXIMM_91_AWCACHE,
    output wire [2:0]                      M_AXIMM_91_AWPROT,
    output wire [3:0]                      M_AXIMM_91_AWREGION,
    output wire [3:0]                      M_AXIMM_91_AWQOS,
    output wire                            M_AXIMM_91_AWVALID,
    input  wire                            M_AXIMM_91_AWREADY,
    output wire [M_AXIMM_91_DATA_WIDTH-1:0]   M_AXIMM_91_WDATA,
    output wire [M_AXIMM_91_DATA_WIDTH/8-1:0] M_AXIMM_91_WSTRB,
    output wire                            M_AXIMM_91_WLAST,
    output wire                            M_AXIMM_91_WVALID,
    input  wire                            M_AXIMM_91_WREADY,
    input  wire [1:0]                      M_AXIMM_91_BRESP,
    input  wire                            M_AXIMM_91_BVALID,
    output wire                            M_AXIMM_91_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_91_ARADDR,
    output wire [7:0]                      M_AXIMM_91_ARLEN,
    output wire [2:0]                      M_AXIMM_91_ARSIZE,
    output wire [1:0]                      M_AXIMM_91_ARBURST,
    output wire [1:0]                      M_AXIMM_91_ARLOCK,
    output wire [3:0]                      M_AXIMM_91_ARCACHE,
    output wire [2:0]                      M_AXIMM_91_ARPROT,
    output wire [3:0]                      M_AXIMM_91_ARREGION,
    output wire [3:0]                      M_AXIMM_91_ARQOS,
    output wire                            M_AXIMM_91_ARVALID,
    input  wire                            M_AXIMM_91_ARREADY,
    input  wire [M_AXIMM_91_DATA_WIDTH-1:0]   M_AXIMM_91_RDATA,
    input  wire [1:0]                      M_AXIMM_91_RRESP,
    input  wire                            M_AXIMM_91_RLAST,
    input  wire                            M_AXIMM_91_RVALID,
    output wire                            M_AXIMM_91_RREADY,
    //AXI-MM pass-through interface 92
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_92_AWADDR,
    input wire [7:0]                      AP_AXIMM_92_AWLEN,
    input wire [2:0]                      AP_AXIMM_92_AWSIZE,
    input wire [1:0]                      AP_AXIMM_92_AWBURST,
    input wire [1:0]                      AP_AXIMM_92_AWLOCK,
    input wire [3:0]                      AP_AXIMM_92_AWCACHE,
    input wire [2:0]                      AP_AXIMM_92_AWPROT,
    input wire [3:0]                      AP_AXIMM_92_AWREGION,
    input wire [3:0]                      AP_AXIMM_92_AWQOS,
    input wire                            AP_AXIMM_92_AWVALID,
    output  wire                            AP_AXIMM_92_AWREADY,
    input wire [M_AXIMM_92_DATA_WIDTH-1:0]   AP_AXIMM_92_WDATA,
    input wire [M_AXIMM_92_DATA_WIDTH/8-1:0] AP_AXIMM_92_WSTRB,
    input wire                            AP_AXIMM_92_WLAST,
    input wire                            AP_AXIMM_92_WVALID,
    output  wire                            AP_AXIMM_92_WREADY,
    output  wire [1:0]                      AP_AXIMM_92_BRESP,
    output  wire                            AP_AXIMM_92_BVALID,
    input wire                            AP_AXIMM_92_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_92_ARADDR,
    input wire [7:0]                      AP_AXIMM_92_ARLEN,
    input wire [2:0]                      AP_AXIMM_92_ARSIZE,
    input wire [1:0]                      AP_AXIMM_92_ARBURST,
    input wire [1:0]                      AP_AXIMM_92_ARLOCK,
    input wire [3:0]                      AP_AXIMM_92_ARCACHE,
    input wire [2:0]                      AP_AXIMM_92_ARPROT,
    input wire [3:0]                      AP_AXIMM_92_ARREGION,
    input wire [3:0]                      AP_AXIMM_92_ARQOS,
    input wire                            AP_AXIMM_92_ARVALID,
    output  wire                            AP_AXIMM_92_ARREADY,
    output  wire [M_AXIMM_92_DATA_WIDTH-1:0]   AP_AXIMM_92_RDATA,
    output  wire [1:0]                      AP_AXIMM_92_RRESP,
    output  wire                            AP_AXIMM_92_RLAST,
    output  wire                            AP_AXIMM_92_RVALID,
    input  wire                            AP_AXIMM_92_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_92_AWADDR,
    output wire [7:0]                      M_AXIMM_92_AWLEN,
    output wire [2:0]                      M_AXIMM_92_AWSIZE,
    output wire [1:0]                      M_AXIMM_92_AWBURST,
    output wire [1:0]                      M_AXIMM_92_AWLOCK,
    output wire [3:0]                      M_AXIMM_92_AWCACHE,
    output wire [2:0]                      M_AXIMM_92_AWPROT,
    output wire [3:0]                      M_AXIMM_92_AWREGION,
    output wire [3:0]                      M_AXIMM_92_AWQOS,
    output wire                            M_AXIMM_92_AWVALID,
    input  wire                            M_AXIMM_92_AWREADY,
    output wire [M_AXIMM_92_DATA_WIDTH-1:0]   M_AXIMM_92_WDATA,
    output wire [M_AXIMM_92_DATA_WIDTH/8-1:0] M_AXIMM_92_WSTRB,
    output wire                            M_AXIMM_92_WLAST,
    output wire                            M_AXIMM_92_WVALID,
    input  wire                            M_AXIMM_92_WREADY,
    input  wire [1:0]                      M_AXIMM_92_BRESP,
    input  wire                            M_AXIMM_92_BVALID,
    output wire                            M_AXIMM_92_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_92_ARADDR,
    output wire [7:0]                      M_AXIMM_92_ARLEN,
    output wire [2:0]                      M_AXIMM_92_ARSIZE,
    output wire [1:0]                      M_AXIMM_92_ARBURST,
    output wire [1:0]                      M_AXIMM_92_ARLOCK,
    output wire [3:0]                      M_AXIMM_92_ARCACHE,
    output wire [2:0]                      M_AXIMM_92_ARPROT,
    output wire [3:0]                      M_AXIMM_92_ARREGION,
    output wire [3:0]                      M_AXIMM_92_ARQOS,
    output wire                            M_AXIMM_92_ARVALID,
    input  wire                            M_AXIMM_92_ARREADY,
    input  wire [M_AXIMM_92_DATA_WIDTH-1:0]   M_AXIMM_92_RDATA,
    input  wire [1:0]                      M_AXIMM_92_RRESP,
    input  wire                            M_AXIMM_92_RLAST,
    input  wire                            M_AXIMM_92_RVALID,
    output wire                            M_AXIMM_92_RREADY,
    //AXI-MM pass-through interface 93
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_93_AWADDR,
    input wire [7:0]                      AP_AXIMM_93_AWLEN,
    input wire [2:0]                      AP_AXIMM_93_AWSIZE,
    input wire [1:0]                      AP_AXIMM_93_AWBURST,
    input wire [1:0]                      AP_AXIMM_93_AWLOCK,
    input wire [3:0]                      AP_AXIMM_93_AWCACHE,
    input wire [2:0]                      AP_AXIMM_93_AWPROT,
    input wire [3:0]                      AP_AXIMM_93_AWREGION,
    input wire [3:0]                      AP_AXIMM_93_AWQOS,
    input wire                            AP_AXIMM_93_AWVALID,
    output  wire                            AP_AXIMM_93_AWREADY,
    input wire [M_AXIMM_93_DATA_WIDTH-1:0]   AP_AXIMM_93_WDATA,
    input wire [M_AXIMM_93_DATA_WIDTH/8-1:0] AP_AXIMM_93_WSTRB,
    input wire                            AP_AXIMM_93_WLAST,
    input wire                            AP_AXIMM_93_WVALID,
    output  wire                            AP_AXIMM_93_WREADY,
    output  wire [1:0]                      AP_AXIMM_93_BRESP,
    output  wire                            AP_AXIMM_93_BVALID,
    input wire                            AP_AXIMM_93_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_93_ARADDR,
    input wire [7:0]                      AP_AXIMM_93_ARLEN,
    input wire [2:0]                      AP_AXIMM_93_ARSIZE,
    input wire [1:0]                      AP_AXIMM_93_ARBURST,
    input wire [1:0]                      AP_AXIMM_93_ARLOCK,
    input wire [3:0]                      AP_AXIMM_93_ARCACHE,
    input wire [2:0]                      AP_AXIMM_93_ARPROT,
    input wire [3:0]                      AP_AXIMM_93_ARREGION,
    input wire [3:0]                      AP_AXIMM_93_ARQOS,
    input wire                            AP_AXIMM_93_ARVALID,
    output  wire                            AP_AXIMM_93_ARREADY,
    output  wire [M_AXIMM_93_DATA_WIDTH-1:0]   AP_AXIMM_93_RDATA,
    output  wire [1:0]                      AP_AXIMM_93_RRESP,
    output  wire                            AP_AXIMM_93_RLAST,
    output  wire                            AP_AXIMM_93_RVALID,
    input  wire                            AP_AXIMM_93_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_93_AWADDR,
    output wire [7:0]                      M_AXIMM_93_AWLEN,
    output wire [2:0]                      M_AXIMM_93_AWSIZE,
    output wire [1:0]                      M_AXIMM_93_AWBURST,
    output wire [1:0]                      M_AXIMM_93_AWLOCK,
    output wire [3:0]                      M_AXIMM_93_AWCACHE,
    output wire [2:0]                      M_AXIMM_93_AWPROT,
    output wire [3:0]                      M_AXIMM_93_AWREGION,
    output wire [3:0]                      M_AXIMM_93_AWQOS,
    output wire                            M_AXIMM_93_AWVALID,
    input  wire                            M_AXIMM_93_AWREADY,
    output wire [M_AXIMM_93_DATA_WIDTH-1:0]   M_AXIMM_93_WDATA,
    output wire [M_AXIMM_93_DATA_WIDTH/8-1:0] M_AXIMM_93_WSTRB,
    output wire                            M_AXIMM_93_WLAST,
    output wire                            M_AXIMM_93_WVALID,
    input  wire                            M_AXIMM_93_WREADY,
    input  wire [1:0]                      M_AXIMM_93_BRESP,
    input  wire                            M_AXIMM_93_BVALID,
    output wire                            M_AXIMM_93_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_93_ARADDR,
    output wire [7:0]                      M_AXIMM_93_ARLEN,
    output wire [2:0]                      M_AXIMM_93_ARSIZE,
    output wire [1:0]                      M_AXIMM_93_ARBURST,
    output wire [1:0]                      M_AXIMM_93_ARLOCK,
    output wire [3:0]                      M_AXIMM_93_ARCACHE,
    output wire [2:0]                      M_AXIMM_93_ARPROT,
    output wire [3:0]                      M_AXIMM_93_ARREGION,
    output wire [3:0]                      M_AXIMM_93_ARQOS,
    output wire                            M_AXIMM_93_ARVALID,
    input  wire                            M_AXIMM_93_ARREADY,
    input  wire [M_AXIMM_93_DATA_WIDTH-1:0]   M_AXIMM_93_RDATA,
    input  wire [1:0]                      M_AXIMM_93_RRESP,
    input  wire                            M_AXIMM_93_RLAST,
    input  wire                            M_AXIMM_93_RVALID,
    output wire                            M_AXIMM_93_RREADY,
    //AXI-MM pass-through interface 94
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_94_AWADDR,
    input wire [7:0]                      AP_AXIMM_94_AWLEN,
    input wire [2:0]                      AP_AXIMM_94_AWSIZE,
    input wire [1:0]                      AP_AXIMM_94_AWBURST,
    input wire [1:0]                      AP_AXIMM_94_AWLOCK,
    input wire [3:0]                      AP_AXIMM_94_AWCACHE,
    input wire [2:0]                      AP_AXIMM_94_AWPROT,
    input wire [3:0]                      AP_AXIMM_94_AWREGION,
    input wire [3:0]                      AP_AXIMM_94_AWQOS,
    input wire                            AP_AXIMM_94_AWVALID,
    output  wire                            AP_AXIMM_94_AWREADY,
    input wire [M_AXIMM_94_DATA_WIDTH-1:0]   AP_AXIMM_94_WDATA,
    input wire [M_AXIMM_94_DATA_WIDTH/8-1:0] AP_AXIMM_94_WSTRB,
    input wire                            AP_AXIMM_94_WLAST,
    input wire                            AP_AXIMM_94_WVALID,
    output  wire                            AP_AXIMM_94_WREADY,
    output  wire [1:0]                      AP_AXIMM_94_BRESP,
    output  wire                            AP_AXIMM_94_BVALID,
    input wire                            AP_AXIMM_94_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_94_ARADDR,
    input wire [7:0]                      AP_AXIMM_94_ARLEN,
    input wire [2:0]                      AP_AXIMM_94_ARSIZE,
    input wire [1:0]                      AP_AXIMM_94_ARBURST,
    input wire [1:0]                      AP_AXIMM_94_ARLOCK,
    input wire [3:0]                      AP_AXIMM_94_ARCACHE,
    input wire [2:0]                      AP_AXIMM_94_ARPROT,
    input wire [3:0]                      AP_AXIMM_94_ARREGION,
    input wire [3:0]                      AP_AXIMM_94_ARQOS,
    input wire                            AP_AXIMM_94_ARVALID,
    output  wire                            AP_AXIMM_94_ARREADY,
    output  wire [M_AXIMM_94_DATA_WIDTH-1:0]   AP_AXIMM_94_RDATA,
    output  wire [1:0]                      AP_AXIMM_94_RRESP,
    output  wire                            AP_AXIMM_94_RLAST,
    output  wire                            AP_AXIMM_94_RVALID,
    input  wire                            AP_AXIMM_94_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_94_AWADDR,
    output wire [7:0]                      M_AXIMM_94_AWLEN,
    output wire [2:0]                      M_AXIMM_94_AWSIZE,
    output wire [1:0]                      M_AXIMM_94_AWBURST,
    output wire [1:0]                      M_AXIMM_94_AWLOCK,
    output wire [3:0]                      M_AXIMM_94_AWCACHE,
    output wire [2:0]                      M_AXIMM_94_AWPROT,
    output wire [3:0]                      M_AXIMM_94_AWREGION,
    output wire [3:0]                      M_AXIMM_94_AWQOS,
    output wire                            M_AXIMM_94_AWVALID,
    input  wire                            M_AXIMM_94_AWREADY,
    output wire [M_AXIMM_94_DATA_WIDTH-1:0]   M_AXIMM_94_WDATA,
    output wire [M_AXIMM_94_DATA_WIDTH/8-1:0] M_AXIMM_94_WSTRB,
    output wire                            M_AXIMM_94_WLAST,
    output wire                            M_AXIMM_94_WVALID,
    input  wire                            M_AXIMM_94_WREADY,
    input  wire [1:0]                      M_AXIMM_94_BRESP,
    input  wire                            M_AXIMM_94_BVALID,
    output wire                            M_AXIMM_94_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_94_ARADDR,
    output wire [7:0]                      M_AXIMM_94_ARLEN,
    output wire [2:0]                      M_AXIMM_94_ARSIZE,
    output wire [1:0]                      M_AXIMM_94_ARBURST,
    output wire [1:0]                      M_AXIMM_94_ARLOCK,
    output wire [3:0]                      M_AXIMM_94_ARCACHE,
    output wire [2:0]                      M_AXIMM_94_ARPROT,
    output wire [3:0]                      M_AXIMM_94_ARREGION,
    output wire [3:0]                      M_AXIMM_94_ARQOS,
    output wire                            M_AXIMM_94_ARVALID,
    input  wire                            M_AXIMM_94_ARREADY,
    input  wire [M_AXIMM_94_DATA_WIDTH-1:0]   M_AXIMM_94_RDATA,
    input  wire [1:0]                      M_AXIMM_94_RRESP,
    input  wire                            M_AXIMM_94_RLAST,
    input  wire                            M_AXIMM_94_RVALID,
    output wire                            M_AXIMM_94_RREADY,
    //AXI-MM pass-through interface 95
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_95_AWADDR,
    input wire [7:0]                      AP_AXIMM_95_AWLEN,
    input wire [2:0]                      AP_AXIMM_95_AWSIZE,
    input wire [1:0]                      AP_AXIMM_95_AWBURST,
    input wire [1:0]                      AP_AXIMM_95_AWLOCK,
    input wire [3:0]                      AP_AXIMM_95_AWCACHE,
    input wire [2:0]                      AP_AXIMM_95_AWPROT,
    input wire [3:0]                      AP_AXIMM_95_AWREGION,
    input wire [3:0]                      AP_AXIMM_95_AWQOS,
    input wire                            AP_AXIMM_95_AWVALID,
    output  wire                            AP_AXIMM_95_AWREADY,
    input wire [M_AXIMM_95_DATA_WIDTH-1:0]   AP_AXIMM_95_WDATA,
    input wire [M_AXIMM_95_DATA_WIDTH/8-1:0] AP_AXIMM_95_WSTRB,
    input wire                            AP_AXIMM_95_WLAST,
    input wire                            AP_AXIMM_95_WVALID,
    output  wire                            AP_AXIMM_95_WREADY,
    output  wire [1:0]                      AP_AXIMM_95_BRESP,
    output  wire                            AP_AXIMM_95_BVALID,
    input wire                            AP_AXIMM_95_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_95_ARADDR,
    input wire [7:0]                      AP_AXIMM_95_ARLEN,
    input wire [2:0]                      AP_AXIMM_95_ARSIZE,
    input wire [1:0]                      AP_AXIMM_95_ARBURST,
    input wire [1:0]                      AP_AXIMM_95_ARLOCK,
    input wire [3:0]                      AP_AXIMM_95_ARCACHE,
    input wire [2:0]                      AP_AXIMM_95_ARPROT,
    input wire [3:0]                      AP_AXIMM_95_ARREGION,
    input wire [3:0]                      AP_AXIMM_95_ARQOS,
    input wire                            AP_AXIMM_95_ARVALID,
    output  wire                            AP_AXIMM_95_ARREADY,
    output  wire [M_AXIMM_95_DATA_WIDTH-1:0]   AP_AXIMM_95_RDATA,
    output  wire [1:0]                      AP_AXIMM_95_RRESP,
    output  wire                            AP_AXIMM_95_RLAST,
    output  wire                            AP_AXIMM_95_RVALID,
    input  wire                            AP_AXIMM_95_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_95_AWADDR,
    output wire [7:0]                      M_AXIMM_95_AWLEN,
    output wire [2:0]                      M_AXIMM_95_AWSIZE,
    output wire [1:0]                      M_AXIMM_95_AWBURST,
    output wire [1:0]                      M_AXIMM_95_AWLOCK,
    output wire [3:0]                      M_AXIMM_95_AWCACHE,
    output wire [2:0]                      M_AXIMM_95_AWPROT,
    output wire [3:0]                      M_AXIMM_95_AWREGION,
    output wire [3:0]                      M_AXIMM_95_AWQOS,
    output wire                            M_AXIMM_95_AWVALID,
    input  wire                            M_AXIMM_95_AWREADY,
    output wire [M_AXIMM_95_DATA_WIDTH-1:0]   M_AXIMM_95_WDATA,
    output wire [M_AXIMM_95_DATA_WIDTH/8-1:0] M_AXIMM_95_WSTRB,
    output wire                            M_AXIMM_95_WLAST,
    output wire                            M_AXIMM_95_WVALID,
    input  wire                            M_AXIMM_95_WREADY,
    input  wire [1:0]                      M_AXIMM_95_BRESP,
    input  wire                            M_AXIMM_95_BVALID,
    output wire                            M_AXIMM_95_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_95_ARADDR,
    output wire [7:0]                      M_AXIMM_95_ARLEN,
    output wire [2:0]                      M_AXIMM_95_ARSIZE,
    output wire [1:0]                      M_AXIMM_95_ARBURST,
    output wire [1:0]                      M_AXIMM_95_ARLOCK,
    output wire [3:0]                      M_AXIMM_95_ARCACHE,
    output wire [2:0]                      M_AXIMM_95_ARPROT,
    output wire [3:0]                      M_AXIMM_95_ARREGION,
    output wire [3:0]                      M_AXIMM_95_ARQOS,
    output wire                            M_AXIMM_95_ARVALID,
    input  wire                            M_AXIMM_95_ARREADY,
    input  wire [M_AXIMM_95_DATA_WIDTH-1:0]   M_AXIMM_95_RDATA,
    input  wire [1:0]                      M_AXIMM_95_RRESP,
    input  wire                            M_AXIMM_95_RLAST,
    input  wire                            M_AXIMM_95_RVALID,
    output wire                            M_AXIMM_95_RREADY,
    //AXI-MM pass-through interface 96
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_96_AWADDR,
    input wire [7:0]                      AP_AXIMM_96_AWLEN,
    input wire [2:0]                      AP_AXIMM_96_AWSIZE,
    input wire [1:0]                      AP_AXIMM_96_AWBURST,
    input wire [1:0]                      AP_AXIMM_96_AWLOCK,
    input wire [3:0]                      AP_AXIMM_96_AWCACHE,
    input wire [2:0]                      AP_AXIMM_96_AWPROT,
    input wire [3:0]                      AP_AXIMM_96_AWREGION,
    input wire [3:0]                      AP_AXIMM_96_AWQOS,
    input wire                            AP_AXIMM_96_AWVALID,
    output  wire                            AP_AXIMM_96_AWREADY,
    input wire [M_AXIMM_96_DATA_WIDTH-1:0]   AP_AXIMM_96_WDATA,
    input wire [M_AXIMM_96_DATA_WIDTH/8-1:0] AP_AXIMM_96_WSTRB,
    input wire                            AP_AXIMM_96_WLAST,
    input wire                            AP_AXIMM_96_WVALID,
    output  wire                            AP_AXIMM_96_WREADY,
    output  wire [1:0]                      AP_AXIMM_96_BRESP,
    output  wire                            AP_AXIMM_96_BVALID,
    input wire                            AP_AXIMM_96_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_96_ARADDR,
    input wire [7:0]                      AP_AXIMM_96_ARLEN,
    input wire [2:0]                      AP_AXIMM_96_ARSIZE,
    input wire [1:0]                      AP_AXIMM_96_ARBURST,
    input wire [1:0]                      AP_AXIMM_96_ARLOCK,
    input wire [3:0]                      AP_AXIMM_96_ARCACHE,
    input wire [2:0]                      AP_AXIMM_96_ARPROT,
    input wire [3:0]                      AP_AXIMM_96_ARREGION,
    input wire [3:0]                      AP_AXIMM_96_ARQOS,
    input wire                            AP_AXIMM_96_ARVALID,
    output  wire                            AP_AXIMM_96_ARREADY,
    output  wire [M_AXIMM_96_DATA_WIDTH-1:0]   AP_AXIMM_96_RDATA,
    output  wire [1:0]                      AP_AXIMM_96_RRESP,
    output  wire                            AP_AXIMM_96_RLAST,
    output  wire                            AP_AXIMM_96_RVALID,
    input  wire                            AP_AXIMM_96_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_96_AWADDR,
    output wire [7:0]                      M_AXIMM_96_AWLEN,
    output wire [2:0]                      M_AXIMM_96_AWSIZE,
    output wire [1:0]                      M_AXIMM_96_AWBURST,
    output wire [1:0]                      M_AXIMM_96_AWLOCK,
    output wire [3:0]                      M_AXIMM_96_AWCACHE,
    output wire [2:0]                      M_AXIMM_96_AWPROT,
    output wire [3:0]                      M_AXIMM_96_AWREGION,
    output wire [3:0]                      M_AXIMM_96_AWQOS,
    output wire                            M_AXIMM_96_AWVALID,
    input  wire                            M_AXIMM_96_AWREADY,
    output wire [M_AXIMM_96_DATA_WIDTH-1:0]   M_AXIMM_96_WDATA,
    output wire [M_AXIMM_96_DATA_WIDTH/8-1:0] M_AXIMM_96_WSTRB,
    output wire                            M_AXIMM_96_WLAST,
    output wire                            M_AXIMM_96_WVALID,
    input  wire                            M_AXIMM_96_WREADY,
    input  wire [1:0]                      M_AXIMM_96_BRESP,
    input  wire                            M_AXIMM_96_BVALID,
    output wire                            M_AXIMM_96_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_96_ARADDR,
    output wire [7:0]                      M_AXIMM_96_ARLEN,
    output wire [2:0]                      M_AXIMM_96_ARSIZE,
    output wire [1:0]                      M_AXIMM_96_ARBURST,
    output wire [1:0]                      M_AXIMM_96_ARLOCK,
    output wire [3:0]                      M_AXIMM_96_ARCACHE,
    output wire [2:0]                      M_AXIMM_96_ARPROT,
    output wire [3:0]                      M_AXIMM_96_ARREGION,
    output wire [3:0]                      M_AXIMM_96_ARQOS,
    output wire                            M_AXIMM_96_ARVALID,
    input  wire                            M_AXIMM_96_ARREADY,
    input  wire [M_AXIMM_96_DATA_WIDTH-1:0]   M_AXIMM_96_RDATA,
    input  wire [1:0]                      M_AXIMM_96_RRESP,
    input  wire                            M_AXIMM_96_RLAST,
    input  wire                            M_AXIMM_96_RVALID,
    output wire                            M_AXIMM_96_RREADY,
    //AXI-MM pass-through interface 97
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_97_AWADDR,
    input wire [7:0]                      AP_AXIMM_97_AWLEN,
    input wire [2:0]                      AP_AXIMM_97_AWSIZE,
    input wire [1:0]                      AP_AXIMM_97_AWBURST,
    input wire [1:0]                      AP_AXIMM_97_AWLOCK,
    input wire [3:0]                      AP_AXIMM_97_AWCACHE,
    input wire [2:0]                      AP_AXIMM_97_AWPROT,
    input wire [3:0]                      AP_AXIMM_97_AWREGION,
    input wire [3:0]                      AP_AXIMM_97_AWQOS,
    input wire                            AP_AXIMM_97_AWVALID,
    output  wire                            AP_AXIMM_97_AWREADY,
    input wire [M_AXIMM_97_DATA_WIDTH-1:0]   AP_AXIMM_97_WDATA,
    input wire [M_AXIMM_97_DATA_WIDTH/8-1:0] AP_AXIMM_97_WSTRB,
    input wire                            AP_AXIMM_97_WLAST,
    input wire                            AP_AXIMM_97_WVALID,
    output  wire                            AP_AXIMM_97_WREADY,
    output  wire [1:0]                      AP_AXIMM_97_BRESP,
    output  wire                            AP_AXIMM_97_BVALID,
    input wire                            AP_AXIMM_97_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_97_ARADDR,
    input wire [7:0]                      AP_AXIMM_97_ARLEN,
    input wire [2:0]                      AP_AXIMM_97_ARSIZE,
    input wire [1:0]                      AP_AXIMM_97_ARBURST,
    input wire [1:0]                      AP_AXIMM_97_ARLOCK,
    input wire [3:0]                      AP_AXIMM_97_ARCACHE,
    input wire [2:0]                      AP_AXIMM_97_ARPROT,
    input wire [3:0]                      AP_AXIMM_97_ARREGION,
    input wire [3:0]                      AP_AXIMM_97_ARQOS,
    input wire                            AP_AXIMM_97_ARVALID,
    output  wire                            AP_AXIMM_97_ARREADY,
    output  wire [M_AXIMM_97_DATA_WIDTH-1:0]   AP_AXIMM_97_RDATA,
    output  wire [1:0]                      AP_AXIMM_97_RRESP,
    output  wire                            AP_AXIMM_97_RLAST,
    output  wire                            AP_AXIMM_97_RVALID,
    input  wire                            AP_AXIMM_97_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_97_AWADDR,
    output wire [7:0]                      M_AXIMM_97_AWLEN,
    output wire [2:0]                      M_AXIMM_97_AWSIZE,
    output wire [1:0]                      M_AXIMM_97_AWBURST,
    output wire [1:0]                      M_AXIMM_97_AWLOCK,
    output wire [3:0]                      M_AXIMM_97_AWCACHE,
    output wire [2:0]                      M_AXIMM_97_AWPROT,
    output wire [3:0]                      M_AXIMM_97_AWREGION,
    output wire [3:0]                      M_AXIMM_97_AWQOS,
    output wire                            M_AXIMM_97_AWVALID,
    input  wire                            M_AXIMM_97_AWREADY,
    output wire [M_AXIMM_97_DATA_WIDTH-1:0]   M_AXIMM_97_WDATA,
    output wire [M_AXIMM_97_DATA_WIDTH/8-1:0] M_AXIMM_97_WSTRB,
    output wire                            M_AXIMM_97_WLAST,
    output wire                            M_AXIMM_97_WVALID,
    input  wire                            M_AXIMM_97_WREADY,
    input  wire [1:0]                      M_AXIMM_97_BRESP,
    input  wire                            M_AXIMM_97_BVALID,
    output wire                            M_AXIMM_97_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_97_ARADDR,
    output wire [7:0]                      M_AXIMM_97_ARLEN,
    output wire [2:0]                      M_AXIMM_97_ARSIZE,
    output wire [1:0]                      M_AXIMM_97_ARBURST,
    output wire [1:0]                      M_AXIMM_97_ARLOCK,
    output wire [3:0]                      M_AXIMM_97_ARCACHE,
    output wire [2:0]                      M_AXIMM_97_ARPROT,
    output wire [3:0]                      M_AXIMM_97_ARREGION,
    output wire [3:0]                      M_AXIMM_97_ARQOS,
    output wire                            M_AXIMM_97_ARVALID,
    input  wire                            M_AXIMM_97_ARREADY,
    input  wire [M_AXIMM_97_DATA_WIDTH-1:0]   M_AXIMM_97_RDATA,
    input  wire [1:0]                      M_AXIMM_97_RRESP,
    input  wire                            M_AXIMM_97_RLAST,
    input  wire                            M_AXIMM_97_RVALID,
    output wire                            M_AXIMM_97_RREADY,
    //AXI-MM pass-through interface 98
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_98_AWADDR,
    input wire [7:0]                      AP_AXIMM_98_AWLEN,
    input wire [2:0]                      AP_AXIMM_98_AWSIZE,
    input wire [1:0]                      AP_AXIMM_98_AWBURST,
    input wire [1:0]                      AP_AXIMM_98_AWLOCK,
    input wire [3:0]                      AP_AXIMM_98_AWCACHE,
    input wire [2:0]                      AP_AXIMM_98_AWPROT,
    input wire [3:0]                      AP_AXIMM_98_AWREGION,
    input wire [3:0]                      AP_AXIMM_98_AWQOS,
    input wire                            AP_AXIMM_98_AWVALID,
    output  wire                            AP_AXIMM_98_AWREADY,
    input wire [M_AXIMM_98_DATA_WIDTH-1:0]   AP_AXIMM_98_WDATA,
    input wire [M_AXIMM_98_DATA_WIDTH/8-1:0] AP_AXIMM_98_WSTRB,
    input wire                            AP_AXIMM_98_WLAST,
    input wire                            AP_AXIMM_98_WVALID,
    output  wire                            AP_AXIMM_98_WREADY,
    output  wire [1:0]                      AP_AXIMM_98_BRESP,
    output  wire                            AP_AXIMM_98_BVALID,
    input wire                            AP_AXIMM_98_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_98_ARADDR,
    input wire [7:0]                      AP_AXIMM_98_ARLEN,
    input wire [2:0]                      AP_AXIMM_98_ARSIZE,
    input wire [1:0]                      AP_AXIMM_98_ARBURST,
    input wire [1:0]                      AP_AXIMM_98_ARLOCK,
    input wire [3:0]                      AP_AXIMM_98_ARCACHE,
    input wire [2:0]                      AP_AXIMM_98_ARPROT,
    input wire [3:0]                      AP_AXIMM_98_ARREGION,
    input wire [3:0]                      AP_AXIMM_98_ARQOS,
    input wire                            AP_AXIMM_98_ARVALID,
    output  wire                            AP_AXIMM_98_ARREADY,
    output  wire [M_AXIMM_98_DATA_WIDTH-1:0]   AP_AXIMM_98_RDATA,
    output  wire [1:0]                      AP_AXIMM_98_RRESP,
    output  wire                            AP_AXIMM_98_RLAST,
    output  wire                            AP_AXIMM_98_RVALID,
    input  wire                            AP_AXIMM_98_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_98_AWADDR,
    output wire [7:0]                      M_AXIMM_98_AWLEN,
    output wire [2:0]                      M_AXIMM_98_AWSIZE,
    output wire [1:0]                      M_AXIMM_98_AWBURST,
    output wire [1:0]                      M_AXIMM_98_AWLOCK,
    output wire [3:0]                      M_AXIMM_98_AWCACHE,
    output wire [2:0]                      M_AXIMM_98_AWPROT,
    output wire [3:0]                      M_AXIMM_98_AWREGION,
    output wire [3:0]                      M_AXIMM_98_AWQOS,
    output wire                            M_AXIMM_98_AWVALID,
    input  wire                            M_AXIMM_98_AWREADY,
    output wire [M_AXIMM_98_DATA_WIDTH-1:0]   M_AXIMM_98_WDATA,
    output wire [M_AXIMM_98_DATA_WIDTH/8-1:0] M_AXIMM_98_WSTRB,
    output wire                            M_AXIMM_98_WLAST,
    output wire                            M_AXIMM_98_WVALID,
    input  wire                            M_AXIMM_98_WREADY,
    input  wire [1:0]                      M_AXIMM_98_BRESP,
    input  wire                            M_AXIMM_98_BVALID,
    output wire                            M_AXIMM_98_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_98_ARADDR,
    output wire [7:0]                      M_AXIMM_98_ARLEN,
    output wire [2:0]                      M_AXIMM_98_ARSIZE,
    output wire [1:0]                      M_AXIMM_98_ARBURST,
    output wire [1:0]                      M_AXIMM_98_ARLOCK,
    output wire [3:0]                      M_AXIMM_98_ARCACHE,
    output wire [2:0]                      M_AXIMM_98_ARPROT,
    output wire [3:0]                      M_AXIMM_98_ARREGION,
    output wire [3:0]                      M_AXIMM_98_ARQOS,
    output wire                            M_AXIMM_98_ARVALID,
    input  wire                            M_AXIMM_98_ARREADY,
    input  wire [M_AXIMM_98_DATA_WIDTH-1:0]   M_AXIMM_98_RDATA,
    input  wire [1:0]                      M_AXIMM_98_RRESP,
    input  wire                            M_AXIMM_98_RLAST,
    input  wire                            M_AXIMM_98_RVALID,
    output wire                            M_AXIMM_98_RREADY,
    //AXI-MM pass-through interface 99
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_99_AWADDR,
    input wire [7:0]                      AP_AXIMM_99_AWLEN,
    input wire [2:0]                      AP_AXIMM_99_AWSIZE,
    input wire [1:0]                      AP_AXIMM_99_AWBURST,
    input wire [1:0]                      AP_AXIMM_99_AWLOCK,
    input wire [3:0]                      AP_AXIMM_99_AWCACHE,
    input wire [2:0]                      AP_AXIMM_99_AWPROT,
    input wire [3:0]                      AP_AXIMM_99_AWREGION,
    input wire [3:0]                      AP_AXIMM_99_AWQOS,
    input wire                            AP_AXIMM_99_AWVALID,
    output  wire                            AP_AXIMM_99_AWREADY,
    input wire [M_AXIMM_99_DATA_WIDTH-1:0]   AP_AXIMM_99_WDATA,
    input wire [M_AXIMM_99_DATA_WIDTH/8-1:0] AP_AXIMM_99_WSTRB,
    input wire                            AP_AXIMM_99_WLAST,
    input wire                            AP_AXIMM_99_WVALID,
    output  wire                            AP_AXIMM_99_WREADY,
    output  wire [1:0]                      AP_AXIMM_99_BRESP,
    output  wire                            AP_AXIMM_99_BVALID,
    input wire                            AP_AXIMM_99_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_99_ARADDR,
    input wire [7:0]                      AP_AXIMM_99_ARLEN,
    input wire [2:0]                      AP_AXIMM_99_ARSIZE,
    input wire [1:0]                      AP_AXIMM_99_ARBURST,
    input wire [1:0]                      AP_AXIMM_99_ARLOCK,
    input wire [3:0]                      AP_AXIMM_99_ARCACHE,
    input wire [2:0]                      AP_AXIMM_99_ARPROT,
    input wire [3:0]                      AP_AXIMM_99_ARREGION,
    input wire [3:0]                      AP_AXIMM_99_ARQOS,
    input wire                            AP_AXIMM_99_ARVALID,
    output  wire                            AP_AXIMM_99_ARREADY,
    output  wire [M_AXIMM_99_DATA_WIDTH-1:0]   AP_AXIMM_99_RDATA,
    output  wire [1:0]                      AP_AXIMM_99_RRESP,
    output  wire                            AP_AXIMM_99_RLAST,
    output  wire                            AP_AXIMM_99_RVALID,
    input  wire                            AP_AXIMM_99_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_99_AWADDR,
    output wire [7:0]                      M_AXIMM_99_AWLEN,
    output wire [2:0]                      M_AXIMM_99_AWSIZE,
    output wire [1:0]                      M_AXIMM_99_AWBURST,
    output wire [1:0]                      M_AXIMM_99_AWLOCK,
    output wire [3:0]                      M_AXIMM_99_AWCACHE,
    output wire [2:0]                      M_AXIMM_99_AWPROT,
    output wire [3:0]                      M_AXIMM_99_AWREGION,
    output wire [3:0]                      M_AXIMM_99_AWQOS,
    output wire                            M_AXIMM_99_AWVALID,
    input  wire                            M_AXIMM_99_AWREADY,
    output wire [M_AXIMM_99_DATA_WIDTH-1:0]   M_AXIMM_99_WDATA,
    output wire [M_AXIMM_99_DATA_WIDTH/8-1:0] M_AXIMM_99_WSTRB,
    output wire                            M_AXIMM_99_WLAST,
    output wire                            M_AXIMM_99_WVALID,
    input  wire                            M_AXIMM_99_WREADY,
    input  wire [1:0]                      M_AXIMM_99_BRESP,
    input  wire                            M_AXIMM_99_BVALID,
    output wire                            M_AXIMM_99_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_99_ARADDR,
    output wire [7:0]                      M_AXIMM_99_ARLEN,
    output wire [2:0]                      M_AXIMM_99_ARSIZE,
    output wire [1:0]                      M_AXIMM_99_ARBURST,
    output wire [1:0]                      M_AXIMM_99_ARLOCK,
    output wire [3:0]                      M_AXIMM_99_ARCACHE,
    output wire [2:0]                      M_AXIMM_99_ARPROT,
    output wire [3:0]                      M_AXIMM_99_ARREGION,
    output wire [3:0]                      M_AXIMM_99_ARQOS,
    output wire                            M_AXIMM_99_ARVALID,
    input  wire                            M_AXIMM_99_ARREADY,
    input  wire [M_AXIMM_99_DATA_WIDTH-1:0]   M_AXIMM_99_RDATA,
    input  wire [1:0]                      M_AXIMM_99_RRESP,
    input  wire                            M_AXIMM_99_RLAST,
    input  wire                            M_AXIMM_99_RVALID,
    output wire                            M_AXIMM_99_RREADY,
    //AXI-MM pass-through interface 100
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_100_AWADDR,
    input wire [7:0]                      AP_AXIMM_100_AWLEN,
    input wire [2:0]                      AP_AXIMM_100_AWSIZE,
    input wire [1:0]                      AP_AXIMM_100_AWBURST,
    input wire [1:0]                      AP_AXIMM_100_AWLOCK,
    input wire [3:0]                      AP_AXIMM_100_AWCACHE,
    input wire [2:0]                      AP_AXIMM_100_AWPROT,
    input wire [3:0]                      AP_AXIMM_100_AWREGION,
    input wire [3:0]                      AP_AXIMM_100_AWQOS,
    input wire                            AP_AXIMM_100_AWVALID,
    output  wire                            AP_AXIMM_100_AWREADY,
    input wire [M_AXIMM_100_DATA_WIDTH-1:0]   AP_AXIMM_100_WDATA,
    input wire [M_AXIMM_100_DATA_WIDTH/8-1:0] AP_AXIMM_100_WSTRB,
    input wire                            AP_AXIMM_100_WLAST,
    input wire                            AP_AXIMM_100_WVALID,
    output  wire                            AP_AXIMM_100_WREADY,
    output  wire [1:0]                      AP_AXIMM_100_BRESP,
    output  wire                            AP_AXIMM_100_BVALID,
    input wire                            AP_AXIMM_100_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_100_ARADDR,
    input wire [7:0]                      AP_AXIMM_100_ARLEN,
    input wire [2:0]                      AP_AXIMM_100_ARSIZE,
    input wire [1:0]                      AP_AXIMM_100_ARBURST,
    input wire [1:0]                      AP_AXIMM_100_ARLOCK,
    input wire [3:0]                      AP_AXIMM_100_ARCACHE,
    input wire [2:0]                      AP_AXIMM_100_ARPROT,
    input wire [3:0]                      AP_AXIMM_100_ARREGION,
    input wire [3:0]                      AP_AXIMM_100_ARQOS,
    input wire                            AP_AXIMM_100_ARVALID,
    output  wire                            AP_AXIMM_100_ARREADY,
    output  wire [M_AXIMM_100_DATA_WIDTH-1:0]   AP_AXIMM_100_RDATA,
    output  wire [1:0]                      AP_AXIMM_100_RRESP,
    output  wire                            AP_AXIMM_100_RLAST,
    output  wire                            AP_AXIMM_100_RVALID,
    input  wire                            AP_AXIMM_100_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_100_AWADDR,
    output wire [7:0]                      M_AXIMM_100_AWLEN,
    output wire [2:0]                      M_AXIMM_100_AWSIZE,
    output wire [1:0]                      M_AXIMM_100_AWBURST,
    output wire [1:0]                      M_AXIMM_100_AWLOCK,
    output wire [3:0]                      M_AXIMM_100_AWCACHE,
    output wire [2:0]                      M_AXIMM_100_AWPROT,
    output wire [3:0]                      M_AXIMM_100_AWREGION,
    output wire [3:0]                      M_AXIMM_100_AWQOS,
    output wire                            M_AXIMM_100_AWVALID,
    input  wire                            M_AXIMM_100_AWREADY,
    output wire [M_AXIMM_100_DATA_WIDTH-1:0]   M_AXIMM_100_WDATA,
    output wire [M_AXIMM_100_DATA_WIDTH/8-1:0] M_AXIMM_100_WSTRB,
    output wire                            M_AXIMM_100_WLAST,
    output wire                            M_AXIMM_100_WVALID,
    input  wire                            M_AXIMM_100_WREADY,
    input  wire [1:0]                      M_AXIMM_100_BRESP,
    input  wire                            M_AXIMM_100_BVALID,
    output wire                            M_AXIMM_100_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_100_ARADDR,
    output wire [7:0]                      M_AXIMM_100_ARLEN,
    output wire [2:0]                      M_AXIMM_100_ARSIZE,
    output wire [1:0]                      M_AXIMM_100_ARBURST,
    output wire [1:0]                      M_AXIMM_100_ARLOCK,
    output wire [3:0]                      M_AXIMM_100_ARCACHE,
    output wire [2:0]                      M_AXIMM_100_ARPROT,
    output wire [3:0]                      M_AXIMM_100_ARREGION,
    output wire [3:0]                      M_AXIMM_100_ARQOS,
    output wire                            M_AXIMM_100_ARVALID,
    input  wire                            M_AXIMM_100_ARREADY,
    input  wire [M_AXIMM_100_DATA_WIDTH-1:0]   M_AXIMM_100_RDATA,
    input  wire [1:0]                      M_AXIMM_100_RRESP,
    input  wire                            M_AXIMM_100_RLAST,
    input  wire                            M_AXIMM_100_RVALID,
    output wire                            M_AXIMM_100_RREADY,
    //AXI-MM pass-through interface 101
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_101_AWADDR,
    input wire [7:0]                      AP_AXIMM_101_AWLEN,
    input wire [2:0]                      AP_AXIMM_101_AWSIZE,
    input wire [1:0]                      AP_AXIMM_101_AWBURST,
    input wire [1:0]                      AP_AXIMM_101_AWLOCK,
    input wire [3:0]                      AP_AXIMM_101_AWCACHE,
    input wire [2:0]                      AP_AXIMM_101_AWPROT,
    input wire [3:0]                      AP_AXIMM_101_AWREGION,
    input wire [3:0]                      AP_AXIMM_101_AWQOS,
    input wire                            AP_AXIMM_101_AWVALID,
    output  wire                            AP_AXIMM_101_AWREADY,
    input wire [M_AXIMM_101_DATA_WIDTH-1:0]   AP_AXIMM_101_WDATA,
    input wire [M_AXIMM_101_DATA_WIDTH/8-1:0] AP_AXIMM_101_WSTRB,
    input wire                            AP_AXIMM_101_WLAST,
    input wire                            AP_AXIMM_101_WVALID,
    output  wire                            AP_AXIMM_101_WREADY,
    output  wire [1:0]                      AP_AXIMM_101_BRESP,
    output  wire                            AP_AXIMM_101_BVALID,
    input wire                            AP_AXIMM_101_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_101_ARADDR,
    input wire [7:0]                      AP_AXIMM_101_ARLEN,
    input wire [2:0]                      AP_AXIMM_101_ARSIZE,
    input wire [1:0]                      AP_AXIMM_101_ARBURST,
    input wire [1:0]                      AP_AXIMM_101_ARLOCK,
    input wire [3:0]                      AP_AXIMM_101_ARCACHE,
    input wire [2:0]                      AP_AXIMM_101_ARPROT,
    input wire [3:0]                      AP_AXIMM_101_ARREGION,
    input wire [3:0]                      AP_AXIMM_101_ARQOS,
    input wire                            AP_AXIMM_101_ARVALID,
    output  wire                            AP_AXIMM_101_ARREADY,
    output  wire [M_AXIMM_101_DATA_WIDTH-1:0]   AP_AXIMM_101_RDATA,
    output  wire [1:0]                      AP_AXIMM_101_RRESP,
    output  wire                            AP_AXIMM_101_RLAST,
    output  wire                            AP_AXIMM_101_RVALID,
    input  wire                            AP_AXIMM_101_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_101_AWADDR,
    output wire [7:0]                      M_AXIMM_101_AWLEN,
    output wire [2:0]                      M_AXIMM_101_AWSIZE,
    output wire [1:0]                      M_AXIMM_101_AWBURST,
    output wire [1:0]                      M_AXIMM_101_AWLOCK,
    output wire [3:0]                      M_AXIMM_101_AWCACHE,
    output wire [2:0]                      M_AXIMM_101_AWPROT,
    output wire [3:0]                      M_AXIMM_101_AWREGION,
    output wire [3:0]                      M_AXIMM_101_AWQOS,
    output wire                            M_AXIMM_101_AWVALID,
    input  wire                            M_AXIMM_101_AWREADY,
    output wire [M_AXIMM_101_DATA_WIDTH-1:0]   M_AXIMM_101_WDATA,
    output wire [M_AXIMM_101_DATA_WIDTH/8-1:0] M_AXIMM_101_WSTRB,
    output wire                            M_AXIMM_101_WLAST,
    output wire                            M_AXIMM_101_WVALID,
    input  wire                            M_AXIMM_101_WREADY,
    input  wire [1:0]                      M_AXIMM_101_BRESP,
    input  wire                            M_AXIMM_101_BVALID,
    output wire                            M_AXIMM_101_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_101_ARADDR,
    output wire [7:0]                      M_AXIMM_101_ARLEN,
    output wire [2:0]                      M_AXIMM_101_ARSIZE,
    output wire [1:0]                      M_AXIMM_101_ARBURST,
    output wire [1:0]                      M_AXIMM_101_ARLOCK,
    output wire [3:0]                      M_AXIMM_101_ARCACHE,
    output wire [2:0]                      M_AXIMM_101_ARPROT,
    output wire [3:0]                      M_AXIMM_101_ARREGION,
    output wire [3:0]                      M_AXIMM_101_ARQOS,
    output wire                            M_AXIMM_101_ARVALID,
    input  wire                            M_AXIMM_101_ARREADY,
    input  wire [M_AXIMM_101_DATA_WIDTH-1:0]   M_AXIMM_101_RDATA,
    input  wire [1:0]                      M_AXIMM_101_RRESP,
    input  wire                            M_AXIMM_101_RLAST,
    input  wire                            M_AXIMM_101_RVALID,
    output wire                            M_AXIMM_101_RREADY,
    //AXI-MM pass-through interface 102
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_102_AWADDR,
    input wire [7:0]                      AP_AXIMM_102_AWLEN,
    input wire [2:0]                      AP_AXIMM_102_AWSIZE,
    input wire [1:0]                      AP_AXIMM_102_AWBURST,
    input wire [1:0]                      AP_AXIMM_102_AWLOCK,
    input wire [3:0]                      AP_AXIMM_102_AWCACHE,
    input wire [2:0]                      AP_AXIMM_102_AWPROT,
    input wire [3:0]                      AP_AXIMM_102_AWREGION,
    input wire [3:0]                      AP_AXIMM_102_AWQOS,
    input wire                            AP_AXIMM_102_AWVALID,
    output  wire                            AP_AXIMM_102_AWREADY,
    input wire [M_AXIMM_102_DATA_WIDTH-1:0]   AP_AXIMM_102_WDATA,
    input wire [M_AXIMM_102_DATA_WIDTH/8-1:0] AP_AXIMM_102_WSTRB,
    input wire                            AP_AXIMM_102_WLAST,
    input wire                            AP_AXIMM_102_WVALID,
    output  wire                            AP_AXIMM_102_WREADY,
    output  wire [1:0]                      AP_AXIMM_102_BRESP,
    output  wire                            AP_AXIMM_102_BVALID,
    input wire                            AP_AXIMM_102_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_102_ARADDR,
    input wire [7:0]                      AP_AXIMM_102_ARLEN,
    input wire [2:0]                      AP_AXIMM_102_ARSIZE,
    input wire [1:0]                      AP_AXIMM_102_ARBURST,
    input wire [1:0]                      AP_AXIMM_102_ARLOCK,
    input wire [3:0]                      AP_AXIMM_102_ARCACHE,
    input wire [2:0]                      AP_AXIMM_102_ARPROT,
    input wire [3:0]                      AP_AXIMM_102_ARREGION,
    input wire [3:0]                      AP_AXIMM_102_ARQOS,
    input wire                            AP_AXIMM_102_ARVALID,
    output  wire                            AP_AXIMM_102_ARREADY,
    output  wire [M_AXIMM_102_DATA_WIDTH-1:0]   AP_AXIMM_102_RDATA,
    output  wire [1:0]                      AP_AXIMM_102_RRESP,
    output  wire                            AP_AXIMM_102_RLAST,
    output  wire                            AP_AXIMM_102_RVALID,
    input  wire                            AP_AXIMM_102_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_102_AWADDR,
    output wire [7:0]                      M_AXIMM_102_AWLEN,
    output wire [2:0]                      M_AXIMM_102_AWSIZE,
    output wire [1:0]                      M_AXIMM_102_AWBURST,
    output wire [1:0]                      M_AXIMM_102_AWLOCK,
    output wire [3:0]                      M_AXIMM_102_AWCACHE,
    output wire [2:0]                      M_AXIMM_102_AWPROT,
    output wire [3:0]                      M_AXIMM_102_AWREGION,
    output wire [3:0]                      M_AXIMM_102_AWQOS,
    output wire                            M_AXIMM_102_AWVALID,
    input  wire                            M_AXIMM_102_AWREADY,
    output wire [M_AXIMM_102_DATA_WIDTH-1:0]   M_AXIMM_102_WDATA,
    output wire [M_AXIMM_102_DATA_WIDTH/8-1:0] M_AXIMM_102_WSTRB,
    output wire                            M_AXIMM_102_WLAST,
    output wire                            M_AXIMM_102_WVALID,
    input  wire                            M_AXIMM_102_WREADY,
    input  wire [1:0]                      M_AXIMM_102_BRESP,
    input  wire                            M_AXIMM_102_BVALID,
    output wire                            M_AXIMM_102_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_102_ARADDR,
    output wire [7:0]                      M_AXIMM_102_ARLEN,
    output wire [2:0]                      M_AXIMM_102_ARSIZE,
    output wire [1:0]                      M_AXIMM_102_ARBURST,
    output wire [1:0]                      M_AXIMM_102_ARLOCK,
    output wire [3:0]                      M_AXIMM_102_ARCACHE,
    output wire [2:0]                      M_AXIMM_102_ARPROT,
    output wire [3:0]                      M_AXIMM_102_ARREGION,
    output wire [3:0]                      M_AXIMM_102_ARQOS,
    output wire                            M_AXIMM_102_ARVALID,
    input  wire                            M_AXIMM_102_ARREADY,
    input  wire [M_AXIMM_102_DATA_WIDTH-1:0]   M_AXIMM_102_RDATA,
    input  wire [1:0]                      M_AXIMM_102_RRESP,
    input  wire                            M_AXIMM_102_RLAST,
    input  wire                            M_AXIMM_102_RVALID,
    output wire                            M_AXIMM_102_RREADY,
    //AXI-MM pass-through interface 103
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_103_AWADDR,
    input wire [7:0]                      AP_AXIMM_103_AWLEN,
    input wire [2:0]                      AP_AXIMM_103_AWSIZE,
    input wire [1:0]                      AP_AXIMM_103_AWBURST,
    input wire [1:0]                      AP_AXIMM_103_AWLOCK,
    input wire [3:0]                      AP_AXIMM_103_AWCACHE,
    input wire [2:0]                      AP_AXIMM_103_AWPROT,
    input wire [3:0]                      AP_AXIMM_103_AWREGION,
    input wire [3:0]                      AP_AXIMM_103_AWQOS,
    input wire                            AP_AXIMM_103_AWVALID,
    output  wire                            AP_AXIMM_103_AWREADY,
    input wire [M_AXIMM_103_DATA_WIDTH-1:0]   AP_AXIMM_103_WDATA,
    input wire [M_AXIMM_103_DATA_WIDTH/8-1:0] AP_AXIMM_103_WSTRB,
    input wire                            AP_AXIMM_103_WLAST,
    input wire                            AP_AXIMM_103_WVALID,
    output  wire                            AP_AXIMM_103_WREADY,
    output  wire [1:0]                      AP_AXIMM_103_BRESP,
    output  wire                            AP_AXIMM_103_BVALID,
    input wire                            AP_AXIMM_103_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_103_ARADDR,
    input wire [7:0]                      AP_AXIMM_103_ARLEN,
    input wire [2:0]                      AP_AXIMM_103_ARSIZE,
    input wire [1:0]                      AP_AXIMM_103_ARBURST,
    input wire [1:0]                      AP_AXIMM_103_ARLOCK,
    input wire [3:0]                      AP_AXIMM_103_ARCACHE,
    input wire [2:0]                      AP_AXIMM_103_ARPROT,
    input wire [3:0]                      AP_AXIMM_103_ARREGION,
    input wire [3:0]                      AP_AXIMM_103_ARQOS,
    input wire                            AP_AXIMM_103_ARVALID,
    output  wire                            AP_AXIMM_103_ARREADY,
    output  wire [M_AXIMM_103_DATA_WIDTH-1:0]   AP_AXIMM_103_RDATA,
    output  wire [1:0]                      AP_AXIMM_103_RRESP,
    output  wire                            AP_AXIMM_103_RLAST,
    output  wire                            AP_AXIMM_103_RVALID,
    input  wire                            AP_AXIMM_103_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_103_AWADDR,
    output wire [7:0]                      M_AXIMM_103_AWLEN,
    output wire [2:0]                      M_AXIMM_103_AWSIZE,
    output wire [1:0]                      M_AXIMM_103_AWBURST,
    output wire [1:0]                      M_AXIMM_103_AWLOCK,
    output wire [3:0]                      M_AXIMM_103_AWCACHE,
    output wire [2:0]                      M_AXIMM_103_AWPROT,
    output wire [3:0]                      M_AXIMM_103_AWREGION,
    output wire [3:0]                      M_AXIMM_103_AWQOS,
    output wire                            M_AXIMM_103_AWVALID,
    input  wire                            M_AXIMM_103_AWREADY,
    output wire [M_AXIMM_103_DATA_WIDTH-1:0]   M_AXIMM_103_WDATA,
    output wire [M_AXIMM_103_DATA_WIDTH/8-1:0] M_AXIMM_103_WSTRB,
    output wire                            M_AXIMM_103_WLAST,
    output wire                            M_AXIMM_103_WVALID,
    input  wire                            M_AXIMM_103_WREADY,
    input  wire [1:0]                      M_AXIMM_103_BRESP,
    input  wire                            M_AXIMM_103_BVALID,
    output wire                            M_AXIMM_103_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_103_ARADDR,
    output wire [7:0]                      M_AXIMM_103_ARLEN,
    output wire [2:0]                      M_AXIMM_103_ARSIZE,
    output wire [1:0]                      M_AXIMM_103_ARBURST,
    output wire [1:0]                      M_AXIMM_103_ARLOCK,
    output wire [3:0]                      M_AXIMM_103_ARCACHE,
    output wire [2:0]                      M_AXIMM_103_ARPROT,
    output wire [3:0]                      M_AXIMM_103_ARREGION,
    output wire [3:0]                      M_AXIMM_103_ARQOS,
    output wire                            M_AXIMM_103_ARVALID,
    input  wire                            M_AXIMM_103_ARREADY,
    input  wire [M_AXIMM_103_DATA_WIDTH-1:0]   M_AXIMM_103_RDATA,
    input  wire [1:0]                      M_AXIMM_103_RRESP,
    input  wire                            M_AXIMM_103_RLAST,
    input  wire                            M_AXIMM_103_RVALID,
    output wire                            M_AXIMM_103_RREADY,
    //AXI-MM pass-through interface 104
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_104_AWADDR,
    input wire [7:0]                      AP_AXIMM_104_AWLEN,
    input wire [2:0]                      AP_AXIMM_104_AWSIZE,
    input wire [1:0]                      AP_AXIMM_104_AWBURST,
    input wire [1:0]                      AP_AXIMM_104_AWLOCK,
    input wire [3:0]                      AP_AXIMM_104_AWCACHE,
    input wire [2:0]                      AP_AXIMM_104_AWPROT,
    input wire [3:0]                      AP_AXIMM_104_AWREGION,
    input wire [3:0]                      AP_AXIMM_104_AWQOS,
    input wire                            AP_AXIMM_104_AWVALID,
    output  wire                            AP_AXIMM_104_AWREADY,
    input wire [M_AXIMM_104_DATA_WIDTH-1:0]   AP_AXIMM_104_WDATA,
    input wire [M_AXIMM_104_DATA_WIDTH/8-1:0] AP_AXIMM_104_WSTRB,
    input wire                            AP_AXIMM_104_WLAST,
    input wire                            AP_AXIMM_104_WVALID,
    output  wire                            AP_AXIMM_104_WREADY,
    output  wire [1:0]                      AP_AXIMM_104_BRESP,
    output  wire                            AP_AXIMM_104_BVALID,
    input wire                            AP_AXIMM_104_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_104_ARADDR,
    input wire [7:0]                      AP_AXIMM_104_ARLEN,
    input wire [2:0]                      AP_AXIMM_104_ARSIZE,
    input wire [1:0]                      AP_AXIMM_104_ARBURST,
    input wire [1:0]                      AP_AXIMM_104_ARLOCK,
    input wire [3:0]                      AP_AXIMM_104_ARCACHE,
    input wire [2:0]                      AP_AXIMM_104_ARPROT,
    input wire [3:0]                      AP_AXIMM_104_ARREGION,
    input wire [3:0]                      AP_AXIMM_104_ARQOS,
    input wire                            AP_AXIMM_104_ARVALID,
    output  wire                            AP_AXIMM_104_ARREADY,
    output  wire [M_AXIMM_104_DATA_WIDTH-1:0]   AP_AXIMM_104_RDATA,
    output  wire [1:0]                      AP_AXIMM_104_RRESP,
    output  wire                            AP_AXIMM_104_RLAST,
    output  wire                            AP_AXIMM_104_RVALID,
    input  wire                            AP_AXIMM_104_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_104_AWADDR,
    output wire [7:0]                      M_AXIMM_104_AWLEN,
    output wire [2:0]                      M_AXIMM_104_AWSIZE,
    output wire [1:0]                      M_AXIMM_104_AWBURST,
    output wire [1:0]                      M_AXIMM_104_AWLOCK,
    output wire [3:0]                      M_AXIMM_104_AWCACHE,
    output wire [2:0]                      M_AXIMM_104_AWPROT,
    output wire [3:0]                      M_AXIMM_104_AWREGION,
    output wire [3:0]                      M_AXIMM_104_AWQOS,
    output wire                            M_AXIMM_104_AWVALID,
    input  wire                            M_AXIMM_104_AWREADY,
    output wire [M_AXIMM_104_DATA_WIDTH-1:0]   M_AXIMM_104_WDATA,
    output wire [M_AXIMM_104_DATA_WIDTH/8-1:0] M_AXIMM_104_WSTRB,
    output wire                            M_AXIMM_104_WLAST,
    output wire                            M_AXIMM_104_WVALID,
    input  wire                            M_AXIMM_104_WREADY,
    input  wire [1:0]                      M_AXIMM_104_BRESP,
    input  wire                            M_AXIMM_104_BVALID,
    output wire                            M_AXIMM_104_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_104_ARADDR,
    output wire [7:0]                      M_AXIMM_104_ARLEN,
    output wire [2:0]                      M_AXIMM_104_ARSIZE,
    output wire [1:0]                      M_AXIMM_104_ARBURST,
    output wire [1:0]                      M_AXIMM_104_ARLOCK,
    output wire [3:0]                      M_AXIMM_104_ARCACHE,
    output wire [2:0]                      M_AXIMM_104_ARPROT,
    output wire [3:0]                      M_AXIMM_104_ARREGION,
    output wire [3:0]                      M_AXIMM_104_ARQOS,
    output wire                            M_AXIMM_104_ARVALID,
    input  wire                            M_AXIMM_104_ARREADY,
    input  wire [M_AXIMM_104_DATA_WIDTH-1:0]   M_AXIMM_104_RDATA,
    input  wire [1:0]                      M_AXIMM_104_RRESP,
    input  wire                            M_AXIMM_104_RLAST,
    input  wire                            M_AXIMM_104_RVALID,
    output wire                            M_AXIMM_104_RREADY,
    //AXI-MM pass-through interface 105
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_105_AWADDR,
    input wire [7:0]                      AP_AXIMM_105_AWLEN,
    input wire [2:0]                      AP_AXIMM_105_AWSIZE,
    input wire [1:0]                      AP_AXIMM_105_AWBURST,
    input wire [1:0]                      AP_AXIMM_105_AWLOCK,
    input wire [3:0]                      AP_AXIMM_105_AWCACHE,
    input wire [2:0]                      AP_AXIMM_105_AWPROT,
    input wire [3:0]                      AP_AXIMM_105_AWREGION,
    input wire [3:0]                      AP_AXIMM_105_AWQOS,
    input wire                            AP_AXIMM_105_AWVALID,
    output  wire                            AP_AXIMM_105_AWREADY,
    input wire [M_AXIMM_105_DATA_WIDTH-1:0]   AP_AXIMM_105_WDATA,
    input wire [M_AXIMM_105_DATA_WIDTH/8-1:0] AP_AXIMM_105_WSTRB,
    input wire                            AP_AXIMM_105_WLAST,
    input wire                            AP_AXIMM_105_WVALID,
    output  wire                            AP_AXIMM_105_WREADY,
    output  wire [1:0]                      AP_AXIMM_105_BRESP,
    output  wire                            AP_AXIMM_105_BVALID,
    input wire                            AP_AXIMM_105_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_105_ARADDR,
    input wire [7:0]                      AP_AXIMM_105_ARLEN,
    input wire [2:0]                      AP_AXIMM_105_ARSIZE,
    input wire [1:0]                      AP_AXIMM_105_ARBURST,
    input wire [1:0]                      AP_AXIMM_105_ARLOCK,
    input wire [3:0]                      AP_AXIMM_105_ARCACHE,
    input wire [2:0]                      AP_AXIMM_105_ARPROT,
    input wire [3:0]                      AP_AXIMM_105_ARREGION,
    input wire [3:0]                      AP_AXIMM_105_ARQOS,
    input wire                            AP_AXIMM_105_ARVALID,
    output  wire                            AP_AXIMM_105_ARREADY,
    output  wire [M_AXIMM_105_DATA_WIDTH-1:0]   AP_AXIMM_105_RDATA,
    output  wire [1:0]                      AP_AXIMM_105_RRESP,
    output  wire                            AP_AXIMM_105_RLAST,
    output  wire                            AP_AXIMM_105_RVALID,
    input  wire                            AP_AXIMM_105_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_105_AWADDR,
    output wire [7:0]                      M_AXIMM_105_AWLEN,
    output wire [2:0]                      M_AXIMM_105_AWSIZE,
    output wire [1:0]                      M_AXIMM_105_AWBURST,
    output wire [1:0]                      M_AXIMM_105_AWLOCK,
    output wire [3:0]                      M_AXIMM_105_AWCACHE,
    output wire [2:0]                      M_AXIMM_105_AWPROT,
    output wire [3:0]                      M_AXIMM_105_AWREGION,
    output wire [3:0]                      M_AXIMM_105_AWQOS,
    output wire                            M_AXIMM_105_AWVALID,
    input  wire                            M_AXIMM_105_AWREADY,
    output wire [M_AXIMM_105_DATA_WIDTH-1:0]   M_AXIMM_105_WDATA,
    output wire [M_AXIMM_105_DATA_WIDTH/8-1:0] M_AXIMM_105_WSTRB,
    output wire                            M_AXIMM_105_WLAST,
    output wire                            M_AXIMM_105_WVALID,
    input  wire                            M_AXIMM_105_WREADY,
    input  wire [1:0]                      M_AXIMM_105_BRESP,
    input  wire                            M_AXIMM_105_BVALID,
    output wire                            M_AXIMM_105_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_105_ARADDR,
    output wire [7:0]                      M_AXIMM_105_ARLEN,
    output wire [2:0]                      M_AXIMM_105_ARSIZE,
    output wire [1:0]                      M_AXIMM_105_ARBURST,
    output wire [1:0]                      M_AXIMM_105_ARLOCK,
    output wire [3:0]                      M_AXIMM_105_ARCACHE,
    output wire [2:0]                      M_AXIMM_105_ARPROT,
    output wire [3:0]                      M_AXIMM_105_ARREGION,
    output wire [3:0]                      M_AXIMM_105_ARQOS,
    output wire                            M_AXIMM_105_ARVALID,
    input  wire                            M_AXIMM_105_ARREADY,
    input  wire [M_AXIMM_105_DATA_WIDTH-1:0]   M_AXIMM_105_RDATA,
    input  wire [1:0]                      M_AXIMM_105_RRESP,
    input  wire                            M_AXIMM_105_RLAST,
    input  wire                            M_AXIMM_105_RVALID,
    output wire                            M_AXIMM_105_RREADY,
    //AXI-MM pass-through interface 106
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_106_AWADDR,
    input wire [7:0]                      AP_AXIMM_106_AWLEN,
    input wire [2:0]                      AP_AXIMM_106_AWSIZE,
    input wire [1:0]                      AP_AXIMM_106_AWBURST,
    input wire [1:0]                      AP_AXIMM_106_AWLOCK,
    input wire [3:0]                      AP_AXIMM_106_AWCACHE,
    input wire [2:0]                      AP_AXIMM_106_AWPROT,
    input wire [3:0]                      AP_AXIMM_106_AWREGION,
    input wire [3:0]                      AP_AXIMM_106_AWQOS,
    input wire                            AP_AXIMM_106_AWVALID,
    output  wire                            AP_AXIMM_106_AWREADY,
    input wire [M_AXIMM_106_DATA_WIDTH-1:0]   AP_AXIMM_106_WDATA,
    input wire [M_AXIMM_106_DATA_WIDTH/8-1:0] AP_AXIMM_106_WSTRB,
    input wire                            AP_AXIMM_106_WLAST,
    input wire                            AP_AXIMM_106_WVALID,
    output  wire                            AP_AXIMM_106_WREADY,
    output  wire [1:0]                      AP_AXIMM_106_BRESP,
    output  wire                            AP_AXIMM_106_BVALID,
    input wire                            AP_AXIMM_106_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_106_ARADDR,
    input wire [7:0]                      AP_AXIMM_106_ARLEN,
    input wire [2:0]                      AP_AXIMM_106_ARSIZE,
    input wire [1:0]                      AP_AXIMM_106_ARBURST,
    input wire [1:0]                      AP_AXIMM_106_ARLOCK,
    input wire [3:0]                      AP_AXIMM_106_ARCACHE,
    input wire [2:0]                      AP_AXIMM_106_ARPROT,
    input wire [3:0]                      AP_AXIMM_106_ARREGION,
    input wire [3:0]                      AP_AXIMM_106_ARQOS,
    input wire                            AP_AXIMM_106_ARVALID,
    output  wire                            AP_AXIMM_106_ARREADY,
    output  wire [M_AXIMM_106_DATA_WIDTH-1:0]   AP_AXIMM_106_RDATA,
    output  wire [1:0]                      AP_AXIMM_106_RRESP,
    output  wire                            AP_AXIMM_106_RLAST,
    output  wire                            AP_AXIMM_106_RVALID,
    input  wire                            AP_AXIMM_106_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_106_AWADDR,
    output wire [7:0]                      M_AXIMM_106_AWLEN,
    output wire [2:0]                      M_AXIMM_106_AWSIZE,
    output wire [1:0]                      M_AXIMM_106_AWBURST,
    output wire [1:0]                      M_AXIMM_106_AWLOCK,
    output wire [3:0]                      M_AXIMM_106_AWCACHE,
    output wire [2:0]                      M_AXIMM_106_AWPROT,
    output wire [3:0]                      M_AXIMM_106_AWREGION,
    output wire [3:0]                      M_AXIMM_106_AWQOS,
    output wire                            M_AXIMM_106_AWVALID,
    input  wire                            M_AXIMM_106_AWREADY,
    output wire [M_AXIMM_106_DATA_WIDTH-1:0]   M_AXIMM_106_WDATA,
    output wire [M_AXIMM_106_DATA_WIDTH/8-1:0] M_AXIMM_106_WSTRB,
    output wire                            M_AXIMM_106_WLAST,
    output wire                            M_AXIMM_106_WVALID,
    input  wire                            M_AXIMM_106_WREADY,
    input  wire [1:0]                      M_AXIMM_106_BRESP,
    input  wire                            M_AXIMM_106_BVALID,
    output wire                            M_AXIMM_106_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_106_ARADDR,
    output wire [7:0]                      M_AXIMM_106_ARLEN,
    output wire [2:0]                      M_AXIMM_106_ARSIZE,
    output wire [1:0]                      M_AXIMM_106_ARBURST,
    output wire [1:0]                      M_AXIMM_106_ARLOCK,
    output wire [3:0]                      M_AXIMM_106_ARCACHE,
    output wire [2:0]                      M_AXIMM_106_ARPROT,
    output wire [3:0]                      M_AXIMM_106_ARREGION,
    output wire [3:0]                      M_AXIMM_106_ARQOS,
    output wire                            M_AXIMM_106_ARVALID,
    input  wire                            M_AXIMM_106_ARREADY,
    input  wire [M_AXIMM_106_DATA_WIDTH-1:0]   M_AXIMM_106_RDATA,
    input  wire [1:0]                      M_AXIMM_106_RRESP,
    input  wire                            M_AXIMM_106_RLAST,
    input  wire                            M_AXIMM_106_RVALID,
    output wire                            M_AXIMM_106_RREADY,
    //AXI-MM pass-through interface 107
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_107_AWADDR,
    input wire [7:0]                      AP_AXIMM_107_AWLEN,
    input wire [2:0]                      AP_AXIMM_107_AWSIZE,
    input wire [1:0]                      AP_AXIMM_107_AWBURST,
    input wire [1:0]                      AP_AXIMM_107_AWLOCK,
    input wire [3:0]                      AP_AXIMM_107_AWCACHE,
    input wire [2:0]                      AP_AXIMM_107_AWPROT,
    input wire [3:0]                      AP_AXIMM_107_AWREGION,
    input wire [3:0]                      AP_AXIMM_107_AWQOS,
    input wire                            AP_AXIMM_107_AWVALID,
    output  wire                            AP_AXIMM_107_AWREADY,
    input wire [M_AXIMM_107_DATA_WIDTH-1:0]   AP_AXIMM_107_WDATA,
    input wire [M_AXIMM_107_DATA_WIDTH/8-1:0] AP_AXIMM_107_WSTRB,
    input wire                            AP_AXIMM_107_WLAST,
    input wire                            AP_AXIMM_107_WVALID,
    output  wire                            AP_AXIMM_107_WREADY,
    output  wire [1:0]                      AP_AXIMM_107_BRESP,
    output  wire                            AP_AXIMM_107_BVALID,
    input wire                            AP_AXIMM_107_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_107_ARADDR,
    input wire [7:0]                      AP_AXIMM_107_ARLEN,
    input wire [2:0]                      AP_AXIMM_107_ARSIZE,
    input wire [1:0]                      AP_AXIMM_107_ARBURST,
    input wire [1:0]                      AP_AXIMM_107_ARLOCK,
    input wire [3:0]                      AP_AXIMM_107_ARCACHE,
    input wire [2:0]                      AP_AXIMM_107_ARPROT,
    input wire [3:0]                      AP_AXIMM_107_ARREGION,
    input wire [3:0]                      AP_AXIMM_107_ARQOS,
    input wire                            AP_AXIMM_107_ARVALID,
    output  wire                            AP_AXIMM_107_ARREADY,
    output  wire [M_AXIMM_107_DATA_WIDTH-1:0]   AP_AXIMM_107_RDATA,
    output  wire [1:0]                      AP_AXIMM_107_RRESP,
    output  wire                            AP_AXIMM_107_RLAST,
    output  wire                            AP_AXIMM_107_RVALID,
    input  wire                            AP_AXIMM_107_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_107_AWADDR,
    output wire [7:0]                      M_AXIMM_107_AWLEN,
    output wire [2:0]                      M_AXIMM_107_AWSIZE,
    output wire [1:0]                      M_AXIMM_107_AWBURST,
    output wire [1:0]                      M_AXIMM_107_AWLOCK,
    output wire [3:0]                      M_AXIMM_107_AWCACHE,
    output wire [2:0]                      M_AXIMM_107_AWPROT,
    output wire [3:0]                      M_AXIMM_107_AWREGION,
    output wire [3:0]                      M_AXIMM_107_AWQOS,
    output wire                            M_AXIMM_107_AWVALID,
    input  wire                            M_AXIMM_107_AWREADY,
    output wire [M_AXIMM_107_DATA_WIDTH-1:0]   M_AXIMM_107_WDATA,
    output wire [M_AXIMM_107_DATA_WIDTH/8-1:0] M_AXIMM_107_WSTRB,
    output wire                            M_AXIMM_107_WLAST,
    output wire                            M_AXIMM_107_WVALID,
    input  wire                            M_AXIMM_107_WREADY,
    input  wire [1:0]                      M_AXIMM_107_BRESP,
    input  wire                            M_AXIMM_107_BVALID,
    output wire                            M_AXIMM_107_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_107_ARADDR,
    output wire [7:0]                      M_AXIMM_107_ARLEN,
    output wire [2:0]                      M_AXIMM_107_ARSIZE,
    output wire [1:0]                      M_AXIMM_107_ARBURST,
    output wire [1:0]                      M_AXIMM_107_ARLOCK,
    output wire [3:0]                      M_AXIMM_107_ARCACHE,
    output wire [2:0]                      M_AXIMM_107_ARPROT,
    output wire [3:0]                      M_AXIMM_107_ARREGION,
    output wire [3:0]                      M_AXIMM_107_ARQOS,
    output wire                            M_AXIMM_107_ARVALID,
    input  wire                            M_AXIMM_107_ARREADY,
    input  wire [M_AXIMM_107_DATA_WIDTH-1:0]   M_AXIMM_107_RDATA,
    input  wire [1:0]                      M_AXIMM_107_RRESP,
    input  wire                            M_AXIMM_107_RLAST,
    input  wire                            M_AXIMM_107_RVALID,
    output wire                            M_AXIMM_107_RREADY,
    //AXI-MM pass-through interface 108
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_108_AWADDR,
    input wire [7:0]                      AP_AXIMM_108_AWLEN,
    input wire [2:0]                      AP_AXIMM_108_AWSIZE,
    input wire [1:0]                      AP_AXIMM_108_AWBURST,
    input wire [1:0]                      AP_AXIMM_108_AWLOCK,
    input wire [3:0]                      AP_AXIMM_108_AWCACHE,
    input wire [2:0]                      AP_AXIMM_108_AWPROT,
    input wire [3:0]                      AP_AXIMM_108_AWREGION,
    input wire [3:0]                      AP_AXIMM_108_AWQOS,
    input wire                            AP_AXIMM_108_AWVALID,
    output  wire                            AP_AXIMM_108_AWREADY,
    input wire [M_AXIMM_108_DATA_WIDTH-1:0]   AP_AXIMM_108_WDATA,
    input wire [M_AXIMM_108_DATA_WIDTH/8-1:0] AP_AXIMM_108_WSTRB,
    input wire                            AP_AXIMM_108_WLAST,
    input wire                            AP_AXIMM_108_WVALID,
    output  wire                            AP_AXIMM_108_WREADY,
    output  wire [1:0]                      AP_AXIMM_108_BRESP,
    output  wire                            AP_AXIMM_108_BVALID,
    input wire                            AP_AXIMM_108_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_108_ARADDR,
    input wire [7:0]                      AP_AXIMM_108_ARLEN,
    input wire [2:0]                      AP_AXIMM_108_ARSIZE,
    input wire [1:0]                      AP_AXIMM_108_ARBURST,
    input wire [1:0]                      AP_AXIMM_108_ARLOCK,
    input wire [3:0]                      AP_AXIMM_108_ARCACHE,
    input wire [2:0]                      AP_AXIMM_108_ARPROT,
    input wire [3:0]                      AP_AXIMM_108_ARREGION,
    input wire [3:0]                      AP_AXIMM_108_ARQOS,
    input wire                            AP_AXIMM_108_ARVALID,
    output  wire                            AP_AXIMM_108_ARREADY,
    output  wire [M_AXIMM_108_DATA_WIDTH-1:0]   AP_AXIMM_108_RDATA,
    output  wire [1:0]                      AP_AXIMM_108_RRESP,
    output  wire                            AP_AXIMM_108_RLAST,
    output  wire                            AP_AXIMM_108_RVALID,
    input  wire                            AP_AXIMM_108_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_108_AWADDR,
    output wire [7:0]                      M_AXIMM_108_AWLEN,
    output wire [2:0]                      M_AXIMM_108_AWSIZE,
    output wire [1:0]                      M_AXIMM_108_AWBURST,
    output wire [1:0]                      M_AXIMM_108_AWLOCK,
    output wire [3:0]                      M_AXIMM_108_AWCACHE,
    output wire [2:0]                      M_AXIMM_108_AWPROT,
    output wire [3:0]                      M_AXIMM_108_AWREGION,
    output wire [3:0]                      M_AXIMM_108_AWQOS,
    output wire                            M_AXIMM_108_AWVALID,
    input  wire                            M_AXIMM_108_AWREADY,
    output wire [M_AXIMM_108_DATA_WIDTH-1:0]   M_AXIMM_108_WDATA,
    output wire [M_AXIMM_108_DATA_WIDTH/8-1:0] M_AXIMM_108_WSTRB,
    output wire                            M_AXIMM_108_WLAST,
    output wire                            M_AXIMM_108_WVALID,
    input  wire                            M_AXIMM_108_WREADY,
    input  wire [1:0]                      M_AXIMM_108_BRESP,
    input  wire                            M_AXIMM_108_BVALID,
    output wire                            M_AXIMM_108_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_108_ARADDR,
    output wire [7:0]                      M_AXIMM_108_ARLEN,
    output wire [2:0]                      M_AXIMM_108_ARSIZE,
    output wire [1:0]                      M_AXIMM_108_ARBURST,
    output wire [1:0]                      M_AXIMM_108_ARLOCK,
    output wire [3:0]                      M_AXIMM_108_ARCACHE,
    output wire [2:0]                      M_AXIMM_108_ARPROT,
    output wire [3:0]                      M_AXIMM_108_ARREGION,
    output wire [3:0]                      M_AXIMM_108_ARQOS,
    output wire                            M_AXIMM_108_ARVALID,
    input  wire                            M_AXIMM_108_ARREADY,
    input  wire [M_AXIMM_108_DATA_WIDTH-1:0]   M_AXIMM_108_RDATA,
    input  wire [1:0]                      M_AXIMM_108_RRESP,
    input  wire                            M_AXIMM_108_RLAST,
    input  wire                            M_AXIMM_108_RVALID,
    output wire                            M_AXIMM_108_RREADY,
    //AXI-MM pass-through interface 109
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_109_AWADDR,
    input wire [7:0]                      AP_AXIMM_109_AWLEN,
    input wire [2:0]                      AP_AXIMM_109_AWSIZE,
    input wire [1:0]                      AP_AXIMM_109_AWBURST,
    input wire [1:0]                      AP_AXIMM_109_AWLOCK,
    input wire [3:0]                      AP_AXIMM_109_AWCACHE,
    input wire [2:0]                      AP_AXIMM_109_AWPROT,
    input wire [3:0]                      AP_AXIMM_109_AWREGION,
    input wire [3:0]                      AP_AXIMM_109_AWQOS,
    input wire                            AP_AXIMM_109_AWVALID,
    output  wire                            AP_AXIMM_109_AWREADY,
    input wire [M_AXIMM_109_DATA_WIDTH-1:0]   AP_AXIMM_109_WDATA,
    input wire [M_AXIMM_109_DATA_WIDTH/8-1:0] AP_AXIMM_109_WSTRB,
    input wire                            AP_AXIMM_109_WLAST,
    input wire                            AP_AXIMM_109_WVALID,
    output  wire                            AP_AXIMM_109_WREADY,
    output  wire [1:0]                      AP_AXIMM_109_BRESP,
    output  wire                            AP_AXIMM_109_BVALID,
    input wire                            AP_AXIMM_109_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_109_ARADDR,
    input wire [7:0]                      AP_AXIMM_109_ARLEN,
    input wire [2:0]                      AP_AXIMM_109_ARSIZE,
    input wire [1:0]                      AP_AXIMM_109_ARBURST,
    input wire [1:0]                      AP_AXIMM_109_ARLOCK,
    input wire [3:0]                      AP_AXIMM_109_ARCACHE,
    input wire [2:0]                      AP_AXIMM_109_ARPROT,
    input wire [3:0]                      AP_AXIMM_109_ARREGION,
    input wire [3:0]                      AP_AXIMM_109_ARQOS,
    input wire                            AP_AXIMM_109_ARVALID,
    output  wire                            AP_AXIMM_109_ARREADY,
    output  wire [M_AXIMM_109_DATA_WIDTH-1:0]   AP_AXIMM_109_RDATA,
    output  wire [1:0]                      AP_AXIMM_109_RRESP,
    output  wire                            AP_AXIMM_109_RLAST,
    output  wire                            AP_AXIMM_109_RVALID,
    input  wire                            AP_AXIMM_109_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_109_AWADDR,
    output wire [7:0]                      M_AXIMM_109_AWLEN,
    output wire [2:0]                      M_AXIMM_109_AWSIZE,
    output wire [1:0]                      M_AXIMM_109_AWBURST,
    output wire [1:0]                      M_AXIMM_109_AWLOCK,
    output wire [3:0]                      M_AXIMM_109_AWCACHE,
    output wire [2:0]                      M_AXIMM_109_AWPROT,
    output wire [3:0]                      M_AXIMM_109_AWREGION,
    output wire [3:0]                      M_AXIMM_109_AWQOS,
    output wire                            M_AXIMM_109_AWVALID,
    input  wire                            M_AXIMM_109_AWREADY,
    output wire [M_AXIMM_109_DATA_WIDTH-1:0]   M_AXIMM_109_WDATA,
    output wire [M_AXIMM_109_DATA_WIDTH/8-1:0] M_AXIMM_109_WSTRB,
    output wire                            M_AXIMM_109_WLAST,
    output wire                            M_AXIMM_109_WVALID,
    input  wire                            M_AXIMM_109_WREADY,
    input  wire [1:0]                      M_AXIMM_109_BRESP,
    input  wire                            M_AXIMM_109_BVALID,
    output wire                            M_AXIMM_109_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_109_ARADDR,
    output wire [7:0]                      M_AXIMM_109_ARLEN,
    output wire [2:0]                      M_AXIMM_109_ARSIZE,
    output wire [1:0]                      M_AXIMM_109_ARBURST,
    output wire [1:0]                      M_AXIMM_109_ARLOCK,
    output wire [3:0]                      M_AXIMM_109_ARCACHE,
    output wire [2:0]                      M_AXIMM_109_ARPROT,
    output wire [3:0]                      M_AXIMM_109_ARREGION,
    output wire [3:0]                      M_AXIMM_109_ARQOS,
    output wire                            M_AXIMM_109_ARVALID,
    input  wire                            M_AXIMM_109_ARREADY,
    input  wire [M_AXIMM_109_DATA_WIDTH-1:0]   M_AXIMM_109_RDATA,
    input  wire [1:0]                      M_AXIMM_109_RRESP,
    input  wire                            M_AXIMM_109_RLAST,
    input  wire                            M_AXIMM_109_RVALID,
    output wire                            M_AXIMM_109_RREADY,
    //AXI-MM pass-through interface 110
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_110_AWADDR,
    input wire [7:0]                      AP_AXIMM_110_AWLEN,
    input wire [2:0]                      AP_AXIMM_110_AWSIZE,
    input wire [1:0]                      AP_AXIMM_110_AWBURST,
    input wire [1:0]                      AP_AXIMM_110_AWLOCK,
    input wire [3:0]                      AP_AXIMM_110_AWCACHE,
    input wire [2:0]                      AP_AXIMM_110_AWPROT,
    input wire [3:0]                      AP_AXIMM_110_AWREGION,
    input wire [3:0]                      AP_AXIMM_110_AWQOS,
    input wire                            AP_AXIMM_110_AWVALID,
    output  wire                            AP_AXIMM_110_AWREADY,
    input wire [M_AXIMM_110_DATA_WIDTH-1:0]   AP_AXIMM_110_WDATA,
    input wire [M_AXIMM_110_DATA_WIDTH/8-1:0] AP_AXIMM_110_WSTRB,
    input wire                            AP_AXIMM_110_WLAST,
    input wire                            AP_AXIMM_110_WVALID,
    output  wire                            AP_AXIMM_110_WREADY,
    output  wire [1:0]                      AP_AXIMM_110_BRESP,
    output  wire                            AP_AXIMM_110_BVALID,
    input wire                            AP_AXIMM_110_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_110_ARADDR,
    input wire [7:0]                      AP_AXIMM_110_ARLEN,
    input wire [2:0]                      AP_AXIMM_110_ARSIZE,
    input wire [1:0]                      AP_AXIMM_110_ARBURST,
    input wire [1:0]                      AP_AXIMM_110_ARLOCK,
    input wire [3:0]                      AP_AXIMM_110_ARCACHE,
    input wire [2:0]                      AP_AXIMM_110_ARPROT,
    input wire [3:0]                      AP_AXIMM_110_ARREGION,
    input wire [3:0]                      AP_AXIMM_110_ARQOS,
    input wire                            AP_AXIMM_110_ARVALID,
    output  wire                            AP_AXIMM_110_ARREADY,
    output  wire [M_AXIMM_110_DATA_WIDTH-1:0]   AP_AXIMM_110_RDATA,
    output  wire [1:0]                      AP_AXIMM_110_RRESP,
    output  wire                            AP_AXIMM_110_RLAST,
    output  wire                            AP_AXIMM_110_RVALID,
    input  wire                            AP_AXIMM_110_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_110_AWADDR,
    output wire [7:0]                      M_AXIMM_110_AWLEN,
    output wire [2:0]                      M_AXIMM_110_AWSIZE,
    output wire [1:0]                      M_AXIMM_110_AWBURST,
    output wire [1:0]                      M_AXIMM_110_AWLOCK,
    output wire [3:0]                      M_AXIMM_110_AWCACHE,
    output wire [2:0]                      M_AXIMM_110_AWPROT,
    output wire [3:0]                      M_AXIMM_110_AWREGION,
    output wire [3:0]                      M_AXIMM_110_AWQOS,
    output wire                            M_AXIMM_110_AWVALID,
    input  wire                            M_AXIMM_110_AWREADY,
    output wire [M_AXIMM_110_DATA_WIDTH-1:0]   M_AXIMM_110_WDATA,
    output wire [M_AXIMM_110_DATA_WIDTH/8-1:0] M_AXIMM_110_WSTRB,
    output wire                            M_AXIMM_110_WLAST,
    output wire                            M_AXIMM_110_WVALID,
    input  wire                            M_AXIMM_110_WREADY,
    input  wire [1:0]                      M_AXIMM_110_BRESP,
    input  wire                            M_AXIMM_110_BVALID,
    output wire                            M_AXIMM_110_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_110_ARADDR,
    output wire [7:0]                      M_AXIMM_110_ARLEN,
    output wire [2:0]                      M_AXIMM_110_ARSIZE,
    output wire [1:0]                      M_AXIMM_110_ARBURST,
    output wire [1:0]                      M_AXIMM_110_ARLOCK,
    output wire [3:0]                      M_AXIMM_110_ARCACHE,
    output wire [2:0]                      M_AXIMM_110_ARPROT,
    output wire [3:0]                      M_AXIMM_110_ARREGION,
    output wire [3:0]                      M_AXIMM_110_ARQOS,
    output wire                            M_AXIMM_110_ARVALID,
    input  wire                            M_AXIMM_110_ARREADY,
    input  wire [M_AXIMM_110_DATA_WIDTH-1:0]   M_AXIMM_110_RDATA,
    input  wire [1:0]                      M_AXIMM_110_RRESP,
    input  wire                            M_AXIMM_110_RLAST,
    input  wire                            M_AXIMM_110_RVALID,
    output wire                            M_AXIMM_110_RREADY,
    //AXI-MM pass-through interface 111
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_111_AWADDR,
    input wire [7:0]                      AP_AXIMM_111_AWLEN,
    input wire [2:0]                      AP_AXIMM_111_AWSIZE,
    input wire [1:0]                      AP_AXIMM_111_AWBURST,
    input wire [1:0]                      AP_AXIMM_111_AWLOCK,
    input wire [3:0]                      AP_AXIMM_111_AWCACHE,
    input wire [2:0]                      AP_AXIMM_111_AWPROT,
    input wire [3:0]                      AP_AXIMM_111_AWREGION,
    input wire [3:0]                      AP_AXIMM_111_AWQOS,
    input wire                            AP_AXIMM_111_AWVALID,
    output  wire                            AP_AXIMM_111_AWREADY,
    input wire [M_AXIMM_111_DATA_WIDTH-1:0]   AP_AXIMM_111_WDATA,
    input wire [M_AXIMM_111_DATA_WIDTH/8-1:0] AP_AXIMM_111_WSTRB,
    input wire                            AP_AXIMM_111_WLAST,
    input wire                            AP_AXIMM_111_WVALID,
    output  wire                            AP_AXIMM_111_WREADY,
    output  wire [1:0]                      AP_AXIMM_111_BRESP,
    output  wire                            AP_AXIMM_111_BVALID,
    input wire                            AP_AXIMM_111_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_111_ARADDR,
    input wire [7:0]                      AP_AXIMM_111_ARLEN,
    input wire [2:0]                      AP_AXIMM_111_ARSIZE,
    input wire [1:0]                      AP_AXIMM_111_ARBURST,
    input wire [1:0]                      AP_AXIMM_111_ARLOCK,
    input wire [3:0]                      AP_AXIMM_111_ARCACHE,
    input wire [2:0]                      AP_AXIMM_111_ARPROT,
    input wire [3:0]                      AP_AXIMM_111_ARREGION,
    input wire [3:0]                      AP_AXIMM_111_ARQOS,
    input wire                            AP_AXIMM_111_ARVALID,
    output  wire                            AP_AXIMM_111_ARREADY,
    output  wire [M_AXIMM_111_DATA_WIDTH-1:0]   AP_AXIMM_111_RDATA,
    output  wire [1:0]                      AP_AXIMM_111_RRESP,
    output  wire                            AP_AXIMM_111_RLAST,
    output  wire                            AP_AXIMM_111_RVALID,
    input  wire                            AP_AXIMM_111_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_111_AWADDR,
    output wire [7:0]                      M_AXIMM_111_AWLEN,
    output wire [2:0]                      M_AXIMM_111_AWSIZE,
    output wire [1:0]                      M_AXIMM_111_AWBURST,
    output wire [1:0]                      M_AXIMM_111_AWLOCK,
    output wire [3:0]                      M_AXIMM_111_AWCACHE,
    output wire [2:0]                      M_AXIMM_111_AWPROT,
    output wire [3:0]                      M_AXIMM_111_AWREGION,
    output wire [3:0]                      M_AXIMM_111_AWQOS,
    output wire                            M_AXIMM_111_AWVALID,
    input  wire                            M_AXIMM_111_AWREADY,
    output wire [M_AXIMM_111_DATA_WIDTH-1:0]   M_AXIMM_111_WDATA,
    output wire [M_AXIMM_111_DATA_WIDTH/8-1:0] M_AXIMM_111_WSTRB,
    output wire                            M_AXIMM_111_WLAST,
    output wire                            M_AXIMM_111_WVALID,
    input  wire                            M_AXIMM_111_WREADY,
    input  wire [1:0]                      M_AXIMM_111_BRESP,
    input  wire                            M_AXIMM_111_BVALID,
    output wire                            M_AXIMM_111_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_111_ARADDR,
    output wire [7:0]                      M_AXIMM_111_ARLEN,
    output wire [2:0]                      M_AXIMM_111_ARSIZE,
    output wire [1:0]                      M_AXIMM_111_ARBURST,
    output wire [1:0]                      M_AXIMM_111_ARLOCK,
    output wire [3:0]                      M_AXIMM_111_ARCACHE,
    output wire [2:0]                      M_AXIMM_111_ARPROT,
    output wire [3:0]                      M_AXIMM_111_ARREGION,
    output wire [3:0]                      M_AXIMM_111_ARQOS,
    output wire                            M_AXIMM_111_ARVALID,
    input  wire                            M_AXIMM_111_ARREADY,
    input  wire [M_AXIMM_111_DATA_WIDTH-1:0]   M_AXIMM_111_RDATA,
    input  wire [1:0]                      M_AXIMM_111_RRESP,
    input  wire                            M_AXIMM_111_RLAST,
    input  wire                            M_AXIMM_111_RVALID,
    output wire                            M_AXIMM_111_RREADY,
    //AXI-MM pass-through interface 112
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_112_AWADDR,
    input wire [7:0]                      AP_AXIMM_112_AWLEN,
    input wire [2:0]                      AP_AXIMM_112_AWSIZE,
    input wire [1:0]                      AP_AXIMM_112_AWBURST,
    input wire [1:0]                      AP_AXIMM_112_AWLOCK,
    input wire [3:0]                      AP_AXIMM_112_AWCACHE,
    input wire [2:0]                      AP_AXIMM_112_AWPROT,
    input wire [3:0]                      AP_AXIMM_112_AWREGION,
    input wire [3:0]                      AP_AXIMM_112_AWQOS,
    input wire                            AP_AXIMM_112_AWVALID,
    output  wire                            AP_AXIMM_112_AWREADY,
    input wire [M_AXIMM_112_DATA_WIDTH-1:0]   AP_AXIMM_112_WDATA,
    input wire [M_AXIMM_112_DATA_WIDTH/8-1:0] AP_AXIMM_112_WSTRB,
    input wire                            AP_AXIMM_112_WLAST,
    input wire                            AP_AXIMM_112_WVALID,
    output  wire                            AP_AXIMM_112_WREADY,
    output  wire [1:0]                      AP_AXIMM_112_BRESP,
    output  wire                            AP_AXIMM_112_BVALID,
    input wire                            AP_AXIMM_112_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_112_ARADDR,
    input wire [7:0]                      AP_AXIMM_112_ARLEN,
    input wire [2:0]                      AP_AXIMM_112_ARSIZE,
    input wire [1:0]                      AP_AXIMM_112_ARBURST,
    input wire [1:0]                      AP_AXIMM_112_ARLOCK,
    input wire [3:0]                      AP_AXIMM_112_ARCACHE,
    input wire [2:0]                      AP_AXIMM_112_ARPROT,
    input wire [3:0]                      AP_AXIMM_112_ARREGION,
    input wire [3:0]                      AP_AXIMM_112_ARQOS,
    input wire                            AP_AXIMM_112_ARVALID,
    output  wire                            AP_AXIMM_112_ARREADY,
    output  wire [M_AXIMM_112_DATA_WIDTH-1:0]   AP_AXIMM_112_RDATA,
    output  wire [1:0]                      AP_AXIMM_112_RRESP,
    output  wire                            AP_AXIMM_112_RLAST,
    output  wire                            AP_AXIMM_112_RVALID,
    input  wire                            AP_AXIMM_112_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_112_AWADDR,
    output wire [7:0]                      M_AXIMM_112_AWLEN,
    output wire [2:0]                      M_AXIMM_112_AWSIZE,
    output wire [1:0]                      M_AXIMM_112_AWBURST,
    output wire [1:0]                      M_AXIMM_112_AWLOCK,
    output wire [3:0]                      M_AXIMM_112_AWCACHE,
    output wire [2:0]                      M_AXIMM_112_AWPROT,
    output wire [3:0]                      M_AXIMM_112_AWREGION,
    output wire [3:0]                      M_AXIMM_112_AWQOS,
    output wire                            M_AXIMM_112_AWVALID,
    input  wire                            M_AXIMM_112_AWREADY,
    output wire [M_AXIMM_112_DATA_WIDTH-1:0]   M_AXIMM_112_WDATA,
    output wire [M_AXIMM_112_DATA_WIDTH/8-1:0] M_AXIMM_112_WSTRB,
    output wire                            M_AXIMM_112_WLAST,
    output wire                            M_AXIMM_112_WVALID,
    input  wire                            M_AXIMM_112_WREADY,
    input  wire [1:0]                      M_AXIMM_112_BRESP,
    input  wire                            M_AXIMM_112_BVALID,
    output wire                            M_AXIMM_112_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_112_ARADDR,
    output wire [7:0]                      M_AXIMM_112_ARLEN,
    output wire [2:0]                      M_AXIMM_112_ARSIZE,
    output wire [1:0]                      M_AXIMM_112_ARBURST,
    output wire [1:0]                      M_AXIMM_112_ARLOCK,
    output wire [3:0]                      M_AXIMM_112_ARCACHE,
    output wire [2:0]                      M_AXIMM_112_ARPROT,
    output wire [3:0]                      M_AXIMM_112_ARREGION,
    output wire [3:0]                      M_AXIMM_112_ARQOS,
    output wire                            M_AXIMM_112_ARVALID,
    input  wire                            M_AXIMM_112_ARREADY,
    input  wire [M_AXIMM_112_DATA_WIDTH-1:0]   M_AXIMM_112_RDATA,
    input  wire [1:0]                      M_AXIMM_112_RRESP,
    input  wire                            M_AXIMM_112_RLAST,
    input  wire                            M_AXIMM_112_RVALID,
    output wire                            M_AXIMM_112_RREADY,
    //AXI-MM pass-through interface 113
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_113_AWADDR,
    input wire [7:0]                      AP_AXIMM_113_AWLEN,
    input wire [2:0]                      AP_AXIMM_113_AWSIZE,
    input wire [1:0]                      AP_AXIMM_113_AWBURST,
    input wire [1:0]                      AP_AXIMM_113_AWLOCK,
    input wire [3:0]                      AP_AXIMM_113_AWCACHE,
    input wire [2:0]                      AP_AXIMM_113_AWPROT,
    input wire [3:0]                      AP_AXIMM_113_AWREGION,
    input wire [3:0]                      AP_AXIMM_113_AWQOS,
    input wire                            AP_AXIMM_113_AWVALID,
    output  wire                            AP_AXIMM_113_AWREADY,
    input wire [M_AXIMM_113_DATA_WIDTH-1:0]   AP_AXIMM_113_WDATA,
    input wire [M_AXIMM_113_DATA_WIDTH/8-1:0] AP_AXIMM_113_WSTRB,
    input wire                            AP_AXIMM_113_WLAST,
    input wire                            AP_AXIMM_113_WVALID,
    output  wire                            AP_AXIMM_113_WREADY,
    output  wire [1:0]                      AP_AXIMM_113_BRESP,
    output  wire                            AP_AXIMM_113_BVALID,
    input wire                            AP_AXIMM_113_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_113_ARADDR,
    input wire [7:0]                      AP_AXIMM_113_ARLEN,
    input wire [2:0]                      AP_AXIMM_113_ARSIZE,
    input wire [1:0]                      AP_AXIMM_113_ARBURST,
    input wire [1:0]                      AP_AXIMM_113_ARLOCK,
    input wire [3:0]                      AP_AXIMM_113_ARCACHE,
    input wire [2:0]                      AP_AXIMM_113_ARPROT,
    input wire [3:0]                      AP_AXIMM_113_ARREGION,
    input wire [3:0]                      AP_AXIMM_113_ARQOS,
    input wire                            AP_AXIMM_113_ARVALID,
    output  wire                            AP_AXIMM_113_ARREADY,
    output  wire [M_AXIMM_113_DATA_WIDTH-1:0]   AP_AXIMM_113_RDATA,
    output  wire [1:0]                      AP_AXIMM_113_RRESP,
    output  wire                            AP_AXIMM_113_RLAST,
    output  wire                            AP_AXIMM_113_RVALID,
    input  wire                            AP_AXIMM_113_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_113_AWADDR,
    output wire [7:0]                      M_AXIMM_113_AWLEN,
    output wire [2:0]                      M_AXIMM_113_AWSIZE,
    output wire [1:0]                      M_AXIMM_113_AWBURST,
    output wire [1:0]                      M_AXIMM_113_AWLOCK,
    output wire [3:0]                      M_AXIMM_113_AWCACHE,
    output wire [2:0]                      M_AXIMM_113_AWPROT,
    output wire [3:0]                      M_AXIMM_113_AWREGION,
    output wire [3:0]                      M_AXIMM_113_AWQOS,
    output wire                            M_AXIMM_113_AWVALID,
    input  wire                            M_AXIMM_113_AWREADY,
    output wire [M_AXIMM_113_DATA_WIDTH-1:0]   M_AXIMM_113_WDATA,
    output wire [M_AXIMM_113_DATA_WIDTH/8-1:0] M_AXIMM_113_WSTRB,
    output wire                            M_AXIMM_113_WLAST,
    output wire                            M_AXIMM_113_WVALID,
    input  wire                            M_AXIMM_113_WREADY,
    input  wire [1:0]                      M_AXIMM_113_BRESP,
    input  wire                            M_AXIMM_113_BVALID,
    output wire                            M_AXIMM_113_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_113_ARADDR,
    output wire [7:0]                      M_AXIMM_113_ARLEN,
    output wire [2:0]                      M_AXIMM_113_ARSIZE,
    output wire [1:0]                      M_AXIMM_113_ARBURST,
    output wire [1:0]                      M_AXIMM_113_ARLOCK,
    output wire [3:0]                      M_AXIMM_113_ARCACHE,
    output wire [2:0]                      M_AXIMM_113_ARPROT,
    output wire [3:0]                      M_AXIMM_113_ARREGION,
    output wire [3:0]                      M_AXIMM_113_ARQOS,
    output wire                            M_AXIMM_113_ARVALID,
    input  wire                            M_AXIMM_113_ARREADY,
    input  wire [M_AXIMM_113_DATA_WIDTH-1:0]   M_AXIMM_113_RDATA,
    input  wire [1:0]                      M_AXIMM_113_RRESP,
    input  wire                            M_AXIMM_113_RLAST,
    input  wire                            M_AXIMM_113_RVALID,
    output wire                            M_AXIMM_113_RREADY,
    //AXI-MM pass-through interface 114
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_114_AWADDR,
    input wire [7:0]                      AP_AXIMM_114_AWLEN,
    input wire [2:0]                      AP_AXIMM_114_AWSIZE,
    input wire [1:0]                      AP_AXIMM_114_AWBURST,
    input wire [1:0]                      AP_AXIMM_114_AWLOCK,
    input wire [3:0]                      AP_AXIMM_114_AWCACHE,
    input wire [2:0]                      AP_AXIMM_114_AWPROT,
    input wire [3:0]                      AP_AXIMM_114_AWREGION,
    input wire [3:0]                      AP_AXIMM_114_AWQOS,
    input wire                            AP_AXIMM_114_AWVALID,
    output  wire                            AP_AXIMM_114_AWREADY,
    input wire [M_AXIMM_114_DATA_WIDTH-1:0]   AP_AXIMM_114_WDATA,
    input wire [M_AXIMM_114_DATA_WIDTH/8-1:0] AP_AXIMM_114_WSTRB,
    input wire                            AP_AXIMM_114_WLAST,
    input wire                            AP_AXIMM_114_WVALID,
    output  wire                            AP_AXIMM_114_WREADY,
    output  wire [1:0]                      AP_AXIMM_114_BRESP,
    output  wire                            AP_AXIMM_114_BVALID,
    input wire                            AP_AXIMM_114_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_114_ARADDR,
    input wire [7:0]                      AP_AXIMM_114_ARLEN,
    input wire [2:0]                      AP_AXIMM_114_ARSIZE,
    input wire [1:0]                      AP_AXIMM_114_ARBURST,
    input wire [1:0]                      AP_AXIMM_114_ARLOCK,
    input wire [3:0]                      AP_AXIMM_114_ARCACHE,
    input wire [2:0]                      AP_AXIMM_114_ARPROT,
    input wire [3:0]                      AP_AXIMM_114_ARREGION,
    input wire [3:0]                      AP_AXIMM_114_ARQOS,
    input wire                            AP_AXIMM_114_ARVALID,
    output  wire                            AP_AXIMM_114_ARREADY,
    output  wire [M_AXIMM_114_DATA_WIDTH-1:0]   AP_AXIMM_114_RDATA,
    output  wire [1:0]                      AP_AXIMM_114_RRESP,
    output  wire                            AP_AXIMM_114_RLAST,
    output  wire                            AP_AXIMM_114_RVALID,
    input  wire                            AP_AXIMM_114_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_114_AWADDR,
    output wire [7:0]                      M_AXIMM_114_AWLEN,
    output wire [2:0]                      M_AXIMM_114_AWSIZE,
    output wire [1:0]                      M_AXIMM_114_AWBURST,
    output wire [1:0]                      M_AXIMM_114_AWLOCK,
    output wire [3:0]                      M_AXIMM_114_AWCACHE,
    output wire [2:0]                      M_AXIMM_114_AWPROT,
    output wire [3:0]                      M_AXIMM_114_AWREGION,
    output wire [3:0]                      M_AXIMM_114_AWQOS,
    output wire                            M_AXIMM_114_AWVALID,
    input  wire                            M_AXIMM_114_AWREADY,
    output wire [M_AXIMM_114_DATA_WIDTH-1:0]   M_AXIMM_114_WDATA,
    output wire [M_AXIMM_114_DATA_WIDTH/8-1:0] M_AXIMM_114_WSTRB,
    output wire                            M_AXIMM_114_WLAST,
    output wire                            M_AXIMM_114_WVALID,
    input  wire                            M_AXIMM_114_WREADY,
    input  wire [1:0]                      M_AXIMM_114_BRESP,
    input  wire                            M_AXIMM_114_BVALID,
    output wire                            M_AXIMM_114_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_114_ARADDR,
    output wire [7:0]                      M_AXIMM_114_ARLEN,
    output wire [2:0]                      M_AXIMM_114_ARSIZE,
    output wire [1:0]                      M_AXIMM_114_ARBURST,
    output wire [1:0]                      M_AXIMM_114_ARLOCK,
    output wire [3:0]                      M_AXIMM_114_ARCACHE,
    output wire [2:0]                      M_AXIMM_114_ARPROT,
    output wire [3:0]                      M_AXIMM_114_ARREGION,
    output wire [3:0]                      M_AXIMM_114_ARQOS,
    output wire                            M_AXIMM_114_ARVALID,
    input  wire                            M_AXIMM_114_ARREADY,
    input  wire [M_AXIMM_114_DATA_WIDTH-1:0]   M_AXIMM_114_RDATA,
    input  wire [1:0]                      M_AXIMM_114_RRESP,
    input  wire                            M_AXIMM_114_RLAST,
    input  wire                            M_AXIMM_114_RVALID,
    output wire                            M_AXIMM_114_RREADY,
    //AXI-MM pass-through interface 115
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_115_AWADDR,
    input wire [7:0]                      AP_AXIMM_115_AWLEN,
    input wire [2:0]                      AP_AXIMM_115_AWSIZE,
    input wire [1:0]                      AP_AXIMM_115_AWBURST,
    input wire [1:0]                      AP_AXIMM_115_AWLOCK,
    input wire [3:0]                      AP_AXIMM_115_AWCACHE,
    input wire [2:0]                      AP_AXIMM_115_AWPROT,
    input wire [3:0]                      AP_AXIMM_115_AWREGION,
    input wire [3:0]                      AP_AXIMM_115_AWQOS,
    input wire                            AP_AXIMM_115_AWVALID,
    output  wire                            AP_AXIMM_115_AWREADY,
    input wire [M_AXIMM_115_DATA_WIDTH-1:0]   AP_AXIMM_115_WDATA,
    input wire [M_AXIMM_115_DATA_WIDTH/8-1:0] AP_AXIMM_115_WSTRB,
    input wire                            AP_AXIMM_115_WLAST,
    input wire                            AP_AXIMM_115_WVALID,
    output  wire                            AP_AXIMM_115_WREADY,
    output  wire [1:0]                      AP_AXIMM_115_BRESP,
    output  wire                            AP_AXIMM_115_BVALID,
    input wire                            AP_AXIMM_115_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_115_ARADDR,
    input wire [7:0]                      AP_AXIMM_115_ARLEN,
    input wire [2:0]                      AP_AXIMM_115_ARSIZE,
    input wire [1:0]                      AP_AXIMM_115_ARBURST,
    input wire [1:0]                      AP_AXIMM_115_ARLOCK,
    input wire [3:0]                      AP_AXIMM_115_ARCACHE,
    input wire [2:0]                      AP_AXIMM_115_ARPROT,
    input wire [3:0]                      AP_AXIMM_115_ARREGION,
    input wire [3:0]                      AP_AXIMM_115_ARQOS,
    input wire                            AP_AXIMM_115_ARVALID,
    output  wire                            AP_AXIMM_115_ARREADY,
    output  wire [M_AXIMM_115_DATA_WIDTH-1:0]   AP_AXIMM_115_RDATA,
    output  wire [1:0]                      AP_AXIMM_115_RRESP,
    output  wire                            AP_AXIMM_115_RLAST,
    output  wire                            AP_AXIMM_115_RVALID,
    input  wire                            AP_AXIMM_115_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_115_AWADDR,
    output wire [7:0]                      M_AXIMM_115_AWLEN,
    output wire [2:0]                      M_AXIMM_115_AWSIZE,
    output wire [1:0]                      M_AXIMM_115_AWBURST,
    output wire [1:0]                      M_AXIMM_115_AWLOCK,
    output wire [3:0]                      M_AXIMM_115_AWCACHE,
    output wire [2:0]                      M_AXIMM_115_AWPROT,
    output wire [3:0]                      M_AXIMM_115_AWREGION,
    output wire [3:0]                      M_AXIMM_115_AWQOS,
    output wire                            M_AXIMM_115_AWVALID,
    input  wire                            M_AXIMM_115_AWREADY,
    output wire [M_AXIMM_115_DATA_WIDTH-1:0]   M_AXIMM_115_WDATA,
    output wire [M_AXIMM_115_DATA_WIDTH/8-1:0] M_AXIMM_115_WSTRB,
    output wire                            M_AXIMM_115_WLAST,
    output wire                            M_AXIMM_115_WVALID,
    input  wire                            M_AXIMM_115_WREADY,
    input  wire [1:0]                      M_AXIMM_115_BRESP,
    input  wire                            M_AXIMM_115_BVALID,
    output wire                            M_AXIMM_115_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_115_ARADDR,
    output wire [7:0]                      M_AXIMM_115_ARLEN,
    output wire [2:0]                      M_AXIMM_115_ARSIZE,
    output wire [1:0]                      M_AXIMM_115_ARBURST,
    output wire [1:0]                      M_AXIMM_115_ARLOCK,
    output wire [3:0]                      M_AXIMM_115_ARCACHE,
    output wire [2:0]                      M_AXIMM_115_ARPROT,
    output wire [3:0]                      M_AXIMM_115_ARREGION,
    output wire [3:0]                      M_AXIMM_115_ARQOS,
    output wire                            M_AXIMM_115_ARVALID,
    input  wire                            M_AXIMM_115_ARREADY,
    input  wire [M_AXIMM_115_DATA_WIDTH-1:0]   M_AXIMM_115_RDATA,
    input  wire [1:0]                      M_AXIMM_115_RRESP,
    input  wire                            M_AXIMM_115_RLAST,
    input  wire                            M_AXIMM_115_RVALID,
    output wire                            M_AXIMM_115_RREADY,
    //AXI-MM pass-through interface 116
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_116_AWADDR,
    input wire [7:0]                      AP_AXIMM_116_AWLEN,
    input wire [2:0]                      AP_AXIMM_116_AWSIZE,
    input wire [1:0]                      AP_AXIMM_116_AWBURST,
    input wire [1:0]                      AP_AXIMM_116_AWLOCK,
    input wire [3:0]                      AP_AXIMM_116_AWCACHE,
    input wire [2:0]                      AP_AXIMM_116_AWPROT,
    input wire [3:0]                      AP_AXIMM_116_AWREGION,
    input wire [3:0]                      AP_AXIMM_116_AWQOS,
    input wire                            AP_AXIMM_116_AWVALID,
    output  wire                            AP_AXIMM_116_AWREADY,
    input wire [M_AXIMM_116_DATA_WIDTH-1:0]   AP_AXIMM_116_WDATA,
    input wire [M_AXIMM_116_DATA_WIDTH/8-1:0] AP_AXIMM_116_WSTRB,
    input wire                            AP_AXIMM_116_WLAST,
    input wire                            AP_AXIMM_116_WVALID,
    output  wire                            AP_AXIMM_116_WREADY,
    output  wire [1:0]                      AP_AXIMM_116_BRESP,
    output  wire                            AP_AXIMM_116_BVALID,
    input wire                            AP_AXIMM_116_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_116_ARADDR,
    input wire [7:0]                      AP_AXIMM_116_ARLEN,
    input wire [2:0]                      AP_AXIMM_116_ARSIZE,
    input wire [1:0]                      AP_AXIMM_116_ARBURST,
    input wire [1:0]                      AP_AXIMM_116_ARLOCK,
    input wire [3:0]                      AP_AXIMM_116_ARCACHE,
    input wire [2:0]                      AP_AXIMM_116_ARPROT,
    input wire [3:0]                      AP_AXIMM_116_ARREGION,
    input wire [3:0]                      AP_AXIMM_116_ARQOS,
    input wire                            AP_AXIMM_116_ARVALID,
    output  wire                            AP_AXIMM_116_ARREADY,
    output  wire [M_AXIMM_116_DATA_WIDTH-1:0]   AP_AXIMM_116_RDATA,
    output  wire [1:0]                      AP_AXIMM_116_RRESP,
    output  wire                            AP_AXIMM_116_RLAST,
    output  wire                            AP_AXIMM_116_RVALID,
    input  wire                            AP_AXIMM_116_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_116_AWADDR,
    output wire [7:0]                      M_AXIMM_116_AWLEN,
    output wire [2:0]                      M_AXIMM_116_AWSIZE,
    output wire [1:0]                      M_AXIMM_116_AWBURST,
    output wire [1:0]                      M_AXIMM_116_AWLOCK,
    output wire [3:0]                      M_AXIMM_116_AWCACHE,
    output wire [2:0]                      M_AXIMM_116_AWPROT,
    output wire [3:0]                      M_AXIMM_116_AWREGION,
    output wire [3:0]                      M_AXIMM_116_AWQOS,
    output wire                            M_AXIMM_116_AWVALID,
    input  wire                            M_AXIMM_116_AWREADY,
    output wire [M_AXIMM_116_DATA_WIDTH-1:0]   M_AXIMM_116_WDATA,
    output wire [M_AXIMM_116_DATA_WIDTH/8-1:0] M_AXIMM_116_WSTRB,
    output wire                            M_AXIMM_116_WLAST,
    output wire                            M_AXIMM_116_WVALID,
    input  wire                            M_AXIMM_116_WREADY,
    input  wire [1:0]                      M_AXIMM_116_BRESP,
    input  wire                            M_AXIMM_116_BVALID,
    output wire                            M_AXIMM_116_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_116_ARADDR,
    output wire [7:0]                      M_AXIMM_116_ARLEN,
    output wire [2:0]                      M_AXIMM_116_ARSIZE,
    output wire [1:0]                      M_AXIMM_116_ARBURST,
    output wire [1:0]                      M_AXIMM_116_ARLOCK,
    output wire [3:0]                      M_AXIMM_116_ARCACHE,
    output wire [2:0]                      M_AXIMM_116_ARPROT,
    output wire [3:0]                      M_AXIMM_116_ARREGION,
    output wire [3:0]                      M_AXIMM_116_ARQOS,
    output wire                            M_AXIMM_116_ARVALID,
    input  wire                            M_AXIMM_116_ARREADY,
    input  wire [M_AXIMM_116_DATA_WIDTH-1:0]   M_AXIMM_116_RDATA,
    input  wire [1:0]                      M_AXIMM_116_RRESP,
    input  wire                            M_AXIMM_116_RLAST,
    input  wire                            M_AXIMM_116_RVALID,
    output wire                            M_AXIMM_116_RREADY,
    //AXI-MM pass-through interface 117
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_117_AWADDR,
    input wire [7:0]                      AP_AXIMM_117_AWLEN,
    input wire [2:0]                      AP_AXIMM_117_AWSIZE,
    input wire [1:0]                      AP_AXIMM_117_AWBURST,
    input wire [1:0]                      AP_AXIMM_117_AWLOCK,
    input wire [3:0]                      AP_AXIMM_117_AWCACHE,
    input wire [2:0]                      AP_AXIMM_117_AWPROT,
    input wire [3:0]                      AP_AXIMM_117_AWREGION,
    input wire [3:0]                      AP_AXIMM_117_AWQOS,
    input wire                            AP_AXIMM_117_AWVALID,
    output  wire                            AP_AXIMM_117_AWREADY,
    input wire [M_AXIMM_117_DATA_WIDTH-1:0]   AP_AXIMM_117_WDATA,
    input wire [M_AXIMM_117_DATA_WIDTH/8-1:0] AP_AXIMM_117_WSTRB,
    input wire                            AP_AXIMM_117_WLAST,
    input wire                            AP_AXIMM_117_WVALID,
    output  wire                            AP_AXIMM_117_WREADY,
    output  wire [1:0]                      AP_AXIMM_117_BRESP,
    output  wire                            AP_AXIMM_117_BVALID,
    input wire                            AP_AXIMM_117_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_117_ARADDR,
    input wire [7:0]                      AP_AXIMM_117_ARLEN,
    input wire [2:0]                      AP_AXIMM_117_ARSIZE,
    input wire [1:0]                      AP_AXIMM_117_ARBURST,
    input wire [1:0]                      AP_AXIMM_117_ARLOCK,
    input wire [3:0]                      AP_AXIMM_117_ARCACHE,
    input wire [2:0]                      AP_AXIMM_117_ARPROT,
    input wire [3:0]                      AP_AXIMM_117_ARREGION,
    input wire [3:0]                      AP_AXIMM_117_ARQOS,
    input wire                            AP_AXIMM_117_ARVALID,
    output  wire                            AP_AXIMM_117_ARREADY,
    output  wire [M_AXIMM_117_DATA_WIDTH-1:0]   AP_AXIMM_117_RDATA,
    output  wire [1:0]                      AP_AXIMM_117_RRESP,
    output  wire                            AP_AXIMM_117_RLAST,
    output  wire                            AP_AXIMM_117_RVALID,
    input  wire                            AP_AXIMM_117_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_117_AWADDR,
    output wire [7:0]                      M_AXIMM_117_AWLEN,
    output wire [2:0]                      M_AXIMM_117_AWSIZE,
    output wire [1:0]                      M_AXIMM_117_AWBURST,
    output wire [1:0]                      M_AXIMM_117_AWLOCK,
    output wire [3:0]                      M_AXIMM_117_AWCACHE,
    output wire [2:0]                      M_AXIMM_117_AWPROT,
    output wire [3:0]                      M_AXIMM_117_AWREGION,
    output wire [3:0]                      M_AXIMM_117_AWQOS,
    output wire                            M_AXIMM_117_AWVALID,
    input  wire                            M_AXIMM_117_AWREADY,
    output wire [M_AXIMM_117_DATA_WIDTH-1:0]   M_AXIMM_117_WDATA,
    output wire [M_AXIMM_117_DATA_WIDTH/8-1:0] M_AXIMM_117_WSTRB,
    output wire                            M_AXIMM_117_WLAST,
    output wire                            M_AXIMM_117_WVALID,
    input  wire                            M_AXIMM_117_WREADY,
    input  wire [1:0]                      M_AXIMM_117_BRESP,
    input  wire                            M_AXIMM_117_BVALID,
    output wire                            M_AXIMM_117_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_117_ARADDR,
    output wire [7:0]                      M_AXIMM_117_ARLEN,
    output wire [2:0]                      M_AXIMM_117_ARSIZE,
    output wire [1:0]                      M_AXIMM_117_ARBURST,
    output wire [1:0]                      M_AXIMM_117_ARLOCK,
    output wire [3:0]                      M_AXIMM_117_ARCACHE,
    output wire [2:0]                      M_AXIMM_117_ARPROT,
    output wire [3:0]                      M_AXIMM_117_ARREGION,
    output wire [3:0]                      M_AXIMM_117_ARQOS,
    output wire                            M_AXIMM_117_ARVALID,
    input  wire                            M_AXIMM_117_ARREADY,
    input  wire [M_AXIMM_117_DATA_WIDTH-1:0]   M_AXIMM_117_RDATA,
    input  wire [1:0]                      M_AXIMM_117_RRESP,
    input  wire                            M_AXIMM_117_RLAST,
    input  wire                            M_AXIMM_117_RVALID,
    output wire                            M_AXIMM_117_RREADY,
    //AXI-MM pass-through interface 118
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_118_AWADDR,
    input wire [7:0]                      AP_AXIMM_118_AWLEN,
    input wire [2:0]                      AP_AXIMM_118_AWSIZE,
    input wire [1:0]                      AP_AXIMM_118_AWBURST,
    input wire [1:0]                      AP_AXIMM_118_AWLOCK,
    input wire [3:0]                      AP_AXIMM_118_AWCACHE,
    input wire [2:0]                      AP_AXIMM_118_AWPROT,
    input wire [3:0]                      AP_AXIMM_118_AWREGION,
    input wire [3:0]                      AP_AXIMM_118_AWQOS,
    input wire                            AP_AXIMM_118_AWVALID,
    output  wire                            AP_AXIMM_118_AWREADY,
    input wire [M_AXIMM_118_DATA_WIDTH-1:0]   AP_AXIMM_118_WDATA,
    input wire [M_AXIMM_118_DATA_WIDTH/8-1:0] AP_AXIMM_118_WSTRB,
    input wire                            AP_AXIMM_118_WLAST,
    input wire                            AP_AXIMM_118_WVALID,
    output  wire                            AP_AXIMM_118_WREADY,
    output  wire [1:0]                      AP_AXIMM_118_BRESP,
    output  wire                            AP_AXIMM_118_BVALID,
    input wire                            AP_AXIMM_118_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_118_ARADDR,
    input wire [7:0]                      AP_AXIMM_118_ARLEN,
    input wire [2:0]                      AP_AXIMM_118_ARSIZE,
    input wire [1:0]                      AP_AXIMM_118_ARBURST,
    input wire [1:0]                      AP_AXIMM_118_ARLOCK,
    input wire [3:0]                      AP_AXIMM_118_ARCACHE,
    input wire [2:0]                      AP_AXIMM_118_ARPROT,
    input wire [3:0]                      AP_AXIMM_118_ARREGION,
    input wire [3:0]                      AP_AXIMM_118_ARQOS,
    input wire                            AP_AXIMM_118_ARVALID,
    output  wire                            AP_AXIMM_118_ARREADY,
    output  wire [M_AXIMM_118_DATA_WIDTH-1:0]   AP_AXIMM_118_RDATA,
    output  wire [1:0]                      AP_AXIMM_118_RRESP,
    output  wire                            AP_AXIMM_118_RLAST,
    output  wire                            AP_AXIMM_118_RVALID,
    input  wire                            AP_AXIMM_118_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_118_AWADDR,
    output wire [7:0]                      M_AXIMM_118_AWLEN,
    output wire [2:0]                      M_AXIMM_118_AWSIZE,
    output wire [1:0]                      M_AXIMM_118_AWBURST,
    output wire [1:0]                      M_AXIMM_118_AWLOCK,
    output wire [3:0]                      M_AXIMM_118_AWCACHE,
    output wire [2:0]                      M_AXIMM_118_AWPROT,
    output wire [3:0]                      M_AXIMM_118_AWREGION,
    output wire [3:0]                      M_AXIMM_118_AWQOS,
    output wire                            M_AXIMM_118_AWVALID,
    input  wire                            M_AXIMM_118_AWREADY,
    output wire [M_AXIMM_118_DATA_WIDTH-1:0]   M_AXIMM_118_WDATA,
    output wire [M_AXIMM_118_DATA_WIDTH/8-1:0] M_AXIMM_118_WSTRB,
    output wire                            M_AXIMM_118_WLAST,
    output wire                            M_AXIMM_118_WVALID,
    input  wire                            M_AXIMM_118_WREADY,
    input  wire [1:0]                      M_AXIMM_118_BRESP,
    input  wire                            M_AXIMM_118_BVALID,
    output wire                            M_AXIMM_118_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_118_ARADDR,
    output wire [7:0]                      M_AXIMM_118_ARLEN,
    output wire [2:0]                      M_AXIMM_118_ARSIZE,
    output wire [1:0]                      M_AXIMM_118_ARBURST,
    output wire [1:0]                      M_AXIMM_118_ARLOCK,
    output wire [3:0]                      M_AXIMM_118_ARCACHE,
    output wire [2:0]                      M_AXIMM_118_ARPROT,
    output wire [3:0]                      M_AXIMM_118_ARREGION,
    output wire [3:0]                      M_AXIMM_118_ARQOS,
    output wire                            M_AXIMM_118_ARVALID,
    input  wire                            M_AXIMM_118_ARREADY,
    input  wire [M_AXIMM_118_DATA_WIDTH-1:0]   M_AXIMM_118_RDATA,
    input  wire [1:0]                      M_AXIMM_118_RRESP,
    input  wire                            M_AXIMM_118_RLAST,
    input  wire                            M_AXIMM_118_RVALID,
    output wire                            M_AXIMM_118_RREADY,
    //AXI-MM pass-through interface 119
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_119_AWADDR,
    input wire [7:0]                      AP_AXIMM_119_AWLEN,
    input wire [2:0]                      AP_AXIMM_119_AWSIZE,
    input wire [1:0]                      AP_AXIMM_119_AWBURST,
    input wire [1:0]                      AP_AXIMM_119_AWLOCK,
    input wire [3:0]                      AP_AXIMM_119_AWCACHE,
    input wire [2:0]                      AP_AXIMM_119_AWPROT,
    input wire [3:0]                      AP_AXIMM_119_AWREGION,
    input wire [3:0]                      AP_AXIMM_119_AWQOS,
    input wire                            AP_AXIMM_119_AWVALID,
    output  wire                            AP_AXIMM_119_AWREADY,
    input wire [M_AXIMM_119_DATA_WIDTH-1:0]   AP_AXIMM_119_WDATA,
    input wire [M_AXIMM_119_DATA_WIDTH/8-1:0] AP_AXIMM_119_WSTRB,
    input wire                            AP_AXIMM_119_WLAST,
    input wire                            AP_AXIMM_119_WVALID,
    output  wire                            AP_AXIMM_119_WREADY,
    output  wire [1:0]                      AP_AXIMM_119_BRESP,
    output  wire                            AP_AXIMM_119_BVALID,
    input wire                            AP_AXIMM_119_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_119_ARADDR,
    input wire [7:0]                      AP_AXIMM_119_ARLEN,
    input wire [2:0]                      AP_AXIMM_119_ARSIZE,
    input wire [1:0]                      AP_AXIMM_119_ARBURST,
    input wire [1:0]                      AP_AXIMM_119_ARLOCK,
    input wire [3:0]                      AP_AXIMM_119_ARCACHE,
    input wire [2:0]                      AP_AXIMM_119_ARPROT,
    input wire [3:0]                      AP_AXIMM_119_ARREGION,
    input wire [3:0]                      AP_AXIMM_119_ARQOS,
    input wire                            AP_AXIMM_119_ARVALID,
    output  wire                            AP_AXIMM_119_ARREADY,
    output  wire [M_AXIMM_119_DATA_WIDTH-1:0]   AP_AXIMM_119_RDATA,
    output  wire [1:0]                      AP_AXIMM_119_RRESP,
    output  wire                            AP_AXIMM_119_RLAST,
    output  wire                            AP_AXIMM_119_RVALID,
    input  wire                            AP_AXIMM_119_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_119_AWADDR,
    output wire [7:0]                      M_AXIMM_119_AWLEN,
    output wire [2:0]                      M_AXIMM_119_AWSIZE,
    output wire [1:0]                      M_AXIMM_119_AWBURST,
    output wire [1:0]                      M_AXIMM_119_AWLOCK,
    output wire [3:0]                      M_AXIMM_119_AWCACHE,
    output wire [2:0]                      M_AXIMM_119_AWPROT,
    output wire [3:0]                      M_AXIMM_119_AWREGION,
    output wire [3:0]                      M_AXIMM_119_AWQOS,
    output wire                            M_AXIMM_119_AWVALID,
    input  wire                            M_AXIMM_119_AWREADY,
    output wire [M_AXIMM_119_DATA_WIDTH-1:0]   M_AXIMM_119_WDATA,
    output wire [M_AXIMM_119_DATA_WIDTH/8-1:0] M_AXIMM_119_WSTRB,
    output wire                            M_AXIMM_119_WLAST,
    output wire                            M_AXIMM_119_WVALID,
    input  wire                            M_AXIMM_119_WREADY,
    input  wire [1:0]                      M_AXIMM_119_BRESP,
    input  wire                            M_AXIMM_119_BVALID,
    output wire                            M_AXIMM_119_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_119_ARADDR,
    output wire [7:0]                      M_AXIMM_119_ARLEN,
    output wire [2:0]                      M_AXIMM_119_ARSIZE,
    output wire [1:0]                      M_AXIMM_119_ARBURST,
    output wire [1:0]                      M_AXIMM_119_ARLOCK,
    output wire [3:0]                      M_AXIMM_119_ARCACHE,
    output wire [2:0]                      M_AXIMM_119_ARPROT,
    output wire [3:0]                      M_AXIMM_119_ARREGION,
    output wire [3:0]                      M_AXIMM_119_ARQOS,
    output wire                            M_AXIMM_119_ARVALID,
    input  wire                            M_AXIMM_119_ARREADY,
    input  wire [M_AXIMM_119_DATA_WIDTH-1:0]   M_AXIMM_119_RDATA,
    input  wire [1:0]                      M_AXIMM_119_RRESP,
    input  wire                            M_AXIMM_119_RLAST,
    input  wire                            M_AXIMM_119_RVALID,
    output wire                            M_AXIMM_119_RREADY,
    //AXI-MM pass-through interface 120
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_120_AWADDR,
    input wire [7:0]                      AP_AXIMM_120_AWLEN,
    input wire [2:0]                      AP_AXIMM_120_AWSIZE,
    input wire [1:0]                      AP_AXIMM_120_AWBURST,
    input wire [1:0]                      AP_AXIMM_120_AWLOCK,
    input wire [3:0]                      AP_AXIMM_120_AWCACHE,
    input wire [2:0]                      AP_AXIMM_120_AWPROT,
    input wire [3:0]                      AP_AXIMM_120_AWREGION,
    input wire [3:0]                      AP_AXIMM_120_AWQOS,
    input wire                            AP_AXIMM_120_AWVALID,
    output  wire                            AP_AXIMM_120_AWREADY,
    input wire [M_AXIMM_120_DATA_WIDTH-1:0]   AP_AXIMM_120_WDATA,
    input wire [M_AXIMM_120_DATA_WIDTH/8-1:0] AP_AXIMM_120_WSTRB,
    input wire                            AP_AXIMM_120_WLAST,
    input wire                            AP_AXIMM_120_WVALID,
    output  wire                            AP_AXIMM_120_WREADY,
    output  wire [1:0]                      AP_AXIMM_120_BRESP,
    output  wire                            AP_AXIMM_120_BVALID,
    input wire                            AP_AXIMM_120_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_120_ARADDR,
    input wire [7:0]                      AP_AXIMM_120_ARLEN,
    input wire [2:0]                      AP_AXIMM_120_ARSIZE,
    input wire [1:0]                      AP_AXIMM_120_ARBURST,
    input wire [1:0]                      AP_AXIMM_120_ARLOCK,
    input wire [3:0]                      AP_AXIMM_120_ARCACHE,
    input wire [2:0]                      AP_AXIMM_120_ARPROT,
    input wire [3:0]                      AP_AXIMM_120_ARREGION,
    input wire [3:0]                      AP_AXIMM_120_ARQOS,
    input wire                            AP_AXIMM_120_ARVALID,
    output  wire                            AP_AXIMM_120_ARREADY,
    output  wire [M_AXIMM_120_DATA_WIDTH-1:0]   AP_AXIMM_120_RDATA,
    output  wire [1:0]                      AP_AXIMM_120_RRESP,
    output  wire                            AP_AXIMM_120_RLAST,
    output  wire                            AP_AXIMM_120_RVALID,
    input  wire                            AP_AXIMM_120_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_120_AWADDR,
    output wire [7:0]                      M_AXIMM_120_AWLEN,
    output wire [2:0]                      M_AXIMM_120_AWSIZE,
    output wire [1:0]                      M_AXIMM_120_AWBURST,
    output wire [1:0]                      M_AXIMM_120_AWLOCK,
    output wire [3:0]                      M_AXIMM_120_AWCACHE,
    output wire [2:0]                      M_AXIMM_120_AWPROT,
    output wire [3:0]                      M_AXIMM_120_AWREGION,
    output wire [3:0]                      M_AXIMM_120_AWQOS,
    output wire                            M_AXIMM_120_AWVALID,
    input  wire                            M_AXIMM_120_AWREADY,
    output wire [M_AXIMM_120_DATA_WIDTH-1:0]   M_AXIMM_120_WDATA,
    output wire [M_AXIMM_120_DATA_WIDTH/8-1:0] M_AXIMM_120_WSTRB,
    output wire                            M_AXIMM_120_WLAST,
    output wire                            M_AXIMM_120_WVALID,
    input  wire                            M_AXIMM_120_WREADY,
    input  wire [1:0]                      M_AXIMM_120_BRESP,
    input  wire                            M_AXIMM_120_BVALID,
    output wire                            M_AXIMM_120_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_120_ARADDR,
    output wire [7:0]                      M_AXIMM_120_ARLEN,
    output wire [2:0]                      M_AXIMM_120_ARSIZE,
    output wire [1:0]                      M_AXIMM_120_ARBURST,
    output wire [1:0]                      M_AXIMM_120_ARLOCK,
    output wire [3:0]                      M_AXIMM_120_ARCACHE,
    output wire [2:0]                      M_AXIMM_120_ARPROT,
    output wire [3:0]                      M_AXIMM_120_ARREGION,
    output wire [3:0]                      M_AXIMM_120_ARQOS,
    output wire                            M_AXIMM_120_ARVALID,
    input  wire                            M_AXIMM_120_ARREADY,
    input  wire [M_AXIMM_120_DATA_WIDTH-1:0]   M_AXIMM_120_RDATA,
    input  wire [1:0]                      M_AXIMM_120_RRESP,
    input  wire                            M_AXIMM_120_RLAST,
    input  wire                            M_AXIMM_120_RVALID,
    output wire                            M_AXIMM_120_RREADY,
    //AXI-MM pass-through interface 121
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_121_AWADDR,
    input wire [7:0]                      AP_AXIMM_121_AWLEN,
    input wire [2:0]                      AP_AXIMM_121_AWSIZE,
    input wire [1:0]                      AP_AXIMM_121_AWBURST,
    input wire [1:0]                      AP_AXIMM_121_AWLOCK,
    input wire [3:0]                      AP_AXIMM_121_AWCACHE,
    input wire [2:0]                      AP_AXIMM_121_AWPROT,
    input wire [3:0]                      AP_AXIMM_121_AWREGION,
    input wire [3:0]                      AP_AXIMM_121_AWQOS,
    input wire                            AP_AXIMM_121_AWVALID,
    output  wire                            AP_AXIMM_121_AWREADY,
    input wire [M_AXIMM_121_DATA_WIDTH-1:0]   AP_AXIMM_121_WDATA,
    input wire [M_AXIMM_121_DATA_WIDTH/8-1:0] AP_AXIMM_121_WSTRB,
    input wire                            AP_AXIMM_121_WLAST,
    input wire                            AP_AXIMM_121_WVALID,
    output  wire                            AP_AXIMM_121_WREADY,
    output  wire [1:0]                      AP_AXIMM_121_BRESP,
    output  wire                            AP_AXIMM_121_BVALID,
    input wire                            AP_AXIMM_121_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_121_ARADDR,
    input wire [7:0]                      AP_AXIMM_121_ARLEN,
    input wire [2:0]                      AP_AXIMM_121_ARSIZE,
    input wire [1:0]                      AP_AXIMM_121_ARBURST,
    input wire [1:0]                      AP_AXIMM_121_ARLOCK,
    input wire [3:0]                      AP_AXIMM_121_ARCACHE,
    input wire [2:0]                      AP_AXIMM_121_ARPROT,
    input wire [3:0]                      AP_AXIMM_121_ARREGION,
    input wire [3:0]                      AP_AXIMM_121_ARQOS,
    input wire                            AP_AXIMM_121_ARVALID,
    output  wire                            AP_AXIMM_121_ARREADY,
    output  wire [M_AXIMM_121_DATA_WIDTH-1:0]   AP_AXIMM_121_RDATA,
    output  wire [1:0]                      AP_AXIMM_121_RRESP,
    output  wire                            AP_AXIMM_121_RLAST,
    output  wire                            AP_AXIMM_121_RVALID,
    input  wire                            AP_AXIMM_121_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_121_AWADDR,
    output wire [7:0]                      M_AXIMM_121_AWLEN,
    output wire [2:0]                      M_AXIMM_121_AWSIZE,
    output wire [1:0]                      M_AXIMM_121_AWBURST,
    output wire [1:0]                      M_AXIMM_121_AWLOCK,
    output wire [3:0]                      M_AXIMM_121_AWCACHE,
    output wire [2:0]                      M_AXIMM_121_AWPROT,
    output wire [3:0]                      M_AXIMM_121_AWREGION,
    output wire [3:0]                      M_AXIMM_121_AWQOS,
    output wire                            M_AXIMM_121_AWVALID,
    input  wire                            M_AXIMM_121_AWREADY,
    output wire [M_AXIMM_121_DATA_WIDTH-1:0]   M_AXIMM_121_WDATA,
    output wire [M_AXIMM_121_DATA_WIDTH/8-1:0] M_AXIMM_121_WSTRB,
    output wire                            M_AXIMM_121_WLAST,
    output wire                            M_AXIMM_121_WVALID,
    input  wire                            M_AXIMM_121_WREADY,
    input  wire [1:0]                      M_AXIMM_121_BRESP,
    input  wire                            M_AXIMM_121_BVALID,
    output wire                            M_AXIMM_121_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_121_ARADDR,
    output wire [7:0]                      M_AXIMM_121_ARLEN,
    output wire [2:0]                      M_AXIMM_121_ARSIZE,
    output wire [1:0]                      M_AXIMM_121_ARBURST,
    output wire [1:0]                      M_AXIMM_121_ARLOCK,
    output wire [3:0]                      M_AXIMM_121_ARCACHE,
    output wire [2:0]                      M_AXIMM_121_ARPROT,
    output wire [3:0]                      M_AXIMM_121_ARREGION,
    output wire [3:0]                      M_AXIMM_121_ARQOS,
    output wire                            M_AXIMM_121_ARVALID,
    input  wire                            M_AXIMM_121_ARREADY,
    input  wire [M_AXIMM_121_DATA_WIDTH-1:0]   M_AXIMM_121_RDATA,
    input  wire [1:0]                      M_AXIMM_121_RRESP,
    input  wire                            M_AXIMM_121_RLAST,
    input  wire                            M_AXIMM_121_RVALID,
    output wire                            M_AXIMM_121_RREADY,
    //AXI-MM pass-through interface 122
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_122_AWADDR,
    input wire [7:0]                      AP_AXIMM_122_AWLEN,
    input wire [2:0]                      AP_AXIMM_122_AWSIZE,
    input wire [1:0]                      AP_AXIMM_122_AWBURST,
    input wire [1:0]                      AP_AXIMM_122_AWLOCK,
    input wire [3:0]                      AP_AXIMM_122_AWCACHE,
    input wire [2:0]                      AP_AXIMM_122_AWPROT,
    input wire [3:0]                      AP_AXIMM_122_AWREGION,
    input wire [3:0]                      AP_AXIMM_122_AWQOS,
    input wire                            AP_AXIMM_122_AWVALID,
    output  wire                            AP_AXIMM_122_AWREADY,
    input wire [M_AXIMM_122_DATA_WIDTH-1:0]   AP_AXIMM_122_WDATA,
    input wire [M_AXIMM_122_DATA_WIDTH/8-1:0] AP_AXIMM_122_WSTRB,
    input wire                            AP_AXIMM_122_WLAST,
    input wire                            AP_AXIMM_122_WVALID,
    output  wire                            AP_AXIMM_122_WREADY,
    output  wire [1:0]                      AP_AXIMM_122_BRESP,
    output  wire                            AP_AXIMM_122_BVALID,
    input wire                            AP_AXIMM_122_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_122_ARADDR,
    input wire [7:0]                      AP_AXIMM_122_ARLEN,
    input wire [2:0]                      AP_AXIMM_122_ARSIZE,
    input wire [1:0]                      AP_AXIMM_122_ARBURST,
    input wire [1:0]                      AP_AXIMM_122_ARLOCK,
    input wire [3:0]                      AP_AXIMM_122_ARCACHE,
    input wire [2:0]                      AP_AXIMM_122_ARPROT,
    input wire [3:0]                      AP_AXIMM_122_ARREGION,
    input wire [3:0]                      AP_AXIMM_122_ARQOS,
    input wire                            AP_AXIMM_122_ARVALID,
    output  wire                            AP_AXIMM_122_ARREADY,
    output  wire [M_AXIMM_122_DATA_WIDTH-1:0]   AP_AXIMM_122_RDATA,
    output  wire [1:0]                      AP_AXIMM_122_RRESP,
    output  wire                            AP_AXIMM_122_RLAST,
    output  wire                            AP_AXIMM_122_RVALID,
    input  wire                            AP_AXIMM_122_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_122_AWADDR,
    output wire [7:0]                      M_AXIMM_122_AWLEN,
    output wire [2:0]                      M_AXIMM_122_AWSIZE,
    output wire [1:0]                      M_AXIMM_122_AWBURST,
    output wire [1:0]                      M_AXIMM_122_AWLOCK,
    output wire [3:0]                      M_AXIMM_122_AWCACHE,
    output wire [2:0]                      M_AXIMM_122_AWPROT,
    output wire [3:0]                      M_AXIMM_122_AWREGION,
    output wire [3:0]                      M_AXIMM_122_AWQOS,
    output wire                            M_AXIMM_122_AWVALID,
    input  wire                            M_AXIMM_122_AWREADY,
    output wire [M_AXIMM_122_DATA_WIDTH-1:0]   M_AXIMM_122_WDATA,
    output wire [M_AXIMM_122_DATA_WIDTH/8-1:0] M_AXIMM_122_WSTRB,
    output wire                            M_AXIMM_122_WLAST,
    output wire                            M_AXIMM_122_WVALID,
    input  wire                            M_AXIMM_122_WREADY,
    input  wire [1:0]                      M_AXIMM_122_BRESP,
    input  wire                            M_AXIMM_122_BVALID,
    output wire                            M_AXIMM_122_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_122_ARADDR,
    output wire [7:0]                      M_AXIMM_122_ARLEN,
    output wire [2:0]                      M_AXIMM_122_ARSIZE,
    output wire [1:0]                      M_AXIMM_122_ARBURST,
    output wire [1:0]                      M_AXIMM_122_ARLOCK,
    output wire [3:0]                      M_AXIMM_122_ARCACHE,
    output wire [2:0]                      M_AXIMM_122_ARPROT,
    output wire [3:0]                      M_AXIMM_122_ARREGION,
    output wire [3:0]                      M_AXIMM_122_ARQOS,
    output wire                            M_AXIMM_122_ARVALID,
    input  wire                            M_AXIMM_122_ARREADY,
    input  wire [M_AXIMM_122_DATA_WIDTH-1:0]   M_AXIMM_122_RDATA,
    input  wire [1:0]                      M_AXIMM_122_RRESP,
    input  wire                            M_AXIMM_122_RLAST,
    input  wire                            M_AXIMM_122_RVALID,
    output wire                            M_AXIMM_122_RREADY,
    //AXI-MM pass-through interface 123
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_123_AWADDR,
    input wire [7:0]                      AP_AXIMM_123_AWLEN,
    input wire [2:0]                      AP_AXIMM_123_AWSIZE,
    input wire [1:0]                      AP_AXIMM_123_AWBURST,
    input wire [1:0]                      AP_AXIMM_123_AWLOCK,
    input wire [3:0]                      AP_AXIMM_123_AWCACHE,
    input wire [2:0]                      AP_AXIMM_123_AWPROT,
    input wire [3:0]                      AP_AXIMM_123_AWREGION,
    input wire [3:0]                      AP_AXIMM_123_AWQOS,
    input wire                            AP_AXIMM_123_AWVALID,
    output  wire                            AP_AXIMM_123_AWREADY,
    input wire [M_AXIMM_123_DATA_WIDTH-1:0]   AP_AXIMM_123_WDATA,
    input wire [M_AXIMM_123_DATA_WIDTH/8-1:0] AP_AXIMM_123_WSTRB,
    input wire                            AP_AXIMM_123_WLAST,
    input wire                            AP_AXIMM_123_WVALID,
    output  wire                            AP_AXIMM_123_WREADY,
    output  wire [1:0]                      AP_AXIMM_123_BRESP,
    output  wire                            AP_AXIMM_123_BVALID,
    input wire                            AP_AXIMM_123_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_123_ARADDR,
    input wire [7:0]                      AP_AXIMM_123_ARLEN,
    input wire [2:0]                      AP_AXIMM_123_ARSIZE,
    input wire [1:0]                      AP_AXIMM_123_ARBURST,
    input wire [1:0]                      AP_AXIMM_123_ARLOCK,
    input wire [3:0]                      AP_AXIMM_123_ARCACHE,
    input wire [2:0]                      AP_AXIMM_123_ARPROT,
    input wire [3:0]                      AP_AXIMM_123_ARREGION,
    input wire [3:0]                      AP_AXIMM_123_ARQOS,
    input wire                            AP_AXIMM_123_ARVALID,
    output  wire                            AP_AXIMM_123_ARREADY,
    output  wire [M_AXIMM_123_DATA_WIDTH-1:0]   AP_AXIMM_123_RDATA,
    output  wire [1:0]                      AP_AXIMM_123_RRESP,
    output  wire                            AP_AXIMM_123_RLAST,
    output  wire                            AP_AXIMM_123_RVALID,
    input  wire                            AP_AXIMM_123_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_123_AWADDR,
    output wire [7:0]                      M_AXIMM_123_AWLEN,
    output wire [2:0]                      M_AXIMM_123_AWSIZE,
    output wire [1:0]                      M_AXIMM_123_AWBURST,
    output wire [1:0]                      M_AXIMM_123_AWLOCK,
    output wire [3:0]                      M_AXIMM_123_AWCACHE,
    output wire [2:0]                      M_AXIMM_123_AWPROT,
    output wire [3:0]                      M_AXIMM_123_AWREGION,
    output wire [3:0]                      M_AXIMM_123_AWQOS,
    output wire                            M_AXIMM_123_AWVALID,
    input  wire                            M_AXIMM_123_AWREADY,
    output wire [M_AXIMM_123_DATA_WIDTH-1:0]   M_AXIMM_123_WDATA,
    output wire [M_AXIMM_123_DATA_WIDTH/8-1:0] M_AXIMM_123_WSTRB,
    output wire                            M_AXIMM_123_WLAST,
    output wire                            M_AXIMM_123_WVALID,
    input  wire                            M_AXIMM_123_WREADY,
    input  wire [1:0]                      M_AXIMM_123_BRESP,
    input  wire                            M_AXIMM_123_BVALID,
    output wire                            M_AXIMM_123_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_123_ARADDR,
    output wire [7:0]                      M_AXIMM_123_ARLEN,
    output wire [2:0]                      M_AXIMM_123_ARSIZE,
    output wire [1:0]                      M_AXIMM_123_ARBURST,
    output wire [1:0]                      M_AXIMM_123_ARLOCK,
    output wire [3:0]                      M_AXIMM_123_ARCACHE,
    output wire [2:0]                      M_AXIMM_123_ARPROT,
    output wire [3:0]                      M_AXIMM_123_ARREGION,
    output wire [3:0]                      M_AXIMM_123_ARQOS,
    output wire                            M_AXIMM_123_ARVALID,
    input  wire                            M_AXIMM_123_ARREADY,
    input  wire [M_AXIMM_123_DATA_WIDTH-1:0]   M_AXIMM_123_RDATA,
    input  wire [1:0]                      M_AXIMM_123_RRESP,
    input  wire                            M_AXIMM_123_RLAST,
    input  wire                            M_AXIMM_123_RVALID,
    output wire                            M_AXIMM_123_RREADY,
    //AXI-MM pass-through interface 124
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_124_AWADDR,
    input wire [7:0]                      AP_AXIMM_124_AWLEN,
    input wire [2:0]                      AP_AXIMM_124_AWSIZE,
    input wire [1:0]                      AP_AXIMM_124_AWBURST,
    input wire [1:0]                      AP_AXIMM_124_AWLOCK,
    input wire [3:0]                      AP_AXIMM_124_AWCACHE,
    input wire [2:0]                      AP_AXIMM_124_AWPROT,
    input wire [3:0]                      AP_AXIMM_124_AWREGION,
    input wire [3:0]                      AP_AXIMM_124_AWQOS,
    input wire                            AP_AXIMM_124_AWVALID,
    output  wire                            AP_AXIMM_124_AWREADY,
    input wire [M_AXIMM_124_DATA_WIDTH-1:0]   AP_AXIMM_124_WDATA,
    input wire [M_AXIMM_124_DATA_WIDTH/8-1:0] AP_AXIMM_124_WSTRB,
    input wire                            AP_AXIMM_124_WLAST,
    input wire                            AP_AXIMM_124_WVALID,
    output  wire                            AP_AXIMM_124_WREADY,
    output  wire [1:0]                      AP_AXIMM_124_BRESP,
    output  wire                            AP_AXIMM_124_BVALID,
    input wire                            AP_AXIMM_124_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_124_ARADDR,
    input wire [7:0]                      AP_AXIMM_124_ARLEN,
    input wire [2:0]                      AP_AXIMM_124_ARSIZE,
    input wire [1:0]                      AP_AXIMM_124_ARBURST,
    input wire [1:0]                      AP_AXIMM_124_ARLOCK,
    input wire [3:0]                      AP_AXIMM_124_ARCACHE,
    input wire [2:0]                      AP_AXIMM_124_ARPROT,
    input wire [3:0]                      AP_AXIMM_124_ARREGION,
    input wire [3:0]                      AP_AXIMM_124_ARQOS,
    input wire                            AP_AXIMM_124_ARVALID,
    output  wire                            AP_AXIMM_124_ARREADY,
    output  wire [M_AXIMM_124_DATA_WIDTH-1:0]   AP_AXIMM_124_RDATA,
    output  wire [1:0]                      AP_AXIMM_124_RRESP,
    output  wire                            AP_AXIMM_124_RLAST,
    output  wire                            AP_AXIMM_124_RVALID,
    input  wire                            AP_AXIMM_124_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_124_AWADDR,
    output wire [7:0]                      M_AXIMM_124_AWLEN,
    output wire [2:0]                      M_AXIMM_124_AWSIZE,
    output wire [1:0]                      M_AXIMM_124_AWBURST,
    output wire [1:0]                      M_AXIMM_124_AWLOCK,
    output wire [3:0]                      M_AXIMM_124_AWCACHE,
    output wire [2:0]                      M_AXIMM_124_AWPROT,
    output wire [3:0]                      M_AXIMM_124_AWREGION,
    output wire [3:0]                      M_AXIMM_124_AWQOS,
    output wire                            M_AXIMM_124_AWVALID,
    input  wire                            M_AXIMM_124_AWREADY,
    output wire [M_AXIMM_124_DATA_WIDTH-1:0]   M_AXIMM_124_WDATA,
    output wire [M_AXIMM_124_DATA_WIDTH/8-1:0] M_AXIMM_124_WSTRB,
    output wire                            M_AXIMM_124_WLAST,
    output wire                            M_AXIMM_124_WVALID,
    input  wire                            M_AXIMM_124_WREADY,
    input  wire [1:0]                      M_AXIMM_124_BRESP,
    input  wire                            M_AXIMM_124_BVALID,
    output wire                            M_AXIMM_124_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_124_ARADDR,
    output wire [7:0]                      M_AXIMM_124_ARLEN,
    output wire [2:0]                      M_AXIMM_124_ARSIZE,
    output wire [1:0]                      M_AXIMM_124_ARBURST,
    output wire [1:0]                      M_AXIMM_124_ARLOCK,
    output wire [3:0]                      M_AXIMM_124_ARCACHE,
    output wire [2:0]                      M_AXIMM_124_ARPROT,
    output wire [3:0]                      M_AXIMM_124_ARREGION,
    output wire [3:0]                      M_AXIMM_124_ARQOS,
    output wire                            M_AXIMM_124_ARVALID,
    input  wire                            M_AXIMM_124_ARREADY,
    input  wire [M_AXIMM_124_DATA_WIDTH-1:0]   M_AXIMM_124_RDATA,
    input  wire [1:0]                      M_AXIMM_124_RRESP,
    input  wire                            M_AXIMM_124_RLAST,
    input  wire                            M_AXIMM_124_RVALID,
    output wire                            M_AXIMM_124_RREADY,
    //AXI-MM pass-through interface 125
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_125_AWADDR,
    input wire [7:0]                      AP_AXIMM_125_AWLEN,
    input wire [2:0]                      AP_AXIMM_125_AWSIZE,
    input wire [1:0]                      AP_AXIMM_125_AWBURST,
    input wire [1:0]                      AP_AXIMM_125_AWLOCK,
    input wire [3:0]                      AP_AXIMM_125_AWCACHE,
    input wire [2:0]                      AP_AXIMM_125_AWPROT,
    input wire [3:0]                      AP_AXIMM_125_AWREGION,
    input wire [3:0]                      AP_AXIMM_125_AWQOS,
    input wire                            AP_AXIMM_125_AWVALID,
    output  wire                            AP_AXIMM_125_AWREADY,
    input wire [M_AXIMM_125_DATA_WIDTH-1:0]   AP_AXIMM_125_WDATA,
    input wire [M_AXIMM_125_DATA_WIDTH/8-1:0] AP_AXIMM_125_WSTRB,
    input wire                            AP_AXIMM_125_WLAST,
    input wire                            AP_AXIMM_125_WVALID,
    output  wire                            AP_AXIMM_125_WREADY,
    output  wire [1:0]                      AP_AXIMM_125_BRESP,
    output  wire                            AP_AXIMM_125_BVALID,
    input wire                            AP_AXIMM_125_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_125_ARADDR,
    input wire [7:0]                      AP_AXIMM_125_ARLEN,
    input wire [2:0]                      AP_AXIMM_125_ARSIZE,
    input wire [1:0]                      AP_AXIMM_125_ARBURST,
    input wire [1:0]                      AP_AXIMM_125_ARLOCK,
    input wire [3:0]                      AP_AXIMM_125_ARCACHE,
    input wire [2:0]                      AP_AXIMM_125_ARPROT,
    input wire [3:0]                      AP_AXIMM_125_ARREGION,
    input wire [3:0]                      AP_AXIMM_125_ARQOS,
    input wire                            AP_AXIMM_125_ARVALID,
    output  wire                            AP_AXIMM_125_ARREADY,
    output  wire [M_AXIMM_125_DATA_WIDTH-1:0]   AP_AXIMM_125_RDATA,
    output  wire [1:0]                      AP_AXIMM_125_RRESP,
    output  wire                            AP_AXIMM_125_RLAST,
    output  wire                            AP_AXIMM_125_RVALID,
    input  wire                            AP_AXIMM_125_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_125_AWADDR,
    output wire [7:0]                      M_AXIMM_125_AWLEN,
    output wire [2:0]                      M_AXIMM_125_AWSIZE,
    output wire [1:0]                      M_AXIMM_125_AWBURST,
    output wire [1:0]                      M_AXIMM_125_AWLOCK,
    output wire [3:0]                      M_AXIMM_125_AWCACHE,
    output wire [2:0]                      M_AXIMM_125_AWPROT,
    output wire [3:0]                      M_AXIMM_125_AWREGION,
    output wire [3:0]                      M_AXIMM_125_AWQOS,
    output wire                            M_AXIMM_125_AWVALID,
    input  wire                            M_AXIMM_125_AWREADY,
    output wire [M_AXIMM_125_DATA_WIDTH-1:0]   M_AXIMM_125_WDATA,
    output wire [M_AXIMM_125_DATA_WIDTH/8-1:0] M_AXIMM_125_WSTRB,
    output wire                            M_AXIMM_125_WLAST,
    output wire                            M_AXIMM_125_WVALID,
    input  wire                            M_AXIMM_125_WREADY,
    input  wire [1:0]                      M_AXIMM_125_BRESP,
    input  wire                            M_AXIMM_125_BVALID,
    output wire                            M_AXIMM_125_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_125_ARADDR,
    output wire [7:0]                      M_AXIMM_125_ARLEN,
    output wire [2:0]                      M_AXIMM_125_ARSIZE,
    output wire [1:0]                      M_AXIMM_125_ARBURST,
    output wire [1:0]                      M_AXIMM_125_ARLOCK,
    output wire [3:0]                      M_AXIMM_125_ARCACHE,
    output wire [2:0]                      M_AXIMM_125_ARPROT,
    output wire [3:0]                      M_AXIMM_125_ARREGION,
    output wire [3:0]                      M_AXIMM_125_ARQOS,
    output wire                            M_AXIMM_125_ARVALID,
    input  wire                            M_AXIMM_125_ARREADY,
    input  wire [M_AXIMM_125_DATA_WIDTH-1:0]   M_AXIMM_125_RDATA,
    input  wire [1:0]                      M_AXIMM_125_RRESP,
    input  wire                            M_AXIMM_125_RLAST,
    input  wire                            M_AXIMM_125_RVALID,
    output wire                            M_AXIMM_125_RREADY,
    //AXI-MM pass-through interface 126
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_126_AWADDR,
    input wire [7:0]                      AP_AXIMM_126_AWLEN,
    input wire [2:0]                      AP_AXIMM_126_AWSIZE,
    input wire [1:0]                      AP_AXIMM_126_AWBURST,
    input wire [1:0]                      AP_AXIMM_126_AWLOCK,
    input wire [3:0]                      AP_AXIMM_126_AWCACHE,
    input wire [2:0]                      AP_AXIMM_126_AWPROT,
    input wire [3:0]                      AP_AXIMM_126_AWREGION,
    input wire [3:0]                      AP_AXIMM_126_AWQOS,
    input wire                            AP_AXIMM_126_AWVALID,
    output  wire                            AP_AXIMM_126_AWREADY,
    input wire [M_AXIMM_126_DATA_WIDTH-1:0]   AP_AXIMM_126_WDATA,
    input wire [M_AXIMM_126_DATA_WIDTH/8-1:0] AP_AXIMM_126_WSTRB,
    input wire                            AP_AXIMM_126_WLAST,
    input wire                            AP_AXIMM_126_WVALID,
    output  wire                            AP_AXIMM_126_WREADY,
    output  wire [1:0]                      AP_AXIMM_126_BRESP,
    output  wire                            AP_AXIMM_126_BVALID,
    input wire                            AP_AXIMM_126_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_126_ARADDR,
    input wire [7:0]                      AP_AXIMM_126_ARLEN,
    input wire [2:0]                      AP_AXIMM_126_ARSIZE,
    input wire [1:0]                      AP_AXIMM_126_ARBURST,
    input wire [1:0]                      AP_AXIMM_126_ARLOCK,
    input wire [3:0]                      AP_AXIMM_126_ARCACHE,
    input wire [2:0]                      AP_AXIMM_126_ARPROT,
    input wire [3:0]                      AP_AXIMM_126_ARREGION,
    input wire [3:0]                      AP_AXIMM_126_ARQOS,
    input wire                            AP_AXIMM_126_ARVALID,
    output  wire                            AP_AXIMM_126_ARREADY,
    output  wire [M_AXIMM_126_DATA_WIDTH-1:0]   AP_AXIMM_126_RDATA,
    output  wire [1:0]                      AP_AXIMM_126_RRESP,
    output  wire                            AP_AXIMM_126_RLAST,
    output  wire                            AP_AXIMM_126_RVALID,
    input  wire                            AP_AXIMM_126_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_126_AWADDR,
    output wire [7:0]                      M_AXIMM_126_AWLEN,
    output wire [2:0]                      M_AXIMM_126_AWSIZE,
    output wire [1:0]                      M_AXIMM_126_AWBURST,
    output wire [1:0]                      M_AXIMM_126_AWLOCK,
    output wire [3:0]                      M_AXIMM_126_AWCACHE,
    output wire [2:0]                      M_AXIMM_126_AWPROT,
    output wire [3:0]                      M_AXIMM_126_AWREGION,
    output wire [3:0]                      M_AXIMM_126_AWQOS,
    output wire                            M_AXIMM_126_AWVALID,
    input  wire                            M_AXIMM_126_AWREADY,
    output wire [M_AXIMM_126_DATA_WIDTH-1:0]   M_AXIMM_126_WDATA,
    output wire [M_AXIMM_126_DATA_WIDTH/8-1:0] M_AXIMM_126_WSTRB,
    output wire                            M_AXIMM_126_WLAST,
    output wire                            M_AXIMM_126_WVALID,
    input  wire                            M_AXIMM_126_WREADY,
    input  wire [1:0]                      M_AXIMM_126_BRESP,
    input  wire                            M_AXIMM_126_BVALID,
    output wire                            M_AXIMM_126_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_126_ARADDR,
    output wire [7:0]                      M_AXIMM_126_ARLEN,
    output wire [2:0]                      M_AXIMM_126_ARSIZE,
    output wire [1:0]                      M_AXIMM_126_ARBURST,
    output wire [1:0]                      M_AXIMM_126_ARLOCK,
    output wire [3:0]                      M_AXIMM_126_ARCACHE,
    output wire [2:0]                      M_AXIMM_126_ARPROT,
    output wire [3:0]                      M_AXIMM_126_ARREGION,
    output wire [3:0]                      M_AXIMM_126_ARQOS,
    output wire                            M_AXIMM_126_ARVALID,
    input  wire                            M_AXIMM_126_ARREADY,
    input  wire [M_AXIMM_126_DATA_WIDTH-1:0]   M_AXIMM_126_RDATA,
    input  wire [1:0]                      M_AXIMM_126_RRESP,
    input  wire                            M_AXIMM_126_RLAST,
    input  wire                            M_AXIMM_126_RVALID,
    output wire                            M_AXIMM_126_RREADY,
    //AXI-MM pass-through interface 127
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_127_AWADDR,
    input wire [7:0]                      AP_AXIMM_127_AWLEN,
    input wire [2:0]                      AP_AXIMM_127_AWSIZE,
    input wire [1:0]                      AP_AXIMM_127_AWBURST,
    input wire [1:0]                      AP_AXIMM_127_AWLOCK,
    input wire [3:0]                      AP_AXIMM_127_AWCACHE,
    input wire [2:0]                      AP_AXIMM_127_AWPROT,
    input wire [3:0]                      AP_AXIMM_127_AWREGION,
    input wire [3:0]                      AP_AXIMM_127_AWQOS,
    input wire                            AP_AXIMM_127_AWVALID,
    output  wire                            AP_AXIMM_127_AWREADY,
    input wire [M_AXIMM_127_DATA_WIDTH-1:0]   AP_AXIMM_127_WDATA,
    input wire [M_AXIMM_127_DATA_WIDTH/8-1:0] AP_AXIMM_127_WSTRB,
    input wire                            AP_AXIMM_127_WLAST,
    input wire                            AP_AXIMM_127_WVALID,
    output  wire                            AP_AXIMM_127_WREADY,
    output  wire [1:0]                      AP_AXIMM_127_BRESP,
    output  wire                            AP_AXIMM_127_BVALID,
    input wire                            AP_AXIMM_127_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_127_ARADDR,
    input wire [7:0]                      AP_AXIMM_127_ARLEN,
    input wire [2:0]                      AP_AXIMM_127_ARSIZE,
    input wire [1:0]                      AP_AXIMM_127_ARBURST,
    input wire [1:0]                      AP_AXIMM_127_ARLOCK,
    input wire [3:0]                      AP_AXIMM_127_ARCACHE,
    input wire [2:0]                      AP_AXIMM_127_ARPROT,
    input wire [3:0]                      AP_AXIMM_127_ARREGION,
    input wire [3:0]                      AP_AXIMM_127_ARQOS,
    input wire                            AP_AXIMM_127_ARVALID,
    output  wire                            AP_AXIMM_127_ARREADY,
    output  wire [M_AXIMM_127_DATA_WIDTH-1:0]   AP_AXIMM_127_RDATA,
    output  wire [1:0]                      AP_AXIMM_127_RRESP,
    output  wire                            AP_AXIMM_127_RLAST,
    output  wire                            AP_AXIMM_127_RVALID,
    input  wire                            AP_AXIMM_127_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_127_AWADDR,
    output wire [7:0]                      M_AXIMM_127_AWLEN,
    output wire [2:0]                      M_AXIMM_127_AWSIZE,
    output wire [1:0]                      M_AXIMM_127_AWBURST,
    output wire [1:0]                      M_AXIMM_127_AWLOCK,
    output wire [3:0]                      M_AXIMM_127_AWCACHE,
    output wire [2:0]                      M_AXIMM_127_AWPROT,
    output wire [3:0]                      M_AXIMM_127_AWREGION,
    output wire [3:0]                      M_AXIMM_127_AWQOS,
    output wire                            M_AXIMM_127_AWVALID,
    input  wire                            M_AXIMM_127_AWREADY,
    output wire [M_AXIMM_127_DATA_WIDTH-1:0]   M_AXIMM_127_WDATA,
    output wire [M_AXIMM_127_DATA_WIDTH/8-1:0] M_AXIMM_127_WSTRB,
    output wire                            M_AXIMM_127_WLAST,
    output wire                            M_AXIMM_127_WVALID,
    input  wire                            M_AXIMM_127_WREADY,
    input  wire [1:0]                      M_AXIMM_127_BRESP,
    input  wire                            M_AXIMM_127_BVALID,
    output wire                            M_AXIMM_127_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_127_ARADDR,
    output wire [7:0]                      M_AXIMM_127_ARLEN,
    output wire [2:0]                      M_AXIMM_127_ARSIZE,
    output wire [1:0]                      M_AXIMM_127_ARBURST,
    output wire [1:0]                      M_AXIMM_127_ARLOCK,
    output wire [3:0]                      M_AXIMM_127_ARCACHE,
    output wire [2:0]                      M_AXIMM_127_ARPROT,
    output wire [3:0]                      M_AXIMM_127_ARREGION,
    output wire [3:0]                      M_AXIMM_127_ARQOS,
    output wire                            M_AXIMM_127_ARVALID,
    input  wire                            M_AXIMM_127_ARREADY,
    input  wire [M_AXIMM_127_DATA_WIDTH-1:0]   M_AXIMM_127_RDATA,
    input  wire [1:0]                      M_AXIMM_127_RRESP,
    input  wire                            M_AXIMM_127_RLAST,
    input  wire                            M_AXIMM_127_RVALID,
    output wire                            M_AXIMM_127_RREADY,
    output wire                                ap_done_irq
);



    //scalar interface 
    wire [31:0] scalar_write_addr;
    wire [31:0] scalar_read_addr;
    wire [31:0] scalar_din;
    wire scalar_we;
    wire scalar_re;
    wire [31:0] scalar_dout;
    wire [C_N_INPUT_SCALARS-1:0] inscalar_next;
    wire [C_N_INPUT_SCALARS-1:0] inscalar_fifo_empty;
    wire [C_N_INPUT_SCALARS-1:0] inscalar_fifo_full;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_fifo_empty;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_fifo_full;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_null_empty;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_null_dout;
    wire [C_N_OUTPUT_SCALARS-1:0] outscalar_null_read;
    
    //wire in bram control interface
    wire inbram_ctrl_allow;
    wire [C_NUM_INPUT_BRAMs-1:0] inbram_ctrl_ready;
    wire [C_NUM_INPUT_BRAMs-1:0] inoutbram_ctrl_ready;
    wire [C_NUM_INPUT_BRAMs*32-1:0] inbram_depth;
    
    //wire in fifo control interface
    wire infifo_ctrl_allow;
    
    //wire out bram control interface
    wire outbram_ctrl_allow;
    wire [C_NUM_OUTPUT_BRAMs-1:0] outbram_ctrl_ready;
    wire [C_NUM_OUTPUT_BRAMs-1:0] outbram_ctrl_canstart;
    wire [C_NUM_OUTPUT_BRAMs*32-1:0] outbram_depth;
    wire [C_NUM_OUTPUT_BRAMs-1:0] outbram_depth_write;
    
    //wire out fifo control interface
    wire outfifo_ctrl_allow;

    //wire in axis control interface
    wire inaxis_ctrl_allow;
    //wire out axis control interface
    wire outaxis_ctrl_allow;

    adapter #(
        .C_ACC_RESET_POLARITY(C_ACC_RESET_POLARITY),
        .C_NUM_INPUT_SCALARS(C_N_INPUT_SCALARS),
        .C_NUM_OUTPUT_SCALARS(C_N_OUTPUT_SCALARS),
        .C_QUEUE_DEPTH(C_QUEUE_DEPTH),
        .C_NUM_INPUT_FIFOs(C_NUM_INPUT_FIFOs),
        .C_NUM_OUTPUT_FIFOs(C_NUM_OUTPUT_FIFOs),
        .C_NUM_INPUT_BRAMs(C_NUM_INPUT_BRAMs),
        .C_NUM_OUTPUT_BRAMs(C_NUM_OUTPUT_BRAMs)
    ) adapter_i (
        .S_AXI_ACLK(s_axi_aclk),
        .S_AXI_ARESETN(s_axi_aresetn),
        .S_AXI_AWADDR(S_AXI_AWADDR),
        .S_AXI_AWPROT(S_AXI_AWPROT),
        .S_AXI_AWVALID(S_AXI_AWVALID),
        .S_AXI_AWREADY(S_AXI_AWREADY),
        .S_AXI_WDATA(S_AXI_WDATA),
        .S_AXI_WSTRB(S_AXI_WSTRB),
        .S_AXI_WVALID(S_AXI_WVALID),
        .S_AXI_WREADY(S_AXI_WREADY),
        .S_AXI_BRESP(S_AXI_BRESP),
        .S_AXI_BVALID(S_AXI_BVALID),
        .S_AXI_BREADY(S_AXI_BREADY),
        .S_AXI_ARADDR(S_AXI_ARADDR),
        .S_AXI_ARPROT(S_AXI_ARPROT),
        .S_AXI_ARVALID(S_AXI_ARVALID),
        .S_AXI_ARREADY(S_AXI_ARREADY),
        .S_AXI_RDATA(S_AXI_RDATA),
        .S_AXI_RRESP(S_AXI_RRESP),
        .S_AXI_RVALID(S_AXI_RVALID),
        .S_AXI_RREADY(S_AXI_RREADY),
        .acc_clk(acc_aclk),
        .acc_rstn(acc_aresetn),
        .ap_rst(ap_resetn),
        .ap_start(ap_start),
        .ap_start_single(ap_start_single),
        .ap_idle(ap_idle),
        .ap_done(ap_done),
        .ap_ready(ap_ready),
        .ap_continue(ap_continue),
        .ap_clk(ap_clk),
        .scalar_write_addr(scalar_write_addr),
        .scalar_read_addr(scalar_read_addr),
        .scalar_din(scalar_din),
        .scalar_we(scalar_we),
        .scalar_re(scalar_re),
        .scalar_dout(scalar_dout),
        .inscalar_next(inscalar_next),
        .inscalar_fifo_empty(inscalar_fifo_empty),
        .inscalar_fifo_full(inscalar_fifo_full),
        .outscalar_fifo_empty(outscalar_fifo_empty),
        .outscalar_fifo_full(outscalar_fifo_full),
        .outscalar_null_empty(outscalar_null_empty),
        .outscalar_null_dout(outscalar_null_dout),
        .outscalar_null_read(outscalar_null_read),
        .inbram_ctrl_allow(inbram_ctrl_allow),
        .inbram_ctrl_ready(inbram_ctrl_ready),
        .inoutbram_ctrl_ready(inoutbram_ctrl_ready),
        .infifo_ctrl_allow(infifo_ctrl_allow),
        .outbram_ctrl_allow(outbram_ctrl_allow),
        .outbram_ctrl_ready(outbram_ctrl_ready),
        .outbram_ctrl_canstart(outbram_ctrl_canstart),
        .outbram_depth(outbram_depth),
        .outbram_depth_write(outbram_depth_write),
        .outfifo_ctrl_allow(outfifo_ctrl_allow),
        .inaxis_ctrl_allow(inaxis_ctrl_allow),
        .outaxis_ctrl_allow(outaxis_ctrl_allow),
        .ap_done_irq(ap_done_irq)
    );
    
    scalar #(
        .C_NUM_INSCALARS(C_N_INPUT_SCALARS),
        .C_NUM_OUTSCALARS(C_N_OUTPUT_SCALARS),
        .C_FIFO_DEPTH(C_FIFO_DEPTH),
        .C_HAS_RETURN(C_HAS_RETURN),
        .C_INSCALAR_0_BITS(C_INPUT_SCALAR_0_WIDTH),
        .C_INSCALAR_1_BITS(C_INPUT_SCALAR_1_WIDTH),
        .C_INSCALAR_2_BITS(C_INPUT_SCALAR_2_WIDTH),
        .C_INSCALAR_3_BITS(C_INPUT_SCALAR_3_WIDTH),
        .C_INSCALAR_4_BITS(C_INPUT_SCALAR_4_WIDTH),
        .C_INSCALAR_5_BITS(C_INPUT_SCALAR_5_WIDTH),
        .C_INSCALAR_6_BITS(C_INPUT_SCALAR_6_WIDTH),
        .C_INSCALAR_7_BITS(C_INPUT_SCALAR_7_WIDTH),
        .C_INSCALAR_8_BITS(C_INPUT_SCALAR_8_WIDTH),
        .C_INSCALAR_9_BITS(C_INPUT_SCALAR_9_WIDTH),
        .C_INSCALAR_10_BITS(C_INPUT_SCALAR_10_WIDTH),
        .C_INSCALAR_11_BITS(C_INPUT_SCALAR_11_WIDTH),
        .C_INSCALAR_12_BITS(C_INPUT_SCALAR_12_WIDTH),
        .C_INSCALAR_13_BITS(C_INPUT_SCALAR_13_WIDTH),
        .C_INSCALAR_14_BITS(C_INPUT_SCALAR_14_WIDTH),
        .C_INSCALAR_15_BITS(C_INPUT_SCALAR_15_WIDTH),
        .C_INSCALAR_16_BITS(C_INPUT_SCALAR_16_WIDTH),
        .C_INSCALAR_17_BITS(C_INPUT_SCALAR_17_WIDTH),
        .C_INSCALAR_18_BITS(C_INPUT_SCALAR_18_WIDTH),
        .C_INSCALAR_19_BITS(C_INPUT_SCALAR_19_WIDTH),
        .C_INSCALAR_20_BITS(C_INPUT_SCALAR_20_WIDTH),
        .C_INSCALAR_21_BITS(C_INPUT_SCALAR_21_WIDTH),
        .C_INSCALAR_22_BITS(C_INPUT_SCALAR_22_WIDTH),
        .C_INSCALAR_23_BITS(C_INPUT_SCALAR_23_WIDTH),
        .C_INSCALAR_24_BITS(C_INPUT_SCALAR_24_WIDTH),
        .C_INSCALAR_25_BITS(C_INPUT_SCALAR_25_WIDTH),
        .C_INSCALAR_26_BITS(C_INPUT_SCALAR_26_WIDTH),
        .C_INSCALAR_27_BITS(C_INPUT_SCALAR_27_WIDTH),
        .C_INSCALAR_28_BITS(C_INPUT_SCALAR_28_WIDTH),
        .C_INSCALAR_29_BITS(C_INPUT_SCALAR_29_WIDTH),
        .C_INSCALAR_30_BITS(C_INPUT_SCALAR_30_WIDTH),
        .C_INSCALAR_31_BITS(C_INPUT_SCALAR_31_WIDTH),
        .C_INSCALAR_32_BITS(C_INPUT_SCALAR_32_WIDTH),
        .C_INSCALAR_33_BITS(C_INPUT_SCALAR_33_WIDTH),
        .C_INSCALAR_34_BITS(C_INPUT_SCALAR_34_WIDTH),
        .C_INSCALAR_35_BITS(C_INPUT_SCALAR_35_WIDTH),
        .C_INSCALAR_36_BITS(C_INPUT_SCALAR_36_WIDTH),
        .C_INSCALAR_37_BITS(C_INPUT_SCALAR_37_WIDTH),
        .C_INSCALAR_38_BITS(C_INPUT_SCALAR_38_WIDTH),
        .C_INSCALAR_39_BITS(C_INPUT_SCALAR_39_WIDTH),
        .C_INSCALAR_40_BITS(C_INPUT_SCALAR_40_WIDTH),
        .C_INSCALAR_41_BITS(C_INPUT_SCALAR_41_WIDTH),
        .C_INSCALAR_42_BITS(C_INPUT_SCALAR_42_WIDTH),
        .C_INSCALAR_43_BITS(C_INPUT_SCALAR_43_WIDTH),
        .C_INSCALAR_44_BITS(C_INPUT_SCALAR_44_WIDTH),
        .C_INSCALAR_45_BITS(C_INPUT_SCALAR_45_WIDTH),
        .C_INSCALAR_46_BITS(C_INPUT_SCALAR_46_WIDTH),
        .C_INSCALAR_47_BITS(C_INPUT_SCALAR_47_WIDTH),
        .C_INSCALAR_48_BITS(C_INPUT_SCALAR_48_WIDTH),
        .C_INSCALAR_49_BITS(C_INPUT_SCALAR_49_WIDTH),
        .C_INSCALAR_50_BITS(C_INPUT_SCALAR_50_WIDTH),
        .C_INSCALAR_51_BITS(C_INPUT_SCALAR_51_WIDTH),
        .C_INSCALAR_52_BITS(C_INPUT_SCALAR_52_WIDTH),
        .C_INSCALAR_53_BITS(C_INPUT_SCALAR_53_WIDTH),
        .C_INSCALAR_54_BITS(C_INPUT_SCALAR_54_WIDTH),
        .C_INSCALAR_55_BITS(C_INPUT_SCALAR_55_WIDTH),
        .C_INSCALAR_56_BITS(C_INPUT_SCALAR_56_WIDTH),
        .C_INSCALAR_57_BITS(C_INPUT_SCALAR_57_WIDTH),
        .C_INSCALAR_58_BITS(C_INPUT_SCALAR_58_WIDTH),
        .C_INSCALAR_59_BITS(C_INPUT_SCALAR_59_WIDTH),
        .C_INSCALAR_60_BITS(C_INPUT_SCALAR_60_WIDTH),
        .C_INSCALAR_61_BITS(C_INPUT_SCALAR_61_WIDTH),
        .C_INSCALAR_62_BITS(C_INPUT_SCALAR_62_WIDTH),
        .C_INSCALAR_63_BITS(C_INPUT_SCALAR_63_WIDTH),
        .C_INSCALAR_64_BITS(C_INPUT_SCALAR_64_WIDTH),
        .C_INSCALAR_65_BITS(C_INPUT_SCALAR_65_WIDTH),
        .C_INSCALAR_66_BITS(C_INPUT_SCALAR_66_WIDTH),
        .C_INSCALAR_67_BITS(C_INPUT_SCALAR_67_WIDTH),
        .C_INSCALAR_68_BITS(C_INPUT_SCALAR_68_WIDTH),
        .C_INSCALAR_69_BITS(C_INPUT_SCALAR_69_WIDTH),
        .C_INSCALAR_70_BITS(C_INPUT_SCALAR_70_WIDTH),
        .C_INSCALAR_71_BITS(C_INPUT_SCALAR_71_WIDTH),
        .C_INSCALAR_72_BITS(C_INPUT_SCALAR_72_WIDTH),
        .C_INSCALAR_73_BITS(C_INPUT_SCALAR_73_WIDTH),
        .C_INSCALAR_74_BITS(C_INPUT_SCALAR_74_WIDTH),
        .C_INSCALAR_75_BITS(C_INPUT_SCALAR_75_WIDTH),
        .C_INSCALAR_76_BITS(C_INPUT_SCALAR_76_WIDTH),
        .C_INSCALAR_77_BITS(C_INPUT_SCALAR_77_WIDTH),
        .C_INSCALAR_78_BITS(C_INPUT_SCALAR_78_WIDTH),
        .C_INSCALAR_79_BITS(C_INPUT_SCALAR_79_WIDTH),
        .C_INSCALAR_80_BITS(C_INPUT_SCALAR_80_WIDTH),
        .C_INSCALAR_81_BITS(C_INPUT_SCALAR_81_WIDTH),
        .C_INSCALAR_82_BITS(C_INPUT_SCALAR_82_WIDTH),
        .C_INSCALAR_83_BITS(C_INPUT_SCALAR_83_WIDTH),
        .C_INSCALAR_84_BITS(C_INPUT_SCALAR_84_WIDTH),
        .C_INSCALAR_85_BITS(C_INPUT_SCALAR_85_WIDTH),
        .C_INSCALAR_86_BITS(C_INPUT_SCALAR_86_WIDTH),
        .C_INSCALAR_87_BITS(C_INPUT_SCALAR_87_WIDTH),
        .C_INSCALAR_88_BITS(C_INPUT_SCALAR_88_WIDTH),
        .C_INSCALAR_89_BITS(C_INPUT_SCALAR_89_WIDTH),
        .C_INSCALAR_90_BITS(C_INPUT_SCALAR_90_WIDTH),
        .C_INSCALAR_91_BITS(C_INPUT_SCALAR_91_WIDTH),
        .C_INSCALAR_92_BITS(C_INPUT_SCALAR_92_WIDTH),
        .C_INSCALAR_93_BITS(C_INPUT_SCALAR_93_WIDTH),
        .C_INSCALAR_94_BITS(C_INPUT_SCALAR_94_WIDTH),
        .C_INSCALAR_95_BITS(C_INPUT_SCALAR_95_WIDTH),
        .C_INSCALAR_96_BITS(C_INPUT_SCALAR_96_WIDTH),
        .C_INSCALAR_97_BITS(C_INPUT_SCALAR_97_WIDTH),
        .C_INSCALAR_98_BITS(C_INPUT_SCALAR_98_WIDTH),
        .C_INSCALAR_99_BITS(C_INPUT_SCALAR_99_WIDTH),
        .C_INSCALAR_100_BITS(C_INPUT_SCALAR_100_WIDTH),
        .C_INSCALAR_101_BITS(C_INPUT_SCALAR_101_WIDTH),
        .C_INSCALAR_102_BITS(C_INPUT_SCALAR_102_WIDTH),
        .C_INSCALAR_103_BITS(C_INPUT_SCALAR_103_WIDTH),
        .C_INSCALAR_104_BITS(C_INPUT_SCALAR_104_WIDTH),
        .C_INSCALAR_105_BITS(C_INPUT_SCALAR_105_WIDTH),
        .C_INSCALAR_106_BITS(C_INPUT_SCALAR_106_WIDTH),
        .C_INSCALAR_107_BITS(C_INPUT_SCALAR_107_WIDTH),
        .C_INSCALAR_108_BITS(C_INPUT_SCALAR_108_WIDTH),
        .C_INSCALAR_109_BITS(C_INPUT_SCALAR_109_WIDTH),
        .C_INSCALAR_110_BITS(C_INPUT_SCALAR_110_WIDTH),
        .C_INSCALAR_111_BITS(C_INPUT_SCALAR_111_WIDTH),
        .C_INSCALAR_112_BITS(C_INPUT_SCALAR_112_WIDTH),
        .C_INSCALAR_113_BITS(C_INPUT_SCALAR_113_WIDTH),
        .C_INSCALAR_114_BITS(C_INPUT_SCALAR_114_WIDTH),
        .C_INSCALAR_115_BITS(C_INPUT_SCALAR_115_WIDTH),
        .C_INSCALAR_116_BITS(C_INPUT_SCALAR_116_WIDTH),
        .C_INSCALAR_117_BITS(C_INPUT_SCALAR_117_WIDTH),
        .C_INSCALAR_118_BITS(C_INPUT_SCALAR_118_WIDTH),
        .C_INSCALAR_119_BITS(C_INPUT_SCALAR_119_WIDTH),
        .C_INSCALAR_120_BITS(C_INPUT_SCALAR_120_WIDTH),
        .C_INSCALAR_121_BITS(C_INPUT_SCALAR_121_WIDTH),
        .C_INSCALAR_122_BITS(C_INPUT_SCALAR_122_WIDTH),
        .C_INSCALAR_123_BITS(C_INPUT_SCALAR_123_WIDTH),
        .C_INSCALAR_124_BITS(C_INPUT_SCALAR_124_WIDTH),
        .C_INSCALAR_125_BITS(C_INPUT_SCALAR_125_WIDTH),
        .C_INSCALAR_126_BITS(C_INPUT_SCALAR_126_WIDTH),
        .C_INSCALAR_127_BITS(C_INPUT_SCALAR_127_WIDTH),
        .S_AXIS_SCALAR_0_IS_DIRECT(S_AXIS_SCALAR_0_IS_DIRECT),
        .S_AXIS_SCALAR_1_IS_DIRECT(S_AXIS_SCALAR_1_IS_DIRECT),
        .S_AXIS_SCALAR_2_IS_DIRECT(S_AXIS_SCALAR_2_IS_DIRECT),
        .S_AXIS_SCALAR_3_IS_DIRECT(S_AXIS_SCALAR_3_IS_DIRECT),
        .S_AXIS_SCALAR_4_IS_DIRECT(S_AXIS_SCALAR_4_IS_DIRECT),
        .S_AXIS_SCALAR_5_IS_DIRECT(S_AXIS_SCALAR_5_IS_DIRECT),
        .S_AXIS_SCALAR_6_IS_DIRECT(S_AXIS_SCALAR_6_IS_DIRECT),
        .S_AXIS_SCALAR_7_IS_DIRECT(S_AXIS_SCALAR_7_IS_DIRECT),
        .S_AXIS_SCALAR_8_IS_DIRECT(S_AXIS_SCALAR_8_IS_DIRECT),
        .S_AXIS_SCALAR_9_IS_DIRECT(S_AXIS_SCALAR_9_IS_DIRECT),
        .S_AXIS_SCALAR_10_IS_DIRECT(S_AXIS_SCALAR_10_IS_DIRECT),
        .S_AXIS_SCALAR_11_IS_DIRECT(S_AXIS_SCALAR_11_IS_DIRECT),
        .S_AXIS_SCALAR_12_IS_DIRECT(S_AXIS_SCALAR_12_IS_DIRECT),
        .S_AXIS_SCALAR_13_IS_DIRECT(S_AXIS_SCALAR_13_IS_DIRECT),
        .S_AXIS_SCALAR_14_IS_DIRECT(S_AXIS_SCALAR_14_IS_DIRECT),
        .S_AXIS_SCALAR_15_IS_DIRECT(S_AXIS_SCALAR_15_IS_DIRECT),
        .S_AXIS_SCALAR_16_IS_DIRECT(S_AXIS_SCALAR_16_IS_DIRECT),
        .S_AXIS_SCALAR_17_IS_DIRECT(S_AXIS_SCALAR_17_IS_DIRECT),
        .S_AXIS_SCALAR_18_IS_DIRECT(S_AXIS_SCALAR_18_IS_DIRECT),
        .S_AXIS_SCALAR_19_IS_DIRECT(S_AXIS_SCALAR_19_IS_DIRECT),
        .S_AXIS_SCALAR_20_IS_DIRECT(S_AXIS_SCALAR_20_IS_DIRECT),
        .S_AXIS_SCALAR_21_IS_DIRECT(S_AXIS_SCALAR_21_IS_DIRECT),
        .S_AXIS_SCALAR_22_IS_DIRECT(S_AXIS_SCALAR_22_IS_DIRECT),
        .S_AXIS_SCALAR_23_IS_DIRECT(S_AXIS_SCALAR_23_IS_DIRECT),
        .S_AXIS_SCALAR_24_IS_DIRECT(S_AXIS_SCALAR_24_IS_DIRECT),
        .S_AXIS_SCALAR_25_IS_DIRECT(S_AXIS_SCALAR_25_IS_DIRECT),
        .S_AXIS_SCALAR_26_IS_DIRECT(S_AXIS_SCALAR_26_IS_DIRECT),
        .S_AXIS_SCALAR_27_IS_DIRECT(S_AXIS_SCALAR_27_IS_DIRECT),
        .S_AXIS_SCALAR_28_IS_DIRECT(S_AXIS_SCALAR_28_IS_DIRECT),
        .S_AXIS_SCALAR_29_IS_DIRECT(S_AXIS_SCALAR_29_IS_DIRECT),
        .S_AXIS_SCALAR_30_IS_DIRECT(S_AXIS_SCALAR_30_IS_DIRECT),
        .S_AXIS_SCALAR_31_IS_DIRECT(S_AXIS_SCALAR_31_IS_DIRECT),
        .S_AXIS_SCALAR_32_IS_DIRECT(S_AXIS_SCALAR_32_IS_DIRECT),
        .S_AXIS_SCALAR_33_IS_DIRECT(S_AXIS_SCALAR_33_IS_DIRECT),
        .S_AXIS_SCALAR_34_IS_DIRECT(S_AXIS_SCALAR_34_IS_DIRECT),
        .S_AXIS_SCALAR_35_IS_DIRECT(S_AXIS_SCALAR_35_IS_DIRECT),
        .S_AXIS_SCALAR_36_IS_DIRECT(S_AXIS_SCALAR_36_IS_DIRECT),
        .S_AXIS_SCALAR_37_IS_DIRECT(S_AXIS_SCALAR_37_IS_DIRECT),
        .S_AXIS_SCALAR_38_IS_DIRECT(S_AXIS_SCALAR_38_IS_DIRECT),
        .S_AXIS_SCALAR_39_IS_DIRECT(S_AXIS_SCALAR_39_IS_DIRECT),
        .S_AXIS_SCALAR_40_IS_DIRECT(S_AXIS_SCALAR_40_IS_DIRECT),
        .S_AXIS_SCALAR_41_IS_DIRECT(S_AXIS_SCALAR_41_IS_DIRECT),
        .S_AXIS_SCALAR_42_IS_DIRECT(S_AXIS_SCALAR_42_IS_DIRECT),
        .S_AXIS_SCALAR_43_IS_DIRECT(S_AXIS_SCALAR_43_IS_DIRECT),
        .S_AXIS_SCALAR_44_IS_DIRECT(S_AXIS_SCALAR_44_IS_DIRECT),
        .S_AXIS_SCALAR_45_IS_DIRECT(S_AXIS_SCALAR_45_IS_DIRECT),
        .S_AXIS_SCALAR_46_IS_DIRECT(S_AXIS_SCALAR_46_IS_DIRECT),
        .S_AXIS_SCALAR_47_IS_DIRECT(S_AXIS_SCALAR_47_IS_DIRECT),
        .S_AXIS_SCALAR_48_IS_DIRECT(S_AXIS_SCALAR_48_IS_DIRECT),
        .S_AXIS_SCALAR_49_IS_DIRECT(S_AXIS_SCALAR_49_IS_DIRECT),
        .S_AXIS_SCALAR_50_IS_DIRECT(S_AXIS_SCALAR_50_IS_DIRECT),
        .S_AXIS_SCALAR_51_IS_DIRECT(S_AXIS_SCALAR_51_IS_DIRECT),
        .S_AXIS_SCALAR_52_IS_DIRECT(S_AXIS_SCALAR_52_IS_DIRECT),
        .S_AXIS_SCALAR_53_IS_DIRECT(S_AXIS_SCALAR_53_IS_DIRECT),
        .S_AXIS_SCALAR_54_IS_DIRECT(S_AXIS_SCALAR_54_IS_DIRECT),
        .S_AXIS_SCALAR_55_IS_DIRECT(S_AXIS_SCALAR_55_IS_DIRECT),
        .S_AXIS_SCALAR_56_IS_DIRECT(S_AXIS_SCALAR_56_IS_DIRECT),
        .S_AXIS_SCALAR_57_IS_DIRECT(S_AXIS_SCALAR_57_IS_DIRECT),
        .S_AXIS_SCALAR_58_IS_DIRECT(S_AXIS_SCALAR_58_IS_DIRECT),
        .S_AXIS_SCALAR_59_IS_DIRECT(S_AXIS_SCALAR_59_IS_DIRECT),
        .S_AXIS_SCALAR_60_IS_DIRECT(S_AXIS_SCALAR_60_IS_DIRECT),
        .S_AXIS_SCALAR_61_IS_DIRECT(S_AXIS_SCALAR_61_IS_DIRECT),
        .S_AXIS_SCALAR_62_IS_DIRECT(S_AXIS_SCALAR_62_IS_DIRECT),
        .S_AXIS_SCALAR_63_IS_DIRECT(S_AXIS_SCALAR_63_IS_DIRECT),
        .S_AXIS_SCALAR_64_IS_DIRECT(S_AXIS_SCALAR_64_IS_DIRECT),
        .S_AXIS_SCALAR_65_IS_DIRECT(S_AXIS_SCALAR_65_IS_DIRECT),
        .S_AXIS_SCALAR_66_IS_DIRECT(S_AXIS_SCALAR_66_IS_DIRECT),
        .S_AXIS_SCALAR_67_IS_DIRECT(S_AXIS_SCALAR_67_IS_DIRECT),
        .S_AXIS_SCALAR_68_IS_DIRECT(S_AXIS_SCALAR_68_IS_DIRECT),
        .S_AXIS_SCALAR_69_IS_DIRECT(S_AXIS_SCALAR_69_IS_DIRECT),
        .S_AXIS_SCALAR_70_IS_DIRECT(S_AXIS_SCALAR_70_IS_DIRECT),
        .S_AXIS_SCALAR_71_IS_DIRECT(S_AXIS_SCALAR_71_IS_DIRECT),
        .S_AXIS_SCALAR_72_IS_DIRECT(S_AXIS_SCALAR_72_IS_DIRECT),
        .S_AXIS_SCALAR_73_IS_DIRECT(S_AXIS_SCALAR_73_IS_DIRECT),
        .S_AXIS_SCALAR_74_IS_DIRECT(S_AXIS_SCALAR_74_IS_DIRECT),
        .S_AXIS_SCALAR_75_IS_DIRECT(S_AXIS_SCALAR_75_IS_DIRECT),
        .S_AXIS_SCALAR_76_IS_DIRECT(S_AXIS_SCALAR_76_IS_DIRECT),
        .S_AXIS_SCALAR_77_IS_DIRECT(S_AXIS_SCALAR_77_IS_DIRECT),
        .S_AXIS_SCALAR_78_IS_DIRECT(S_AXIS_SCALAR_78_IS_DIRECT),
        .S_AXIS_SCALAR_79_IS_DIRECT(S_AXIS_SCALAR_79_IS_DIRECT),
        .S_AXIS_SCALAR_80_IS_DIRECT(S_AXIS_SCALAR_80_IS_DIRECT),
        .S_AXIS_SCALAR_81_IS_DIRECT(S_AXIS_SCALAR_81_IS_DIRECT),
        .S_AXIS_SCALAR_82_IS_DIRECT(S_AXIS_SCALAR_82_IS_DIRECT),
        .S_AXIS_SCALAR_83_IS_DIRECT(S_AXIS_SCALAR_83_IS_DIRECT),
        .S_AXIS_SCALAR_84_IS_DIRECT(S_AXIS_SCALAR_84_IS_DIRECT),
        .S_AXIS_SCALAR_85_IS_DIRECT(S_AXIS_SCALAR_85_IS_DIRECT),
        .S_AXIS_SCALAR_86_IS_DIRECT(S_AXIS_SCALAR_86_IS_DIRECT),
        .S_AXIS_SCALAR_87_IS_DIRECT(S_AXIS_SCALAR_87_IS_DIRECT),
        .S_AXIS_SCALAR_88_IS_DIRECT(S_AXIS_SCALAR_88_IS_DIRECT),
        .S_AXIS_SCALAR_89_IS_DIRECT(S_AXIS_SCALAR_89_IS_DIRECT),
        .S_AXIS_SCALAR_90_IS_DIRECT(S_AXIS_SCALAR_90_IS_DIRECT),
        .S_AXIS_SCALAR_91_IS_DIRECT(S_AXIS_SCALAR_91_IS_DIRECT),
        .S_AXIS_SCALAR_92_IS_DIRECT(S_AXIS_SCALAR_92_IS_DIRECT),
        .S_AXIS_SCALAR_93_IS_DIRECT(S_AXIS_SCALAR_93_IS_DIRECT),
        .S_AXIS_SCALAR_94_IS_DIRECT(S_AXIS_SCALAR_94_IS_DIRECT),
        .S_AXIS_SCALAR_95_IS_DIRECT(S_AXIS_SCALAR_95_IS_DIRECT),
        .S_AXIS_SCALAR_96_IS_DIRECT(S_AXIS_SCALAR_96_IS_DIRECT),
        .S_AXIS_SCALAR_97_IS_DIRECT(S_AXIS_SCALAR_97_IS_DIRECT),
        .S_AXIS_SCALAR_98_IS_DIRECT(S_AXIS_SCALAR_98_IS_DIRECT),
        .S_AXIS_SCALAR_99_IS_DIRECT(S_AXIS_SCALAR_99_IS_DIRECT),
        .S_AXIS_SCALAR_100_IS_DIRECT(S_AXIS_SCALAR_100_IS_DIRECT),
        .S_AXIS_SCALAR_101_IS_DIRECT(S_AXIS_SCALAR_101_IS_DIRECT),
        .S_AXIS_SCALAR_102_IS_DIRECT(S_AXIS_SCALAR_102_IS_DIRECT),
        .S_AXIS_SCALAR_103_IS_DIRECT(S_AXIS_SCALAR_103_IS_DIRECT),
        .S_AXIS_SCALAR_104_IS_DIRECT(S_AXIS_SCALAR_104_IS_DIRECT),
        .S_AXIS_SCALAR_105_IS_DIRECT(S_AXIS_SCALAR_105_IS_DIRECT),
        .S_AXIS_SCALAR_106_IS_DIRECT(S_AXIS_SCALAR_106_IS_DIRECT),
        .S_AXIS_SCALAR_107_IS_DIRECT(S_AXIS_SCALAR_107_IS_DIRECT),
        .S_AXIS_SCALAR_108_IS_DIRECT(S_AXIS_SCALAR_108_IS_DIRECT),
        .S_AXIS_SCALAR_109_IS_DIRECT(S_AXIS_SCALAR_109_IS_DIRECT),
        .S_AXIS_SCALAR_110_IS_DIRECT(S_AXIS_SCALAR_110_IS_DIRECT),
        .S_AXIS_SCALAR_111_IS_DIRECT(S_AXIS_SCALAR_111_IS_DIRECT),
        .S_AXIS_SCALAR_112_IS_DIRECT(S_AXIS_SCALAR_112_IS_DIRECT),
        .S_AXIS_SCALAR_113_IS_DIRECT(S_AXIS_SCALAR_113_IS_DIRECT),
        .S_AXIS_SCALAR_114_IS_DIRECT(S_AXIS_SCALAR_114_IS_DIRECT),
        .S_AXIS_SCALAR_115_IS_DIRECT(S_AXIS_SCALAR_115_IS_DIRECT),
        .S_AXIS_SCALAR_116_IS_DIRECT(S_AXIS_SCALAR_116_IS_DIRECT),
        .S_AXIS_SCALAR_117_IS_DIRECT(S_AXIS_SCALAR_117_IS_DIRECT),
        .S_AXIS_SCALAR_118_IS_DIRECT(S_AXIS_SCALAR_118_IS_DIRECT),
        .S_AXIS_SCALAR_119_IS_DIRECT(S_AXIS_SCALAR_119_IS_DIRECT),
        .S_AXIS_SCALAR_120_IS_DIRECT(S_AXIS_SCALAR_120_IS_DIRECT),
        .S_AXIS_SCALAR_121_IS_DIRECT(S_AXIS_SCALAR_121_IS_DIRECT),
        .S_AXIS_SCALAR_122_IS_DIRECT(S_AXIS_SCALAR_122_IS_DIRECT),
        .S_AXIS_SCALAR_123_IS_DIRECT(S_AXIS_SCALAR_123_IS_DIRECT),
        .S_AXIS_SCALAR_124_IS_DIRECT(S_AXIS_SCALAR_124_IS_DIRECT),
        .S_AXIS_SCALAR_125_IS_DIRECT(S_AXIS_SCALAR_125_IS_DIRECT),
        .S_AXIS_SCALAR_126_IS_DIRECT(S_AXIS_SCALAR_126_IS_DIRECT),
        .S_AXIS_SCALAR_127_IS_DIRECT(S_AXIS_SCALAR_127_IS_DIRECT),
        .S_AXIS_SCALAR_0_DIRECT_DMWIDTH(S_AXIS_SCALAR_0_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_1_DIRECT_DMWIDTH(S_AXIS_SCALAR_1_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_2_DIRECT_DMWIDTH(S_AXIS_SCALAR_2_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_3_DIRECT_DMWIDTH(S_AXIS_SCALAR_3_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_4_DIRECT_DMWIDTH(S_AXIS_SCALAR_4_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_5_DIRECT_DMWIDTH(S_AXIS_SCALAR_5_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_6_DIRECT_DMWIDTH(S_AXIS_SCALAR_6_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_7_DIRECT_DMWIDTH(S_AXIS_SCALAR_7_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_8_DIRECT_DMWIDTH(S_AXIS_SCALAR_8_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_9_DIRECT_DMWIDTH(S_AXIS_SCALAR_9_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_10_DIRECT_DMWIDTH(S_AXIS_SCALAR_10_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_11_DIRECT_DMWIDTH(S_AXIS_SCALAR_11_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_12_DIRECT_DMWIDTH(S_AXIS_SCALAR_12_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_13_DIRECT_DMWIDTH(S_AXIS_SCALAR_13_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_14_DIRECT_DMWIDTH(S_AXIS_SCALAR_14_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_15_DIRECT_DMWIDTH(S_AXIS_SCALAR_15_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_16_DIRECT_DMWIDTH(S_AXIS_SCALAR_16_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_17_DIRECT_DMWIDTH(S_AXIS_SCALAR_17_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_18_DIRECT_DMWIDTH(S_AXIS_SCALAR_18_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_19_DIRECT_DMWIDTH(S_AXIS_SCALAR_19_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_20_DIRECT_DMWIDTH(S_AXIS_SCALAR_20_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_21_DIRECT_DMWIDTH(S_AXIS_SCALAR_21_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_22_DIRECT_DMWIDTH(S_AXIS_SCALAR_22_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_23_DIRECT_DMWIDTH(S_AXIS_SCALAR_23_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_24_DIRECT_DMWIDTH(S_AXIS_SCALAR_24_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_25_DIRECT_DMWIDTH(S_AXIS_SCALAR_25_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_26_DIRECT_DMWIDTH(S_AXIS_SCALAR_26_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_27_DIRECT_DMWIDTH(S_AXIS_SCALAR_27_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_28_DIRECT_DMWIDTH(S_AXIS_SCALAR_28_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_29_DIRECT_DMWIDTH(S_AXIS_SCALAR_29_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_30_DIRECT_DMWIDTH(S_AXIS_SCALAR_30_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_31_DIRECT_DMWIDTH(S_AXIS_SCALAR_31_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_32_DIRECT_DMWIDTH(S_AXIS_SCALAR_32_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_33_DIRECT_DMWIDTH(S_AXIS_SCALAR_33_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_34_DIRECT_DMWIDTH(S_AXIS_SCALAR_34_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_35_DIRECT_DMWIDTH(S_AXIS_SCALAR_35_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_36_DIRECT_DMWIDTH(S_AXIS_SCALAR_36_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_37_DIRECT_DMWIDTH(S_AXIS_SCALAR_37_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_38_DIRECT_DMWIDTH(S_AXIS_SCALAR_38_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_39_DIRECT_DMWIDTH(S_AXIS_SCALAR_39_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_40_DIRECT_DMWIDTH(S_AXIS_SCALAR_40_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_41_DIRECT_DMWIDTH(S_AXIS_SCALAR_41_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_42_DIRECT_DMWIDTH(S_AXIS_SCALAR_42_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_43_DIRECT_DMWIDTH(S_AXIS_SCALAR_43_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_44_DIRECT_DMWIDTH(S_AXIS_SCALAR_44_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_45_DIRECT_DMWIDTH(S_AXIS_SCALAR_45_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_46_DIRECT_DMWIDTH(S_AXIS_SCALAR_46_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_47_DIRECT_DMWIDTH(S_AXIS_SCALAR_47_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_48_DIRECT_DMWIDTH(S_AXIS_SCALAR_48_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_49_DIRECT_DMWIDTH(S_AXIS_SCALAR_49_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_50_DIRECT_DMWIDTH(S_AXIS_SCALAR_50_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_51_DIRECT_DMWIDTH(S_AXIS_SCALAR_51_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_52_DIRECT_DMWIDTH(S_AXIS_SCALAR_52_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_53_DIRECT_DMWIDTH(S_AXIS_SCALAR_53_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_54_DIRECT_DMWIDTH(S_AXIS_SCALAR_54_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_55_DIRECT_DMWIDTH(S_AXIS_SCALAR_55_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_56_DIRECT_DMWIDTH(S_AXIS_SCALAR_56_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_57_DIRECT_DMWIDTH(S_AXIS_SCALAR_57_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_58_DIRECT_DMWIDTH(S_AXIS_SCALAR_58_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_59_DIRECT_DMWIDTH(S_AXIS_SCALAR_59_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_60_DIRECT_DMWIDTH(S_AXIS_SCALAR_60_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_61_DIRECT_DMWIDTH(S_AXIS_SCALAR_61_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_62_DIRECT_DMWIDTH(S_AXIS_SCALAR_62_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_63_DIRECT_DMWIDTH(S_AXIS_SCALAR_63_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_64_DIRECT_DMWIDTH(S_AXIS_SCALAR_64_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_65_DIRECT_DMWIDTH(S_AXIS_SCALAR_65_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_66_DIRECT_DMWIDTH(S_AXIS_SCALAR_66_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_67_DIRECT_DMWIDTH(S_AXIS_SCALAR_67_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_68_DIRECT_DMWIDTH(S_AXIS_SCALAR_68_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_69_DIRECT_DMWIDTH(S_AXIS_SCALAR_69_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_70_DIRECT_DMWIDTH(S_AXIS_SCALAR_70_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_71_DIRECT_DMWIDTH(S_AXIS_SCALAR_71_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_72_DIRECT_DMWIDTH(S_AXIS_SCALAR_72_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_73_DIRECT_DMWIDTH(S_AXIS_SCALAR_73_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_74_DIRECT_DMWIDTH(S_AXIS_SCALAR_74_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_75_DIRECT_DMWIDTH(S_AXIS_SCALAR_75_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_76_DIRECT_DMWIDTH(S_AXIS_SCALAR_76_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_77_DIRECT_DMWIDTH(S_AXIS_SCALAR_77_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_78_DIRECT_DMWIDTH(S_AXIS_SCALAR_78_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_79_DIRECT_DMWIDTH(S_AXIS_SCALAR_79_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_80_DIRECT_DMWIDTH(S_AXIS_SCALAR_80_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_81_DIRECT_DMWIDTH(S_AXIS_SCALAR_81_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_82_DIRECT_DMWIDTH(S_AXIS_SCALAR_82_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_83_DIRECT_DMWIDTH(S_AXIS_SCALAR_83_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_84_DIRECT_DMWIDTH(S_AXIS_SCALAR_84_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_85_DIRECT_DMWIDTH(S_AXIS_SCALAR_85_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_86_DIRECT_DMWIDTH(S_AXIS_SCALAR_86_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_87_DIRECT_DMWIDTH(S_AXIS_SCALAR_87_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_88_DIRECT_DMWIDTH(S_AXIS_SCALAR_88_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_89_DIRECT_DMWIDTH(S_AXIS_SCALAR_89_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_90_DIRECT_DMWIDTH(S_AXIS_SCALAR_90_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_91_DIRECT_DMWIDTH(S_AXIS_SCALAR_91_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_92_DIRECT_DMWIDTH(S_AXIS_SCALAR_92_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_93_DIRECT_DMWIDTH(S_AXIS_SCALAR_93_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_94_DIRECT_DMWIDTH(S_AXIS_SCALAR_94_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_95_DIRECT_DMWIDTH(S_AXIS_SCALAR_95_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_96_DIRECT_DMWIDTH(S_AXIS_SCALAR_96_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_97_DIRECT_DMWIDTH(S_AXIS_SCALAR_97_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_98_DIRECT_DMWIDTH(S_AXIS_SCALAR_98_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_99_DIRECT_DMWIDTH(S_AXIS_SCALAR_99_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_100_DIRECT_DMWIDTH(S_AXIS_SCALAR_100_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_101_DIRECT_DMWIDTH(S_AXIS_SCALAR_101_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_102_DIRECT_DMWIDTH(S_AXIS_SCALAR_102_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_103_DIRECT_DMWIDTH(S_AXIS_SCALAR_103_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_104_DIRECT_DMWIDTH(S_AXIS_SCALAR_104_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_105_DIRECT_DMWIDTH(S_AXIS_SCALAR_105_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_106_DIRECT_DMWIDTH(S_AXIS_SCALAR_106_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_107_DIRECT_DMWIDTH(S_AXIS_SCALAR_107_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_108_DIRECT_DMWIDTH(S_AXIS_SCALAR_108_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_109_DIRECT_DMWIDTH(S_AXIS_SCALAR_109_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_110_DIRECT_DMWIDTH(S_AXIS_SCALAR_110_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_111_DIRECT_DMWIDTH(S_AXIS_SCALAR_111_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_112_DIRECT_DMWIDTH(S_AXIS_SCALAR_112_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_113_DIRECT_DMWIDTH(S_AXIS_SCALAR_113_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_114_DIRECT_DMWIDTH(S_AXIS_SCALAR_114_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_115_DIRECT_DMWIDTH(S_AXIS_SCALAR_115_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_116_DIRECT_DMWIDTH(S_AXIS_SCALAR_116_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_117_DIRECT_DMWIDTH(S_AXIS_SCALAR_117_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_118_DIRECT_DMWIDTH(S_AXIS_SCALAR_118_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_119_DIRECT_DMWIDTH(S_AXIS_SCALAR_119_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_120_DIRECT_DMWIDTH(S_AXIS_SCALAR_120_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_121_DIRECT_DMWIDTH(S_AXIS_SCALAR_121_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_122_DIRECT_DMWIDTH(S_AXIS_SCALAR_122_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_123_DIRECT_DMWIDTH(S_AXIS_SCALAR_123_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_124_DIRECT_DMWIDTH(S_AXIS_SCALAR_124_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_125_DIRECT_DMWIDTH(S_AXIS_SCALAR_125_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_126_DIRECT_DMWIDTH(S_AXIS_SCALAR_126_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_127_DIRECT_DMWIDTH(S_AXIS_SCALAR_127_DIRECT_DMWIDTH),
        .S_AXIS_SCALAR_0_DIRECT_IS_ASYNC(S_AXIS_SCALAR_0_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_1_DIRECT_IS_ASYNC(S_AXIS_SCALAR_1_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_2_DIRECT_IS_ASYNC(S_AXIS_SCALAR_2_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_3_DIRECT_IS_ASYNC(S_AXIS_SCALAR_3_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_4_DIRECT_IS_ASYNC(S_AXIS_SCALAR_4_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_5_DIRECT_IS_ASYNC(S_AXIS_SCALAR_5_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_6_DIRECT_IS_ASYNC(S_AXIS_SCALAR_6_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_7_DIRECT_IS_ASYNC(S_AXIS_SCALAR_7_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_8_DIRECT_IS_ASYNC(S_AXIS_SCALAR_8_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_9_DIRECT_IS_ASYNC(S_AXIS_SCALAR_9_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_10_DIRECT_IS_ASYNC(S_AXIS_SCALAR_10_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_11_DIRECT_IS_ASYNC(S_AXIS_SCALAR_11_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_12_DIRECT_IS_ASYNC(S_AXIS_SCALAR_12_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_13_DIRECT_IS_ASYNC(S_AXIS_SCALAR_13_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_14_DIRECT_IS_ASYNC(S_AXIS_SCALAR_14_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_15_DIRECT_IS_ASYNC(S_AXIS_SCALAR_15_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_16_DIRECT_IS_ASYNC(S_AXIS_SCALAR_16_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_17_DIRECT_IS_ASYNC(S_AXIS_SCALAR_17_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_18_DIRECT_IS_ASYNC(S_AXIS_SCALAR_18_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_19_DIRECT_IS_ASYNC(S_AXIS_SCALAR_19_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_20_DIRECT_IS_ASYNC(S_AXIS_SCALAR_20_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_21_DIRECT_IS_ASYNC(S_AXIS_SCALAR_21_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_22_DIRECT_IS_ASYNC(S_AXIS_SCALAR_22_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_23_DIRECT_IS_ASYNC(S_AXIS_SCALAR_23_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_24_DIRECT_IS_ASYNC(S_AXIS_SCALAR_24_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_25_DIRECT_IS_ASYNC(S_AXIS_SCALAR_25_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_26_DIRECT_IS_ASYNC(S_AXIS_SCALAR_26_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_27_DIRECT_IS_ASYNC(S_AXIS_SCALAR_27_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_28_DIRECT_IS_ASYNC(S_AXIS_SCALAR_28_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_29_DIRECT_IS_ASYNC(S_AXIS_SCALAR_29_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_30_DIRECT_IS_ASYNC(S_AXIS_SCALAR_30_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_31_DIRECT_IS_ASYNC(S_AXIS_SCALAR_31_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_32_DIRECT_IS_ASYNC(S_AXIS_SCALAR_32_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_33_DIRECT_IS_ASYNC(S_AXIS_SCALAR_33_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_34_DIRECT_IS_ASYNC(S_AXIS_SCALAR_34_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_35_DIRECT_IS_ASYNC(S_AXIS_SCALAR_35_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_36_DIRECT_IS_ASYNC(S_AXIS_SCALAR_36_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_37_DIRECT_IS_ASYNC(S_AXIS_SCALAR_37_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_38_DIRECT_IS_ASYNC(S_AXIS_SCALAR_38_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_39_DIRECT_IS_ASYNC(S_AXIS_SCALAR_39_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_40_DIRECT_IS_ASYNC(S_AXIS_SCALAR_40_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_41_DIRECT_IS_ASYNC(S_AXIS_SCALAR_41_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_42_DIRECT_IS_ASYNC(S_AXIS_SCALAR_42_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_43_DIRECT_IS_ASYNC(S_AXIS_SCALAR_43_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_44_DIRECT_IS_ASYNC(S_AXIS_SCALAR_44_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_45_DIRECT_IS_ASYNC(S_AXIS_SCALAR_45_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_46_DIRECT_IS_ASYNC(S_AXIS_SCALAR_46_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_47_DIRECT_IS_ASYNC(S_AXIS_SCALAR_47_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_48_DIRECT_IS_ASYNC(S_AXIS_SCALAR_48_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_49_DIRECT_IS_ASYNC(S_AXIS_SCALAR_49_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_50_DIRECT_IS_ASYNC(S_AXIS_SCALAR_50_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_51_DIRECT_IS_ASYNC(S_AXIS_SCALAR_51_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_52_DIRECT_IS_ASYNC(S_AXIS_SCALAR_52_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_53_DIRECT_IS_ASYNC(S_AXIS_SCALAR_53_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_54_DIRECT_IS_ASYNC(S_AXIS_SCALAR_54_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_55_DIRECT_IS_ASYNC(S_AXIS_SCALAR_55_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_56_DIRECT_IS_ASYNC(S_AXIS_SCALAR_56_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_57_DIRECT_IS_ASYNC(S_AXIS_SCALAR_57_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_58_DIRECT_IS_ASYNC(S_AXIS_SCALAR_58_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_59_DIRECT_IS_ASYNC(S_AXIS_SCALAR_59_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_60_DIRECT_IS_ASYNC(S_AXIS_SCALAR_60_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_61_DIRECT_IS_ASYNC(S_AXIS_SCALAR_61_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_62_DIRECT_IS_ASYNC(S_AXIS_SCALAR_62_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_63_DIRECT_IS_ASYNC(S_AXIS_SCALAR_63_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_64_DIRECT_IS_ASYNC(S_AXIS_SCALAR_64_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_65_DIRECT_IS_ASYNC(S_AXIS_SCALAR_65_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_66_DIRECT_IS_ASYNC(S_AXIS_SCALAR_66_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_67_DIRECT_IS_ASYNC(S_AXIS_SCALAR_67_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_68_DIRECT_IS_ASYNC(S_AXIS_SCALAR_68_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_69_DIRECT_IS_ASYNC(S_AXIS_SCALAR_69_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_70_DIRECT_IS_ASYNC(S_AXIS_SCALAR_70_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_71_DIRECT_IS_ASYNC(S_AXIS_SCALAR_71_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_72_DIRECT_IS_ASYNC(S_AXIS_SCALAR_72_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_73_DIRECT_IS_ASYNC(S_AXIS_SCALAR_73_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_74_DIRECT_IS_ASYNC(S_AXIS_SCALAR_74_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_75_DIRECT_IS_ASYNC(S_AXIS_SCALAR_75_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_76_DIRECT_IS_ASYNC(S_AXIS_SCALAR_76_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_77_DIRECT_IS_ASYNC(S_AXIS_SCALAR_77_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_78_DIRECT_IS_ASYNC(S_AXIS_SCALAR_78_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_79_DIRECT_IS_ASYNC(S_AXIS_SCALAR_79_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_80_DIRECT_IS_ASYNC(S_AXIS_SCALAR_80_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_81_DIRECT_IS_ASYNC(S_AXIS_SCALAR_81_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_82_DIRECT_IS_ASYNC(S_AXIS_SCALAR_82_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_83_DIRECT_IS_ASYNC(S_AXIS_SCALAR_83_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_84_DIRECT_IS_ASYNC(S_AXIS_SCALAR_84_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_85_DIRECT_IS_ASYNC(S_AXIS_SCALAR_85_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_86_DIRECT_IS_ASYNC(S_AXIS_SCALAR_86_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_87_DIRECT_IS_ASYNC(S_AXIS_SCALAR_87_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_88_DIRECT_IS_ASYNC(S_AXIS_SCALAR_88_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_89_DIRECT_IS_ASYNC(S_AXIS_SCALAR_89_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_90_DIRECT_IS_ASYNC(S_AXIS_SCALAR_90_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_91_DIRECT_IS_ASYNC(S_AXIS_SCALAR_91_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_92_DIRECT_IS_ASYNC(S_AXIS_SCALAR_92_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_93_DIRECT_IS_ASYNC(S_AXIS_SCALAR_93_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_94_DIRECT_IS_ASYNC(S_AXIS_SCALAR_94_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_95_DIRECT_IS_ASYNC(S_AXIS_SCALAR_95_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_96_DIRECT_IS_ASYNC(S_AXIS_SCALAR_96_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_97_DIRECT_IS_ASYNC(S_AXIS_SCALAR_97_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_98_DIRECT_IS_ASYNC(S_AXIS_SCALAR_98_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_99_DIRECT_IS_ASYNC(S_AXIS_SCALAR_99_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_100_DIRECT_IS_ASYNC(S_AXIS_SCALAR_100_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_101_DIRECT_IS_ASYNC(S_AXIS_SCALAR_101_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_102_DIRECT_IS_ASYNC(S_AXIS_SCALAR_102_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_103_DIRECT_IS_ASYNC(S_AXIS_SCALAR_103_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_104_DIRECT_IS_ASYNC(S_AXIS_SCALAR_104_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_105_DIRECT_IS_ASYNC(S_AXIS_SCALAR_105_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_106_DIRECT_IS_ASYNC(S_AXIS_SCALAR_106_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_107_DIRECT_IS_ASYNC(S_AXIS_SCALAR_107_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_108_DIRECT_IS_ASYNC(S_AXIS_SCALAR_108_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_109_DIRECT_IS_ASYNC(S_AXIS_SCALAR_109_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_110_DIRECT_IS_ASYNC(S_AXIS_SCALAR_110_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_111_DIRECT_IS_ASYNC(S_AXIS_SCALAR_111_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_112_DIRECT_IS_ASYNC(S_AXIS_SCALAR_112_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_113_DIRECT_IS_ASYNC(S_AXIS_SCALAR_113_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_114_DIRECT_IS_ASYNC(S_AXIS_SCALAR_114_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_115_DIRECT_IS_ASYNC(S_AXIS_SCALAR_115_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_116_DIRECT_IS_ASYNC(S_AXIS_SCALAR_116_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_117_DIRECT_IS_ASYNC(S_AXIS_SCALAR_117_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_118_DIRECT_IS_ASYNC(S_AXIS_SCALAR_118_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_119_DIRECT_IS_ASYNC(S_AXIS_SCALAR_119_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_120_DIRECT_IS_ASYNC(S_AXIS_SCALAR_120_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_121_DIRECT_IS_ASYNC(S_AXIS_SCALAR_121_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_122_DIRECT_IS_ASYNC(S_AXIS_SCALAR_122_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_123_DIRECT_IS_ASYNC(S_AXIS_SCALAR_123_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_124_DIRECT_IS_ASYNC(S_AXIS_SCALAR_124_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_125_DIRECT_IS_ASYNC(S_AXIS_SCALAR_125_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_126_DIRECT_IS_ASYNC(S_AXIS_SCALAR_126_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_127_DIRECT_IS_ASYNC(S_AXIS_SCALAR_127_DIRECT_IS_ASYNC),
        .S_AXIS_SCALAR_0_DIRECT_DEPTH(S_AXIS_SCALAR_0_DIRECT_DEPTH),
        .S_AXIS_SCALAR_1_DIRECT_DEPTH(S_AXIS_SCALAR_1_DIRECT_DEPTH),
        .S_AXIS_SCALAR_2_DIRECT_DEPTH(S_AXIS_SCALAR_2_DIRECT_DEPTH),
        .S_AXIS_SCALAR_3_DIRECT_DEPTH(S_AXIS_SCALAR_3_DIRECT_DEPTH),
        .S_AXIS_SCALAR_4_DIRECT_DEPTH(S_AXIS_SCALAR_4_DIRECT_DEPTH),
        .S_AXIS_SCALAR_5_DIRECT_DEPTH(S_AXIS_SCALAR_5_DIRECT_DEPTH),
        .S_AXIS_SCALAR_6_DIRECT_DEPTH(S_AXIS_SCALAR_6_DIRECT_DEPTH),
        .S_AXIS_SCALAR_7_DIRECT_DEPTH(S_AXIS_SCALAR_7_DIRECT_DEPTH),
        .S_AXIS_SCALAR_8_DIRECT_DEPTH(S_AXIS_SCALAR_8_DIRECT_DEPTH),
        .S_AXIS_SCALAR_9_DIRECT_DEPTH(S_AXIS_SCALAR_9_DIRECT_DEPTH),
        .S_AXIS_SCALAR_10_DIRECT_DEPTH(S_AXIS_SCALAR_10_DIRECT_DEPTH),
        .S_AXIS_SCALAR_11_DIRECT_DEPTH(S_AXIS_SCALAR_11_DIRECT_DEPTH),
        .S_AXIS_SCALAR_12_DIRECT_DEPTH(S_AXIS_SCALAR_12_DIRECT_DEPTH),
        .S_AXIS_SCALAR_13_DIRECT_DEPTH(S_AXIS_SCALAR_13_DIRECT_DEPTH),
        .S_AXIS_SCALAR_14_DIRECT_DEPTH(S_AXIS_SCALAR_14_DIRECT_DEPTH),
        .S_AXIS_SCALAR_15_DIRECT_DEPTH(S_AXIS_SCALAR_15_DIRECT_DEPTH),
        .S_AXIS_SCALAR_16_DIRECT_DEPTH(S_AXIS_SCALAR_16_DIRECT_DEPTH),
        .S_AXIS_SCALAR_17_DIRECT_DEPTH(S_AXIS_SCALAR_17_DIRECT_DEPTH),
        .S_AXIS_SCALAR_18_DIRECT_DEPTH(S_AXIS_SCALAR_18_DIRECT_DEPTH),
        .S_AXIS_SCALAR_19_DIRECT_DEPTH(S_AXIS_SCALAR_19_DIRECT_DEPTH),
        .S_AXIS_SCALAR_20_DIRECT_DEPTH(S_AXIS_SCALAR_20_DIRECT_DEPTH),
        .S_AXIS_SCALAR_21_DIRECT_DEPTH(S_AXIS_SCALAR_21_DIRECT_DEPTH),
        .S_AXIS_SCALAR_22_DIRECT_DEPTH(S_AXIS_SCALAR_22_DIRECT_DEPTH),
        .S_AXIS_SCALAR_23_DIRECT_DEPTH(S_AXIS_SCALAR_23_DIRECT_DEPTH),
        .S_AXIS_SCALAR_24_DIRECT_DEPTH(S_AXIS_SCALAR_24_DIRECT_DEPTH),
        .S_AXIS_SCALAR_25_DIRECT_DEPTH(S_AXIS_SCALAR_25_DIRECT_DEPTH),
        .S_AXIS_SCALAR_26_DIRECT_DEPTH(S_AXIS_SCALAR_26_DIRECT_DEPTH),
        .S_AXIS_SCALAR_27_DIRECT_DEPTH(S_AXIS_SCALAR_27_DIRECT_DEPTH),
        .S_AXIS_SCALAR_28_DIRECT_DEPTH(S_AXIS_SCALAR_28_DIRECT_DEPTH),
        .S_AXIS_SCALAR_29_DIRECT_DEPTH(S_AXIS_SCALAR_29_DIRECT_DEPTH),
        .S_AXIS_SCALAR_30_DIRECT_DEPTH(S_AXIS_SCALAR_30_DIRECT_DEPTH),
        .S_AXIS_SCALAR_31_DIRECT_DEPTH(S_AXIS_SCALAR_31_DIRECT_DEPTH),
        .S_AXIS_SCALAR_32_DIRECT_DEPTH(S_AXIS_SCALAR_32_DIRECT_DEPTH),
        .S_AXIS_SCALAR_33_DIRECT_DEPTH(S_AXIS_SCALAR_33_DIRECT_DEPTH),
        .S_AXIS_SCALAR_34_DIRECT_DEPTH(S_AXIS_SCALAR_34_DIRECT_DEPTH),
        .S_AXIS_SCALAR_35_DIRECT_DEPTH(S_AXIS_SCALAR_35_DIRECT_DEPTH),
        .S_AXIS_SCALAR_36_DIRECT_DEPTH(S_AXIS_SCALAR_36_DIRECT_DEPTH),
        .S_AXIS_SCALAR_37_DIRECT_DEPTH(S_AXIS_SCALAR_37_DIRECT_DEPTH),
        .S_AXIS_SCALAR_38_DIRECT_DEPTH(S_AXIS_SCALAR_38_DIRECT_DEPTH),
        .S_AXIS_SCALAR_39_DIRECT_DEPTH(S_AXIS_SCALAR_39_DIRECT_DEPTH),
        .S_AXIS_SCALAR_40_DIRECT_DEPTH(S_AXIS_SCALAR_40_DIRECT_DEPTH),
        .S_AXIS_SCALAR_41_DIRECT_DEPTH(S_AXIS_SCALAR_41_DIRECT_DEPTH),
        .S_AXIS_SCALAR_42_DIRECT_DEPTH(S_AXIS_SCALAR_42_DIRECT_DEPTH),
        .S_AXIS_SCALAR_43_DIRECT_DEPTH(S_AXIS_SCALAR_43_DIRECT_DEPTH),
        .S_AXIS_SCALAR_44_DIRECT_DEPTH(S_AXIS_SCALAR_44_DIRECT_DEPTH),
        .S_AXIS_SCALAR_45_DIRECT_DEPTH(S_AXIS_SCALAR_45_DIRECT_DEPTH),
        .S_AXIS_SCALAR_46_DIRECT_DEPTH(S_AXIS_SCALAR_46_DIRECT_DEPTH),
        .S_AXIS_SCALAR_47_DIRECT_DEPTH(S_AXIS_SCALAR_47_DIRECT_DEPTH),
        .S_AXIS_SCALAR_48_DIRECT_DEPTH(S_AXIS_SCALAR_48_DIRECT_DEPTH),
        .S_AXIS_SCALAR_49_DIRECT_DEPTH(S_AXIS_SCALAR_49_DIRECT_DEPTH),
        .S_AXIS_SCALAR_50_DIRECT_DEPTH(S_AXIS_SCALAR_50_DIRECT_DEPTH),
        .S_AXIS_SCALAR_51_DIRECT_DEPTH(S_AXIS_SCALAR_51_DIRECT_DEPTH),
        .S_AXIS_SCALAR_52_DIRECT_DEPTH(S_AXIS_SCALAR_52_DIRECT_DEPTH),
        .S_AXIS_SCALAR_53_DIRECT_DEPTH(S_AXIS_SCALAR_53_DIRECT_DEPTH),
        .S_AXIS_SCALAR_54_DIRECT_DEPTH(S_AXIS_SCALAR_54_DIRECT_DEPTH),
        .S_AXIS_SCALAR_55_DIRECT_DEPTH(S_AXIS_SCALAR_55_DIRECT_DEPTH),
        .S_AXIS_SCALAR_56_DIRECT_DEPTH(S_AXIS_SCALAR_56_DIRECT_DEPTH),
        .S_AXIS_SCALAR_57_DIRECT_DEPTH(S_AXIS_SCALAR_57_DIRECT_DEPTH),
        .S_AXIS_SCALAR_58_DIRECT_DEPTH(S_AXIS_SCALAR_58_DIRECT_DEPTH),
        .S_AXIS_SCALAR_59_DIRECT_DEPTH(S_AXIS_SCALAR_59_DIRECT_DEPTH),
        .S_AXIS_SCALAR_60_DIRECT_DEPTH(S_AXIS_SCALAR_60_DIRECT_DEPTH),
        .S_AXIS_SCALAR_61_DIRECT_DEPTH(S_AXIS_SCALAR_61_DIRECT_DEPTH),
        .S_AXIS_SCALAR_62_DIRECT_DEPTH(S_AXIS_SCALAR_62_DIRECT_DEPTH),
        .S_AXIS_SCALAR_63_DIRECT_DEPTH(S_AXIS_SCALAR_63_DIRECT_DEPTH),
        .S_AXIS_SCALAR_64_DIRECT_DEPTH(S_AXIS_SCALAR_64_DIRECT_DEPTH),
        .S_AXIS_SCALAR_65_DIRECT_DEPTH(S_AXIS_SCALAR_65_DIRECT_DEPTH),
        .S_AXIS_SCALAR_66_DIRECT_DEPTH(S_AXIS_SCALAR_66_DIRECT_DEPTH),
        .S_AXIS_SCALAR_67_DIRECT_DEPTH(S_AXIS_SCALAR_67_DIRECT_DEPTH),
        .S_AXIS_SCALAR_68_DIRECT_DEPTH(S_AXIS_SCALAR_68_DIRECT_DEPTH),
        .S_AXIS_SCALAR_69_DIRECT_DEPTH(S_AXIS_SCALAR_69_DIRECT_DEPTH),
        .S_AXIS_SCALAR_70_DIRECT_DEPTH(S_AXIS_SCALAR_70_DIRECT_DEPTH),
        .S_AXIS_SCALAR_71_DIRECT_DEPTH(S_AXIS_SCALAR_71_DIRECT_DEPTH),
        .S_AXIS_SCALAR_72_DIRECT_DEPTH(S_AXIS_SCALAR_72_DIRECT_DEPTH),
        .S_AXIS_SCALAR_73_DIRECT_DEPTH(S_AXIS_SCALAR_73_DIRECT_DEPTH),
        .S_AXIS_SCALAR_74_DIRECT_DEPTH(S_AXIS_SCALAR_74_DIRECT_DEPTH),
        .S_AXIS_SCALAR_75_DIRECT_DEPTH(S_AXIS_SCALAR_75_DIRECT_DEPTH),
        .S_AXIS_SCALAR_76_DIRECT_DEPTH(S_AXIS_SCALAR_76_DIRECT_DEPTH),
        .S_AXIS_SCALAR_77_DIRECT_DEPTH(S_AXIS_SCALAR_77_DIRECT_DEPTH),
        .S_AXIS_SCALAR_78_DIRECT_DEPTH(S_AXIS_SCALAR_78_DIRECT_DEPTH),
        .S_AXIS_SCALAR_79_DIRECT_DEPTH(S_AXIS_SCALAR_79_DIRECT_DEPTH),
        .S_AXIS_SCALAR_80_DIRECT_DEPTH(S_AXIS_SCALAR_80_DIRECT_DEPTH),
        .S_AXIS_SCALAR_81_DIRECT_DEPTH(S_AXIS_SCALAR_81_DIRECT_DEPTH),
        .S_AXIS_SCALAR_82_DIRECT_DEPTH(S_AXIS_SCALAR_82_DIRECT_DEPTH),
        .S_AXIS_SCALAR_83_DIRECT_DEPTH(S_AXIS_SCALAR_83_DIRECT_DEPTH),
        .S_AXIS_SCALAR_84_DIRECT_DEPTH(S_AXIS_SCALAR_84_DIRECT_DEPTH),
        .S_AXIS_SCALAR_85_DIRECT_DEPTH(S_AXIS_SCALAR_85_DIRECT_DEPTH),
        .S_AXIS_SCALAR_86_DIRECT_DEPTH(S_AXIS_SCALAR_86_DIRECT_DEPTH),
        .S_AXIS_SCALAR_87_DIRECT_DEPTH(S_AXIS_SCALAR_87_DIRECT_DEPTH),
        .S_AXIS_SCALAR_88_DIRECT_DEPTH(S_AXIS_SCALAR_88_DIRECT_DEPTH),
        .S_AXIS_SCALAR_89_DIRECT_DEPTH(S_AXIS_SCALAR_89_DIRECT_DEPTH),
        .S_AXIS_SCALAR_90_DIRECT_DEPTH(S_AXIS_SCALAR_90_DIRECT_DEPTH),
        .S_AXIS_SCALAR_91_DIRECT_DEPTH(S_AXIS_SCALAR_91_DIRECT_DEPTH),
        .S_AXIS_SCALAR_92_DIRECT_DEPTH(S_AXIS_SCALAR_92_DIRECT_DEPTH),
        .S_AXIS_SCALAR_93_DIRECT_DEPTH(S_AXIS_SCALAR_93_DIRECT_DEPTH),
        .S_AXIS_SCALAR_94_DIRECT_DEPTH(S_AXIS_SCALAR_94_DIRECT_DEPTH),
        .S_AXIS_SCALAR_95_DIRECT_DEPTH(S_AXIS_SCALAR_95_DIRECT_DEPTH),
        .S_AXIS_SCALAR_96_DIRECT_DEPTH(S_AXIS_SCALAR_96_DIRECT_DEPTH),
        .S_AXIS_SCALAR_97_DIRECT_DEPTH(S_AXIS_SCALAR_97_DIRECT_DEPTH),
        .S_AXIS_SCALAR_98_DIRECT_DEPTH(S_AXIS_SCALAR_98_DIRECT_DEPTH),
        .S_AXIS_SCALAR_99_DIRECT_DEPTH(S_AXIS_SCALAR_99_DIRECT_DEPTH),
        .S_AXIS_SCALAR_100_DIRECT_DEPTH(S_AXIS_SCALAR_100_DIRECT_DEPTH),
        .S_AXIS_SCALAR_101_DIRECT_DEPTH(S_AXIS_SCALAR_101_DIRECT_DEPTH),
        .S_AXIS_SCALAR_102_DIRECT_DEPTH(S_AXIS_SCALAR_102_DIRECT_DEPTH),
        .S_AXIS_SCALAR_103_DIRECT_DEPTH(S_AXIS_SCALAR_103_DIRECT_DEPTH),
        .S_AXIS_SCALAR_104_DIRECT_DEPTH(S_AXIS_SCALAR_104_DIRECT_DEPTH),
        .S_AXIS_SCALAR_105_DIRECT_DEPTH(S_AXIS_SCALAR_105_DIRECT_DEPTH),
        .S_AXIS_SCALAR_106_DIRECT_DEPTH(S_AXIS_SCALAR_106_DIRECT_DEPTH),
        .S_AXIS_SCALAR_107_DIRECT_DEPTH(S_AXIS_SCALAR_107_DIRECT_DEPTH),
        .S_AXIS_SCALAR_108_DIRECT_DEPTH(S_AXIS_SCALAR_108_DIRECT_DEPTH),
        .S_AXIS_SCALAR_109_DIRECT_DEPTH(S_AXIS_SCALAR_109_DIRECT_DEPTH),
        .S_AXIS_SCALAR_110_DIRECT_DEPTH(S_AXIS_SCALAR_110_DIRECT_DEPTH),
        .S_AXIS_SCALAR_111_DIRECT_DEPTH(S_AXIS_SCALAR_111_DIRECT_DEPTH),
        .S_AXIS_SCALAR_112_DIRECT_DEPTH(S_AXIS_SCALAR_112_DIRECT_DEPTH),
        .S_AXIS_SCALAR_113_DIRECT_DEPTH(S_AXIS_SCALAR_113_DIRECT_DEPTH),
        .S_AXIS_SCALAR_114_DIRECT_DEPTH(S_AXIS_SCALAR_114_DIRECT_DEPTH),
        .S_AXIS_SCALAR_115_DIRECT_DEPTH(S_AXIS_SCALAR_115_DIRECT_DEPTH),
        .S_AXIS_SCALAR_116_DIRECT_DEPTH(S_AXIS_SCALAR_116_DIRECT_DEPTH),
        .S_AXIS_SCALAR_117_DIRECT_DEPTH(S_AXIS_SCALAR_117_DIRECT_DEPTH),
        .S_AXIS_SCALAR_118_DIRECT_DEPTH(S_AXIS_SCALAR_118_DIRECT_DEPTH),
        .S_AXIS_SCALAR_119_DIRECT_DEPTH(S_AXIS_SCALAR_119_DIRECT_DEPTH),
        .S_AXIS_SCALAR_120_DIRECT_DEPTH(S_AXIS_SCALAR_120_DIRECT_DEPTH),
        .S_AXIS_SCALAR_121_DIRECT_DEPTH(S_AXIS_SCALAR_121_DIRECT_DEPTH),
        .S_AXIS_SCALAR_122_DIRECT_DEPTH(S_AXIS_SCALAR_122_DIRECT_DEPTH),
        .S_AXIS_SCALAR_123_DIRECT_DEPTH(S_AXIS_SCALAR_123_DIRECT_DEPTH),
        .S_AXIS_SCALAR_124_DIRECT_DEPTH(S_AXIS_SCALAR_124_DIRECT_DEPTH),
        .S_AXIS_SCALAR_125_DIRECT_DEPTH(S_AXIS_SCALAR_125_DIRECT_DEPTH),
        .S_AXIS_SCALAR_126_DIRECT_DEPTH(S_AXIS_SCALAR_126_DIRECT_DEPTH),
        .S_AXIS_SCALAR_127_DIRECT_DEPTH(S_AXIS_SCALAR_127_DIRECT_DEPTH),
        .C_OUTSCALAR_0_BITS(C_OUTPUT_SCALAR_0_WIDTH),
        .C_OUTSCALAR_1_BITS(C_OUTPUT_SCALAR_1_WIDTH),
        .C_OUTSCALAR_2_BITS(C_OUTPUT_SCALAR_2_WIDTH),
        .C_OUTSCALAR_3_BITS(C_OUTPUT_SCALAR_3_WIDTH),
        .C_OUTSCALAR_4_BITS(C_OUTPUT_SCALAR_4_WIDTH),
        .C_OUTSCALAR_5_BITS(C_OUTPUT_SCALAR_5_WIDTH),
        .C_OUTSCALAR_6_BITS(C_OUTPUT_SCALAR_6_WIDTH),
        .C_OUTSCALAR_7_BITS(C_OUTPUT_SCALAR_7_WIDTH),
        .C_OUTSCALAR_8_BITS(C_OUTPUT_SCALAR_8_WIDTH),
        .C_OUTSCALAR_9_BITS(C_OUTPUT_SCALAR_9_WIDTH),
        .C_OUTSCALAR_10_BITS(C_OUTPUT_SCALAR_10_WIDTH),
        .C_OUTSCALAR_11_BITS(C_OUTPUT_SCALAR_11_WIDTH),
        .C_OUTSCALAR_12_BITS(C_OUTPUT_SCALAR_12_WIDTH),
        .C_OUTSCALAR_13_BITS(C_OUTPUT_SCALAR_13_WIDTH),
        .C_OUTSCALAR_14_BITS(C_OUTPUT_SCALAR_14_WIDTH),
        .C_OUTSCALAR_15_BITS(C_OUTPUT_SCALAR_15_WIDTH),
        .C_OUTSCALAR_16_BITS(C_OUTPUT_SCALAR_16_WIDTH),
        .C_OUTSCALAR_17_BITS(C_OUTPUT_SCALAR_17_WIDTH),
        .C_OUTSCALAR_18_BITS(C_OUTPUT_SCALAR_18_WIDTH),
        .C_OUTSCALAR_19_BITS(C_OUTPUT_SCALAR_19_WIDTH),
        .C_OUTSCALAR_20_BITS(C_OUTPUT_SCALAR_20_WIDTH),
        .C_OUTSCALAR_21_BITS(C_OUTPUT_SCALAR_21_WIDTH),
        .C_OUTSCALAR_22_BITS(C_OUTPUT_SCALAR_22_WIDTH),
        .C_OUTSCALAR_23_BITS(C_OUTPUT_SCALAR_23_WIDTH),
        .C_OUTSCALAR_24_BITS(C_OUTPUT_SCALAR_24_WIDTH),
        .C_OUTSCALAR_25_BITS(C_OUTPUT_SCALAR_25_WIDTH),
        .C_OUTSCALAR_26_BITS(C_OUTPUT_SCALAR_26_WIDTH),
        .C_OUTSCALAR_27_BITS(C_OUTPUT_SCALAR_27_WIDTH),
        .C_OUTSCALAR_28_BITS(C_OUTPUT_SCALAR_28_WIDTH),
        .C_OUTSCALAR_29_BITS(C_OUTPUT_SCALAR_29_WIDTH),
        .C_OUTSCALAR_30_BITS(C_OUTPUT_SCALAR_30_WIDTH),
        .C_OUTSCALAR_31_BITS(C_OUTPUT_SCALAR_31_WIDTH),
        .C_OUTSCALAR_32_BITS(C_OUTPUT_SCALAR_32_WIDTH),
        .C_OUTSCALAR_33_BITS(C_OUTPUT_SCALAR_33_WIDTH),
        .C_OUTSCALAR_34_BITS(C_OUTPUT_SCALAR_34_WIDTH),
        .C_OUTSCALAR_35_BITS(C_OUTPUT_SCALAR_35_WIDTH),
        .C_OUTSCALAR_36_BITS(C_OUTPUT_SCALAR_36_WIDTH),
        .C_OUTSCALAR_37_BITS(C_OUTPUT_SCALAR_37_WIDTH),
        .C_OUTSCALAR_38_BITS(C_OUTPUT_SCALAR_38_WIDTH),
        .C_OUTSCALAR_39_BITS(C_OUTPUT_SCALAR_39_WIDTH),
        .C_OUTSCALAR_40_BITS(C_OUTPUT_SCALAR_40_WIDTH),
        .C_OUTSCALAR_41_BITS(C_OUTPUT_SCALAR_41_WIDTH),
        .C_OUTSCALAR_42_BITS(C_OUTPUT_SCALAR_42_WIDTH),
        .C_OUTSCALAR_43_BITS(C_OUTPUT_SCALAR_43_WIDTH),
        .C_OUTSCALAR_44_BITS(C_OUTPUT_SCALAR_44_WIDTH),
        .C_OUTSCALAR_45_BITS(C_OUTPUT_SCALAR_45_WIDTH),
        .C_OUTSCALAR_46_BITS(C_OUTPUT_SCALAR_46_WIDTH),
        .C_OUTSCALAR_47_BITS(C_OUTPUT_SCALAR_47_WIDTH),
        .C_OUTSCALAR_48_BITS(C_OUTPUT_SCALAR_48_WIDTH),
        .C_OUTSCALAR_49_BITS(C_OUTPUT_SCALAR_49_WIDTH),
        .C_OUTSCALAR_50_BITS(C_OUTPUT_SCALAR_50_WIDTH),
        .C_OUTSCALAR_51_BITS(C_OUTPUT_SCALAR_51_WIDTH),
        .C_OUTSCALAR_52_BITS(C_OUTPUT_SCALAR_52_WIDTH),
        .C_OUTSCALAR_53_BITS(C_OUTPUT_SCALAR_53_WIDTH),
        .C_OUTSCALAR_54_BITS(C_OUTPUT_SCALAR_54_WIDTH),
        .C_OUTSCALAR_55_BITS(C_OUTPUT_SCALAR_55_WIDTH),
        .C_OUTSCALAR_56_BITS(C_OUTPUT_SCALAR_56_WIDTH),
        .C_OUTSCALAR_57_BITS(C_OUTPUT_SCALAR_57_WIDTH),
        .C_OUTSCALAR_58_BITS(C_OUTPUT_SCALAR_58_WIDTH),
        .C_OUTSCALAR_59_BITS(C_OUTPUT_SCALAR_59_WIDTH),
        .C_OUTSCALAR_60_BITS(C_OUTPUT_SCALAR_60_WIDTH),
        .C_OUTSCALAR_61_BITS(C_OUTPUT_SCALAR_61_WIDTH),
        .C_OUTSCALAR_62_BITS(C_OUTPUT_SCALAR_62_WIDTH),
        .C_OUTSCALAR_63_BITS(C_OUTPUT_SCALAR_63_WIDTH),
        .C_OUTSCALAR_64_BITS(C_OUTPUT_SCALAR_64_WIDTH),
        .C_OUTSCALAR_65_BITS(C_OUTPUT_SCALAR_65_WIDTH),
        .C_OUTSCALAR_66_BITS(C_OUTPUT_SCALAR_66_WIDTH),
        .C_OUTSCALAR_67_BITS(C_OUTPUT_SCALAR_67_WIDTH),
        .C_OUTSCALAR_68_BITS(C_OUTPUT_SCALAR_68_WIDTH),
        .C_OUTSCALAR_69_BITS(C_OUTPUT_SCALAR_69_WIDTH),
        .C_OUTSCALAR_70_BITS(C_OUTPUT_SCALAR_70_WIDTH),
        .C_OUTSCALAR_71_BITS(C_OUTPUT_SCALAR_71_WIDTH),
        .C_OUTSCALAR_72_BITS(C_OUTPUT_SCALAR_72_WIDTH),
        .C_OUTSCALAR_73_BITS(C_OUTPUT_SCALAR_73_WIDTH),
        .C_OUTSCALAR_74_BITS(C_OUTPUT_SCALAR_74_WIDTH),
        .C_OUTSCALAR_75_BITS(C_OUTPUT_SCALAR_75_WIDTH),
        .C_OUTSCALAR_76_BITS(C_OUTPUT_SCALAR_76_WIDTH),
        .C_OUTSCALAR_77_BITS(C_OUTPUT_SCALAR_77_WIDTH),
        .C_OUTSCALAR_78_BITS(C_OUTPUT_SCALAR_78_WIDTH),
        .C_OUTSCALAR_79_BITS(C_OUTPUT_SCALAR_79_WIDTH),
        .C_OUTSCALAR_80_BITS(C_OUTPUT_SCALAR_80_WIDTH),
        .C_OUTSCALAR_81_BITS(C_OUTPUT_SCALAR_81_WIDTH),
        .C_OUTSCALAR_82_BITS(C_OUTPUT_SCALAR_82_WIDTH),
        .C_OUTSCALAR_83_BITS(C_OUTPUT_SCALAR_83_WIDTH),
        .C_OUTSCALAR_84_BITS(C_OUTPUT_SCALAR_84_WIDTH),
        .C_OUTSCALAR_85_BITS(C_OUTPUT_SCALAR_85_WIDTH),
        .C_OUTSCALAR_86_BITS(C_OUTPUT_SCALAR_86_WIDTH),
        .C_OUTSCALAR_87_BITS(C_OUTPUT_SCALAR_87_WIDTH),
        .C_OUTSCALAR_88_BITS(C_OUTPUT_SCALAR_88_WIDTH),
        .C_OUTSCALAR_89_BITS(C_OUTPUT_SCALAR_89_WIDTH),
        .C_OUTSCALAR_90_BITS(C_OUTPUT_SCALAR_90_WIDTH),
        .C_OUTSCALAR_91_BITS(C_OUTPUT_SCALAR_91_WIDTH),
        .C_OUTSCALAR_92_BITS(C_OUTPUT_SCALAR_92_WIDTH),
        .C_OUTSCALAR_93_BITS(C_OUTPUT_SCALAR_93_WIDTH),
        .C_OUTSCALAR_94_BITS(C_OUTPUT_SCALAR_94_WIDTH),
        .C_OUTSCALAR_95_BITS(C_OUTPUT_SCALAR_95_WIDTH),
        .C_OUTSCALAR_96_BITS(C_OUTPUT_SCALAR_96_WIDTH),
        .C_OUTSCALAR_97_BITS(C_OUTPUT_SCALAR_97_WIDTH),
        .C_OUTSCALAR_98_BITS(C_OUTPUT_SCALAR_98_WIDTH),
        .C_OUTSCALAR_99_BITS(C_OUTPUT_SCALAR_99_WIDTH),
        .C_OUTSCALAR_100_BITS(C_OUTPUT_SCALAR_100_WIDTH),
        .C_OUTSCALAR_101_BITS(C_OUTPUT_SCALAR_101_WIDTH),
        .C_OUTSCALAR_102_BITS(C_OUTPUT_SCALAR_102_WIDTH),
        .C_OUTSCALAR_103_BITS(C_OUTPUT_SCALAR_103_WIDTH),
        .C_OUTSCALAR_104_BITS(C_OUTPUT_SCALAR_104_WIDTH),
        .C_OUTSCALAR_105_BITS(C_OUTPUT_SCALAR_105_WIDTH),
        .C_OUTSCALAR_106_BITS(C_OUTPUT_SCALAR_106_WIDTH),
        .C_OUTSCALAR_107_BITS(C_OUTPUT_SCALAR_107_WIDTH),
        .C_OUTSCALAR_108_BITS(C_OUTPUT_SCALAR_108_WIDTH),
        .C_OUTSCALAR_109_BITS(C_OUTPUT_SCALAR_109_WIDTH),
        .C_OUTSCALAR_110_BITS(C_OUTPUT_SCALAR_110_WIDTH),
        .C_OUTSCALAR_111_BITS(C_OUTPUT_SCALAR_111_WIDTH),
        .C_OUTSCALAR_112_BITS(C_OUTPUT_SCALAR_112_WIDTH),
        .C_OUTSCALAR_113_BITS(C_OUTPUT_SCALAR_113_WIDTH),
        .C_OUTSCALAR_114_BITS(C_OUTPUT_SCALAR_114_WIDTH),
        .C_OUTSCALAR_115_BITS(C_OUTPUT_SCALAR_115_WIDTH),
        .C_OUTSCALAR_116_BITS(C_OUTPUT_SCALAR_116_WIDTH),
        .C_OUTSCALAR_117_BITS(C_OUTPUT_SCALAR_117_WIDTH),
        .C_OUTSCALAR_118_BITS(C_OUTPUT_SCALAR_118_WIDTH),
        .C_OUTSCALAR_119_BITS(C_OUTPUT_SCALAR_119_WIDTH),
        .C_OUTSCALAR_120_BITS(C_OUTPUT_SCALAR_120_WIDTH),
        .C_OUTSCALAR_121_BITS(C_OUTPUT_SCALAR_121_WIDTH),
        .C_OUTSCALAR_122_BITS(C_OUTPUT_SCALAR_122_WIDTH),
        .C_OUTSCALAR_123_BITS(C_OUTPUT_SCALAR_123_WIDTH),
        .C_OUTSCALAR_124_BITS(C_OUTPUT_SCALAR_124_WIDTH),
        .C_OUTSCALAR_125_BITS(C_OUTPUT_SCALAR_125_WIDTH),
        .C_OUTSCALAR_126_BITS(C_OUTPUT_SCALAR_126_WIDTH),
        .C_OUTSCALAR_127_BITS(C_OUTPUT_SCALAR_127_WIDTH),
        .M_AXIS_SCALAR_0_IS_DIRECT(M_AXIS_SCALAR_0_IS_DIRECT),
        .M_AXIS_SCALAR_1_IS_DIRECT(M_AXIS_SCALAR_1_IS_DIRECT),
        .M_AXIS_SCALAR_2_IS_DIRECT(M_AXIS_SCALAR_2_IS_DIRECT),
        .M_AXIS_SCALAR_3_IS_DIRECT(M_AXIS_SCALAR_3_IS_DIRECT),
        .M_AXIS_SCALAR_4_IS_DIRECT(M_AXIS_SCALAR_4_IS_DIRECT),
        .M_AXIS_SCALAR_5_IS_DIRECT(M_AXIS_SCALAR_5_IS_DIRECT),
        .M_AXIS_SCALAR_6_IS_DIRECT(M_AXIS_SCALAR_6_IS_DIRECT),
        .M_AXIS_SCALAR_7_IS_DIRECT(M_AXIS_SCALAR_7_IS_DIRECT),
        .M_AXIS_SCALAR_8_IS_DIRECT(M_AXIS_SCALAR_8_IS_DIRECT),
        .M_AXIS_SCALAR_9_IS_DIRECT(M_AXIS_SCALAR_9_IS_DIRECT),
        .M_AXIS_SCALAR_10_IS_DIRECT(M_AXIS_SCALAR_10_IS_DIRECT),
        .M_AXIS_SCALAR_11_IS_DIRECT(M_AXIS_SCALAR_11_IS_DIRECT),
        .M_AXIS_SCALAR_12_IS_DIRECT(M_AXIS_SCALAR_12_IS_DIRECT),
        .M_AXIS_SCALAR_13_IS_DIRECT(M_AXIS_SCALAR_13_IS_DIRECT),
        .M_AXIS_SCALAR_14_IS_DIRECT(M_AXIS_SCALAR_14_IS_DIRECT),
        .M_AXIS_SCALAR_15_IS_DIRECT(M_AXIS_SCALAR_15_IS_DIRECT),
        .M_AXIS_SCALAR_16_IS_DIRECT(M_AXIS_SCALAR_16_IS_DIRECT),
        .M_AXIS_SCALAR_17_IS_DIRECT(M_AXIS_SCALAR_17_IS_DIRECT),
        .M_AXIS_SCALAR_18_IS_DIRECT(M_AXIS_SCALAR_18_IS_DIRECT),
        .M_AXIS_SCALAR_19_IS_DIRECT(M_AXIS_SCALAR_19_IS_DIRECT),
        .M_AXIS_SCALAR_20_IS_DIRECT(M_AXIS_SCALAR_20_IS_DIRECT),
        .M_AXIS_SCALAR_21_IS_DIRECT(M_AXIS_SCALAR_21_IS_DIRECT),
        .M_AXIS_SCALAR_22_IS_DIRECT(M_AXIS_SCALAR_22_IS_DIRECT),
        .M_AXIS_SCALAR_23_IS_DIRECT(M_AXIS_SCALAR_23_IS_DIRECT),
        .M_AXIS_SCALAR_24_IS_DIRECT(M_AXIS_SCALAR_24_IS_DIRECT),
        .M_AXIS_SCALAR_25_IS_DIRECT(M_AXIS_SCALAR_25_IS_DIRECT),
        .M_AXIS_SCALAR_26_IS_DIRECT(M_AXIS_SCALAR_26_IS_DIRECT),
        .M_AXIS_SCALAR_27_IS_DIRECT(M_AXIS_SCALAR_27_IS_DIRECT),
        .M_AXIS_SCALAR_28_IS_DIRECT(M_AXIS_SCALAR_28_IS_DIRECT),
        .M_AXIS_SCALAR_29_IS_DIRECT(M_AXIS_SCALAR_29_IS_DIRECT),
        .M_AXIS_SCALAR_30_IS_DIRECT(M_AXIS_SCALAR_30_IS_DIRECT),
        .M_AXIS_SCALAR_31_IS_DIRECT(M_AXIS_SCALAR_31_IS_DIRECT),
        .M_AXIS_SCALAR_32_IS_DIRECT(M_AXIS_SCALAR_32_IS_DIRECT),
        .M_AXIS_SCALAR_33_IS_DIRECT(M_AXIS_SCALAR_33_IS_DIRECT),
        .M_AXIS_SCALAR_34_IS_DIRECT(M_AXIS_SCALAR_34_IS_DIRECT),
        .M_AXIS_SCALAR_35_IS_DIRECT(M_AXIS_SCALAR_35_IS_DIRECT),
        .M_AXIS_SCALAR_36_IS_DIRECT(M_AXIS_SCALAR_36_IS_DIRECT),
        .M_AXIS_SCALAR_37_IS_DIRECT(M_AXIS_SCALAR_37_IS_DIRECT),
        .M_AXIS_SCALAR_38_IS_DIRECT(M_AXIS_SCALAR_38_IS_DIRECT),
        .M_AXIS_SCALAR_39_IS_DIRECT(M_AXIS_SCALAR_39_IS_DIRECT),
        .M_AXIS_SCALAR_40_IS_DIRECT(M_AXIS_SCALAR_40_IS_DIRECT),
        .M_AXIS_SCALAR_41_IS_DIRECT(M_AXIS_SCALAR_41_IS_DIRECT),
        .M_AXIS_SCALAR_42_IS_DIRECT(M_AXIS_SCALAR_42_IS_DIRECT),
        .M_AXIS_SCALAR_43_IS_DIRECT(M_AXIS_SCALAR_43_IS_DIRECT),
        .M_AXIS_SCALAR_44_IS_DIRECT(M_AXIS_SCALAR_44_IS_DIRECT),
        .M_AXIS_SCALAR_45_IS_DIRECT(M_AXIS_SCALAR_45_IS_DIRECT),
        .M_AXIS_SCALAR_46_IS_DIRECT(M_AXIS_SCALAR_46_IS_DIRECT),
        .M_AXIS_SCALAR_47_IS_DIRECT(M_AXIS_SCALAR_47_IS_DIRECT),
        .M_AXIS_SCALAR_48_IS_DIRECT(M_AXIS_SCALAR_48_IS_DIRECT),
        .M_AXIS_SCALAR_49_IS_DIRECT(M_AXIS_SCALAR_49_IS_DIRECT),
        .M_AXIS_SCALAR_50_IS_DIRECT(M_AXIS_SCALAR_50_IS_DIRECT),
        .M_AXIS_SCALAR_51_IS_DIRECT(M_AXIS_SCALAR_51_IS_DIRECT),
        .M_AXIS_SCALAR_52_IS_DIRECT(M_AXIS_SCALAR_52_IS_DIRECT),
        .M_AXIS_SCALAR_53_IS_DIRECT(M_AXIS_SCALAR_53_IS_DIRECT),
        .M_AXIS_SCALAR_54_IS_DIRECT(M_AXIS_SCALAR_54_IS_DIRECT),
        .M_AXIS_SCALAR_55_IS_DIRECT(M_AXIS_SCALAR_55_IS_DIRECT),
        .M_AXIS_SCALAR_56_IS_DIRECT(M_AXIS_SCALAR_56_IS_DIRECT),
        .M_AXIS_SCALAR_57_IS_DIRECT(M_AXIS_SCALAR_57_IS_DIRECT),
        .M_AXIS_SCALAR_58_IS_DIRECT(M_AXIS_SCALAR_58_IS_DIRECT),
        .M_AXIS_SCALAR_59_IS_DIRECT(M_AXIS_SCALAR_59_IS_DIRECT),
        .M_AXIS_SCALAR_60_IS_DIRECT(M_AXIS_SCALAR_60_IS_DIRECT),
        .M_AXIS_SCALAR_61_IS_DIRECT(M_AXIS_SCALAR_61_IS_DIRECT),
        .M_AXIS_SCALAR_62_IS_DIRECT(M_AXIS_SCALAR_62_IS_DIRECT),
        .M_AXIS_SCALAR_63_IS_DIRECT(M_AXIS_SCALAR_63_IS_DIRECT),
        .M_AXIS_SCALAR_64_IS_DIRECT(M_AXIS_SCALAR_64_IS_DIRECT),
        .M_AXIS_SCALAR_65_IS_DIRECT(M_AXIS_SCALAR_65_IS_DIRECT),
        .M_AXIS_SCALAR_66_IS_DIRECT(M_AXIS_SCALAR_66_IS_DIRECT),
        .M_AXIS_SCALAR_67_IS_DIRECT(M_AXIS_SCALAR_67_IS_DIRECT),
        .M_AXIS_SCALAR_68_IS_DIRECT(M_AXIS_SCALAR_68_IS_DIRECT),
        .M_AXIS_SCALAR_69_IS_DIRECT(M_AXIS_SCALAR_69_IS_DIRECT),
        .M_AXIS_SCALAR_70_IS_DIRECT(M_AXIS_SCALAR_70_IS_DIRECT),
        .M_AXIS_SCALAR_71_IS_DIRECT(M_AXIS_SCALAR_71_IS_DIRECT),
        .M_AXIS_SCALAR_72_IS_DIRECT(M_AXIS_SCALAR_72_IS_DIRECT),
        .M_AXIS_SCALAR_73_IS_DIRECT(M_AXIS_SCALAR_73_IS_DIRECT),
        .M_AXIS_SCALAR_74_IS_DIRECT(M_AXIS_SCALAR_74_IS_DIRECT),
        .M_AXIS_SCALAR_75_IS_DIRECT(M_AXIS_SCALAR_75_IS_DIRECT),
        .M_AXIS_SCALAR_76_IS_DIRECT(M_AXIS_SCALAR_76_IS_DIRECT),
        .M_AXIS_SCALAR_77_IS_DIRECT(M_AXIS_SCALAR_77_IS_DIRECT),
        .M_AXIS_SCALAR_78_IS_DIRECT(M_AXIS_SCALAR_78_IS_DIRECT),
        .M_AXIS_SCALAR_79_IS_DIRECT(M_AXIS_SCALAR_79_IS_DIRECT),
        .M_AXIS_SCALAR_80_IS_DIRECT(M_AXIS_SCALAR_80_IS_DIRECT),
        .M_AXIS_SCALAR_81_IS_DIRECT(M_AXIS_SCALAR_81_IS_DIRECT),
        .M_AXIS_SCALAR_82_IS_DIRECT(M_AXIS_SCALAR_82_IS_DIRECT),
        .M_AXIS_SCALAR_83_IS_DIRECT(M_AXIS_SCALAR_83_IS_DIRECT),
        .M_AXIS_SCALAR_84_IS_DIRECT(M_AXIS_SCALAR_84_IS_DIRECT),
        .M_AXIS_SCALAR_85_IS_DIRECT(M_AXIS_SCALAR_85_IS_DIRECT),
        .M_AXIS_SCALAR_86_IS_DIRECT(M_AXIS_SCALAR_86_IS_DIRECT),
        .M_AXIS_SCALAR_87_IS_DIRECT(M_AXIS_SCALAR_87_IS_DIRECT),
        .M_AXIS_SCALAR_88_IS_DIRECT(M_AXIS_SCALAR_88_IS_DIRECT),
        .M_AXIS_SCALAR_89_IS_DIRECT(M_AXIS_SCALAR_89_IS_DIRECT),
        .M_AXIS_SCALAR_90_IS_DIRECT(M_AXIS_SCALAR_90_IS_DIRECT),
        .M_AXIS_SCALAR_91_IS_DIRECT(M_AXIS_SCALAR_91_IS_DIRECT),
        .M_AXIS_SCALAR_92_IS_DIRECT(M_AXIS_SCALAR_92_IS_DIRECT),
        .M_AXIS_SCALAR_93_IS_DIRECT(M_AXIS_SCALAR_93_IS_DIRECT),
        .M_AXIS_SCALAR_94_IS_DIRECT(M_AXIS_SCALAR_94_IS_DIRECT),
        .M_AXIS_SCALAR_95_IS_DIRECT(M_AXIS_SCALAR_95_IS_DIRECT),
        .M_AXIS_SCALAR_96_IS_DIRECT(M_AXIS_SCALAR_96_IS_DIRECT),
        .M_AXIS_SCALAR_97_IS_DIRECT(M_AXIS_SCALAR_97_IS_DIRECT),
        .M_AXIS_SCALAR_98_IS_DIRECT(M_AXIS_SCALAR_98_IS_DIRECT),
        .M_AXIS_SCALAR_99_IS_DIRECT(M_AXIS_SCALAR_99_IS_DIRECT),
        .M_AXIS_SCALAR_100_IS_DIRECT(M_AXIS_SCALAR_100_IS_DIRECT),
        .M_AXIS_SCALAR_101_IS_DIRECT(M_AXIS_SCALAR_101_IS_DIRECT),
        .M_AXIS_SCALAR_102_IS_DIRECT(M_AXIS_SCALAR_102_IS_DIRECT),
        .M_AXIS_SCALAR_103_IS_DIRECT(M_AXIS_SCALAR_103_IS_DIRECT),
        .M_AXIS_SCALAR_104_IS_DIRECT(M_AXIS_SCALAR_104_IS_DIRECT),
        .M_AXIS_SCALAR_105_IS_DIRECT(M_AXIS_SCALAR_105_IS_DIRECT),
        .M_AXIS_SCALAR_106_IS_DIRECT(M_AXIS_SCALAR_106_IS_DIRECT),
        .M_AXIS_SCALAR_107_IS_DIRECT(M_AXIS_SCALAR_107_IS_DIRECT),
        .M_AXIS_SCALAR_108_IS_DIRECT(M_AXIS_SCALAR_108_IS_DIRECT),
        .M_AXIS_SCALAR_109_IS_DIRECT(M_AXIS_SCALAR_109_IS_DIRECT),
        .M_AXIS_SCALAR_110_IS_DIRECT(M_AXIS_SCALAR_110_IS_DIRECT),
        .M_AXIS_SCALAR_111_IS_DIRECT(M_AXIS_SCALAR_111_IS_DIRECT),
        .M_AXIS_SCALAR_112_IS_DIRECT(M_AXIS_SCALAR_112_IS_DIRECT),
        .M_AXIS_SCALAR_113_IS_DIRECT(M_AXIS_SCALAR_113_IS_DIRECT),
        .M_AXIS_SCALAR_114_IS_DIRECT(M_AXIS_SCALAR_114_IS_DIRECT),
        .M_AXIS_SCALAR_115_IS_DIRECT(M_AXIS_SCALAR_115_IS_DIRECT),
        .M_AXIS_SCALAR_116_IS_DIRECT(M_AXIS_SCALAR_116_IS_DIRECT),
        .M_AXIS_SCALAR_117_IS_DIRECT(M_AXIS_SCALAR_117_IS_DIRECT),
        .M_AXIS_SCALAR_118_IS_DIRECT(M_AXIS_SCALAR_118_IS_DIRECT),
        .M_AXIS_SCALAR_119_IS_DIRECT(M_AXIS_SCALAR_119_IS_DIRECT),
        .M_AXIS_SCALAR_120_IS_DIRECT(M_AXIS_SCALAR_120_IS_DIRECT),
        .M_AXIS_SCALAR_121_IS_DIRECT(M_AXIS_SCALAR_121_IS_DIRECT),
        .M_AXIS_SCALAR_122_IS_DIRECT(M_AXIS_SCALAR_122_IS_DIRECT),
        .M_AXIS_SCALAR_123_IS_DIRECT(M_AXIS_SCALAR_123_IS_DIRECT),
        .M_AXIS_SCALAR_124_IS_DIRECT(M_AXIS_SCALAR_124_IS_DIRECT),
        .M_AXIS_SCALAR_125_IS_DIRECT(M_AXIS_SCALAR_125_IS_DIRECT),
        .M_AXIS_SCALAR_126_IS_DIRECT(M_AXIS_SCALAR_126_IS_DIRECT),
        .M_AXIS_SCALAR_127_IS_DIRECT(M_AXIS_SCALAR_127_IS_DIRECT),
        .M_AXIS_SCALAR_0_DIRECT_DMWIDTH(M_AXIS_SCALAR_0_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_1_DIRECT_DMWIDTH(M_AXIS_SCALAR_1_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_2_DIRECT_DMWIDTH(M_AXIS_SCALAR_2_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_3_DIRECT_DMWIDTH(M_AXIS_SCALAR_3_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_4_DIRECT_DMWIDTH(M_AXIS_SCALAR_4_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_5_DIRECT_DMWIDTH(M_AXIS_SCALAR_5_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_6_DIRECT_DMWIDTH(M_AXIS_SCALAR_6_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_7_DIRECT_DMWIDTH(M_AXIS_SCALAR_7_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_8_DIRECT_DMWIDTH(M_AXIS_SCALAR_8_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_9_DIRECT_DMWIDTH(M_AXIS_SCALAR_9_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_10_DIRECT_DMWIDTH(M_AXIS_SCALAR_10_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_11_DIRECT_DMWIDTH(M_AXIS_SCALAR_11_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_12_DIRECT_DMWIDTH(M_AXIS_SCALAR_12_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_13_DIRECT_DMWIDTH(M_AXIS_SCALAR_13_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_14_DIRECT_DMWIDTH(M_AXIS_SCALAR_14_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_15_DIRECT_DMWIDTH(M_AXIS_SCALAR_15_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_16_DIRECT_DMWIDTH(M_AXIS_SCALAR_16_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_17_DIRECT_DMWIDTH(M_AXIS_SCALAR_17_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_18_DIRECT_DMWIDTH(M_AXIS_SCALAR_18_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_19_DIRECT_DMWIDTH(M_AXIS_SCALAR_19_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_20_DIRECT_DMWIDTH(M_AXIS_SCALAR_20_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_21_DIRECT_DMWIDTH(M_AXIS_SCALAR_21_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_22_DIRECT_DMWIDTH(M_AXIS_SCALAR_22_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_23_DIRECT_DMWIDTH(M_AXIS_SCALAR_23_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_24_DIRECT_DMWIDTH(M_AXIS_SCALAR_24_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_25_DIRECT_DMWIDTH(M_AXIS_SCALAR_25_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_26_DIRECT_DMWIDTH(M_AXIS_SCALAR_26_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_27_DIRECT_DMWIDTH(M_AXIS_SCALAR_27_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_28_DIRECT_DMWIDTH(M_AXIS_SCALAR_28_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_29_DIRECT_DMWIDTH(M_AXIS_SCALAR_29_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_30_DIRECT_DMWIDTH(M_AXIS_SCALAR_30_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_31_DIRECT_DMWIDTH(M_AXIS_SCALAR_31_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_32_DIRECT_DMWIDTH(M_AXIS_SCALAR_32_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_33_DIRECT_DMWIDTH(M_AXIS_SCALAR_33_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_34_DIRECT_DMWIDTH(M_AXIS_SCALAR_34_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_35_DIRECT_DMWIDTH(M_AXIS_SCALAR_35_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_36_DIRECT_DMWIDTH(M_AXIS_SCALAR_36_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_37_DIRECT_DMWIDTH(M_AXIS_SCALAR_37_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_38_DIRECT_DMWIDTH(M_AXIS_SCALAR_38_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_39_DIRECT_DMWIDTH(M_AXIS_SCALAR_39_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_40_DIRECT_DMWIDTH(M_AXIS_SCALAR_40_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_41_DIRECT_DMWIDTH(M_AXIS_SCALAR_41_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_42_DIRECT_DMWIDTH(M_AXIS_SCALAR_42_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_43_DIRECT_DMWIDTH(M_AXIS_SCALAR_43_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_44_DIRECT_DMWIDTH(M_AXIS_SCALAR_44_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_45_DIRECT_DMWIDTH(M_AXIS_SCALAR_45_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_46_DIRECT_DMWIDTH(M_AXIS_SCALAR_46_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_47_DIRECT_DMWIDTH(M_AXIS_SCALAR_47_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_48_DIRECT_DMWIDTH(M_AXIS_SCALAR_48_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_49_DIRECT_DMWIDTH(M_AXIS_SCALAR_49_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_50_DIRECT_DMWIDTH(M_AXIS_SCALAR_50_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_51_DIRECT_DMWIDTH(M_AXIS_SCALAR_51_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_52_DIRECT_DMWIDTH(M_AXIS_SCALAR_52_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_53_DIRECT_DMWIDTH(M_AXIS_SCALAR_53_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_54_DIRECT_DMWIDTH(M_AXIS_SCALAR_54_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_55_DIRECT_DMWIDTH(M_AXIS_SCALAR_55_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_56_DIRECT_DMWIDTH(M_AXIS_SCALAR_56_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_57_DIRECT_DMWIDTH(M_AXIS_SCALAR_57_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_58_DIRECT_DMWIDTH(M_AXIS_SCALAR_58_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_59_DIRECT_DMWIDTH(M_AXIS_SCALAR_59_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_60_DIRECT_DMWIDTH(M_AXIS_SCALAR_60_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_61_DIRECT_DMWIDTH(M_AXIS_SCALAR_61_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_62_DIRECT_DMWIDTH(M_AXIS_SCALAR_62_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_63_DIRECT_DMWIDTH(M_AXIS_SCALAR_63_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_64_DIRECT_DMWIDTH(M_AXIS_SCALAR_64_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_65_DIRECT_DMWIDTH(M_AXIS_SCALAR_65_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_66_DIRECT_DMWIDTH(M_AXIS_SCALAR_66_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_67_DIRECT_DMWIDTH(M_AXIS_SCALAR_67_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_68_DIRECT_DMWIDTH(M_AXIS_SCALAR_68_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_69_DIRECT_DMWIDTH(M_AXIS_SCALAR_69_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_70_DIRECT_DMWIDTH(M_AXIS_SCALAR_70_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_71_DIRECT_DMWIDTH(M_AXIS_SCALAR_71_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_72_DIRECT_DMWIDTH(M_AXIS_SCALAR_72_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_73_DIRECT_DMWIDTH(M_AXIS_SCALAR_73_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_74_DIRECT_DMWIDTH(M_AXIS_SCALAR_74_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_75_DIRECT_DMWIDTH(M_AXIS_SCALAR_75_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_76_DIRECT_DMWIDTH(M_AXIS_SCALAR_76_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_77_DIRECT_DMWIDTH(M_AXIS_SCALAR_77_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_78_DIRECT_DMWIDTH(M_AXIS_SCALAR_78_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_79_DIRECT_DMWIDTH(M_AXIS_SCALAR_79_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_80_DIRECT_DMWIDTH(M_AXIS_SCALAR_80_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_81_DIRECT_DMWIDTH(M_AXIS_SCALAR_81_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_82_DIRECT_DMWIDTH(M_AXIS_SCALAR_82_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_83_DIRECT_DMWIDTH(M_AXIS_SCALAR_83_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_84_DIRECT_DMWIDTH(M_AXIS_SCALAR_84_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_85_DIRECT_DMWIDTH(M_AXIS_SCALAR_85_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_86_DIRECT_DMWIDTH(M_AXIS_SCALAR_86_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_87_DIRECT_DMWIDTH(M_AXIS_SCALAR_87_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_88_DIRECT_DMWIDTH(M_AXIS_SCALAR_88_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_89_DIRECT_DMWIDTH(M_AXIS_SCALAR_89_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_90_DIRECT_DMWIDTH(M_AXIS_SCALAR_90_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_91_DIRECT_DMWIDTH(M_AXIS_SCALAR_91_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_92_DIRECT_DMWIDTH(M_AXIS_SCALAR_92_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_93_DIRECT_DMWIDTH(M_AXIS_SCALAR_93_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_94_DIRECT_DMWIDTH(M_AXIS_SCALAR_94_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_95_DIRECT_DMWIDTH(M_AXIS_SCALAR_95_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_96_DIRECT_DMWIDTH(M_AXIS_SCALAR_96_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_97_DIRECT_DMWIDTH(M_AXIS_SCALAR_97_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_98_DIRECT_DMWIDTH(M_AXIS_SCALAR_98_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_99_DIRECT_DMWIDTH(M_AXIS_SCALAR_99_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_100_DIRECT_DMWIDTH(M_AXIS_SCALAR_100_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_101_DIRECT_DMWIDTH(M_AXIS_SCALAR_101_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_102_DIRECT_DMWIDTH(M_AXIS_SCALAR_102_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_103_DIRECT_DMWIDTH(M_AXIS_SCALAR_103_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_104_DIRECT_DMWIDTH(M_AXIS_SCALAR_104_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_105_DIRECT_DMWIDTH(M_AXIS_SCALAR_105_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_106_DIRECT_DMWIDTH(M_AXIS_SCALAR_106_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_107_DIRECT_DMWIDTH(M_AXIS_SCALAR_107_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_108_DIRECT_DMWIDTH(M_AXIS_SCALAR_108_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_109_DIRECT_DMWIDTH(M_AXIS_SCALAR_109_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_110_DIRECT_DMWIDTH(M_AXIS_SCALAR_110_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_111_DIRECT_DMWIDTH(M_AXIS_SCALAR_111_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_112_DIRECT_DMWIDTH(M_AXIS_SCALAR_112_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_113_DIRECT_DMWIDTH(M_AXIS_SCALAR_113_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_114_DIRECT_DMWIDTH(M_AXIS_SCALAR_114_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_115_DIRECT_DMWIDTH(M_AXIS_SCALAR_115_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_116_DIRECT_DMWIDTH(M_AXIS_SCALAR_116_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_117_DIRECT_DMWIDTH(M_AXIS_SCALAR_117_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_118_DIRECT_DMWIDTH(M_AXIS_SCALAR_118_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_119_DIRECT_DMWIDTH(M_AXIS_SCALAR_119_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_120_DIRECT_DMWIDTH(M_AXIS_SCALAR_120_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_121_DIRECT_DMWIDTH(M_AXIS_SCALAR_121_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_122_DIRECT_DMWIDTH(M_AXIS_SCALAR_122_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_123_DIRECT_DMWIDTH(M_AXIS_SCALAR_123_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_124_DIRECT_DMWIDTH(M_AXIS_SCALAR_124_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_125_DIRECT_DMWIDTH(M_AXIS_SCALAR_125_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_126_DIRECT_DMWIDTH(M_AXIS_SCALAR_126_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_127_DIRECT_DMWIDTH(M_AXIS_SCALAR_127_DIRECT_DMWIDTH),
        .M_AXIS_SCALAR_0_DIRECT_IS_ASYNC(M_AXIS_SCALAR_0_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_1_DIRECT_IS_ASYNC(M_AXIS_SCALAR_1_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_2_DIRECT_IS_ASYNC(M_AXIS_SCALAR_2_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_3_DIRECT_IS_ASYNC(M_AXIS_SCALAR_3_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_4_DIRECT_IS_ASYNC(M_AXIS_SCALAR_4_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_5_DIRECT_IS_ASYNC(M_AXIS_SCALAR_5_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_6_DIRECT_IS_ASYNC(M_AXIS_SCALAR_6_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_7_DIRECT_IS_ASYNC(M_AXIS_SCALAR_7_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_8_DIRECT_IS_ASYNC(M_AXIS_SCALAR_8_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_9_DIRECT_IS_ASYNC(M_AXIS_SCALAR_9_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_10_DIRECT_IS_ASYNC(M_AXIS_SCALAR_10_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_11_DIRECT_IS_ASYNC(M_AXIS_SCALAR_11_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_12_DIRECT_IS_ASYNC(M_AXIS_SCALAR_12_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_13_DIRECT_IS_ASYNC(M_AXIS_SCALAR_13_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_14_DIRECT_IS_ASYNC(M_AXIS_SCALAR_14_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_15_DIRECT_IS_ASYNC(M_AXIS_SCALAR_15_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_16_DIRECT_IS_ASYNC(M_AXIS_SCALAR_16_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_17_DIRECT_IS_ASYNC(M_AXIS_SCALAR_17_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_18_DIRECT_IS_ASYNC(M_AXIS_SCALAR_18_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_19_DIRECT_IS_ASYNC(M_AXIS_SCALAR_19_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_20_DIRECT_IS_ASYNC(M_AXIS_SCALAR_20_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_21_DIRECT_IS_ASYNC(M_AXIS_SCALAR_21_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_22_DIRECT_IS_ASYNC(M_AXIS_SCALAR_22_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_23_DIRECT_IS_ASYNC(M_AXIS_SCALAR_23_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_24_DIRECT_IS_ASYNC(M_AXIS_SCALAR_24_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_25_DIRECT_IS_ASYNC(M_AXIS_SCALAR_25_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_26_DIRECT_IS_ASYNC(M_AXIS_SCALAR_26_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_27_DIRECT_IS_ASYNC(M_AXIS_SCALAR_27_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_28_DIRECT_IS_ASYNC(M_AXIS_SCALAR_28_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_29_DIRECT_IS_ASYNC(M_AXIS_SCALAR_29_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_30_DIRECT_IS_ASYNC(M_AXIS_SCALAR_30_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_31_DIRECT_IS_ASYNC(M_AXIS_SCALAR_31_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_32_DIRECT_IS_ASYNC(M_AXIS_SCALAR_32_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_33_DIRECT_IS_ASYNC(M_AXIS_SCALAR_33_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_34_DIRECT_IS_ASYNC(M_AXIS_SCALAR_34_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_35_DIRECT_IS_ASYNC(M_AXIS_SCALAR_35_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_36_DIRECT_IS_ASYNC(M_AXIS_SCALAR_36_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_37_DIRECT_IS_ASYNC(M_AXIS_SCALAR_37_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_38_DIRECT_IS_ASYNC(M_AXIS_SCALAR_38_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_39_DIRECT_IS_ASYNC(M_AXIS_SCALAR_39_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_40_DIRECT_IS_ASYNC(M_AXIS_SCALAR_40_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_41_DIRECT_IS_ASYNC(M_AXIS_SCALAR_41_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_42_DIRECT_IS_ASYNC(M_AXIS_SCALAR_42_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_43_DIRECT_IS_ASYNC(M_AXIS_SCALAR_43_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_44_DIRECT_IS_ASYNC(M_AXIS_SCALAR_44_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_45_DIRECT_IS_ASYNC(M_AXIS_SCALAR_45_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_46_DIRECT_IS_ASYNC(M_AXIS_SCALAR_46_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_47_DIRECT_IS_ASYNC(M_AXIS_SCALAR_47_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_48_DIRECT_IS_ASYNC(M_AXIS_SCALAR_48_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_49_DIRECT_IS_ASYNC(M_AXIS_SCALAR_49_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_50_DIRECT_IS_ASYNC(M_AXIS_SCALAR_50_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_51_DIRECT_IS_ASYNC(M_AXIS_SCALAR_51_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_52_DIRECT_IS_ASYNC(M_AXIS_SCALAR_52_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_53_DIRECT_IS_ASYNC(M_AXIS_SCALAR_53_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_54_DIRECT_IS_ASYNC(M_AXIS_SCALAR_54_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_55_DIRECT_IS_ASYNC(M_AXIS_SCALAR_55_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_56_DIRECT_IS_ASYNC(M_AXIS_SCALAR_56_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_57_DIRECT_IS_ASYNC(M_AXIS_SCALAR_57_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_58_DIRECT_IS_ASYNC(M_AXIS_SCALAR_58_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_59_DIRECT_IS_ASYNC(M_AXIS_SCALAR_59_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_60_DIRECT_IS_ASYNC(M_AXIS_SCALAR_60_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_61_DIRECT_IS_ASYNC(M_AXIS_SCALAR_61_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_62_DIRECT_IS_ASYNC(M_AXIS_SCALAR_62_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_63_DIRECT_IS_ASYNC(M_AXIS_SCALAR_63_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_64_DIRECT_IS_ASYNC(M_AXIS_SCALAR_64_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_65_DIRECT_IS_ASYNC(M_AXIS_SCALAR_65_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_66_DIRECT_IS_ASYNC(M_AXIS_SCALAR_66_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_67_DIRECT_IS_ASYNC(M_AXIS_SCALAR_67_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_68_DIRECT_IS_ASYNC(M_AXIS_SCALAR_68_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_69_DIRECT_IS_ASYNC(M_AXIS_SCALAR_69_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_70_DIRECT_IS_ASYNC(M_AXIS_SCALAR_70_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_71_DIRECT_IS_ASYNC(M_AXIS_SCALAR_71_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_72_DIRECT_IS_ASYNC(M_AXIS_SCALAR_72_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_73_DIRECT_IS_ASYNC(M_AXIS_SCALAR_73_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_74_DIRECT_IS_ASYNC(M_AXIS_SCALAR_74_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_75_DIRECT_IS_ASYNC(M_AXIS_SCALAR_75_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_76_DIRECT_IS_ASYNC(M_AXIS_SCALAR_76_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_77_DIRECT_IS_ASYNC(M_AXIS_SCALAR_77_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_78_DIRECT_IS_ASYNC(M_AXIS_SCALAR_78_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_79_DIRECT_IS_ASYNC(M_AXIS_SCALAR_79_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_80_DIRECT_IS_ASYNC(M_AXIS_SCALAR_80_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_81_DIRECT_IS_ASYNC(M_AXIS_SCALAR_81_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_82_DIRECT_IS_ASYNC(M_AXIS_SCALAR_82_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_83_DIRECT_IS_ASYNC(M_AXIS_SCALAR_83_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_84_DIRECT_IS_ASYNC(M_AXIS_SCALAR_84_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_85_DIRECT_IS_ASYNC(M_AXIS_SCALAR_85_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_86_DIRECT_IS_ASYNC(M_AXIS_SCALAR_86_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_87_DIRECT_IS_ASYNC(M_AXIS_SCALAR_87_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_88_DIRECT_IS_ASYNC(M_AXIS_SCALAR_88_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_89_DIRECT_IS_ASYNC(M_AXIS_SCALAR_89_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_90_DIRECT_IS_ASYNC(M_AXIS_SCALAR_90_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_91_DIRECT_IS_ASYNC(M_AXIS_SCALAR_91_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_92_DIRECT_IS_ASYNC(M_AXIS_SCALAR_92_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_93_DIRECT_IS_ASYNC(M_AXIS_SCALAR_93_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_94_DIRECT_IS_ASYNC(M_AXIS_SCALAR_94_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_95_DIRECT_IS_ASYNC(M_AXIS_SCALAR_95_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_96_DIRECT_IS_ASYNC(M_AXIS_SCALAR_96_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_97_DIRECT_IS_ASYNC(M_AXIS_SCALAR_97_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_98_DIRECT_IS_ASYNC(M_AXIS_SCALAR_98_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_99_DIRECT_IS_ASYNC(M_AXIS_SCALAR_99_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_100_DIRECT_IS_ASYNC(M_AXIS_SCALAR_100_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_101_DIRECT_IS_ASYNC(M_AXIS_SCALAR_101_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_102_DIRECT_IS_ASYNC(M_AXIS_SCALAR_102_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_103_DIRECT_IS_ASYNC(M_AXIS_SCALAR_103_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_104_DIRECT_IS_ASYNC(M_AXIS_SCALAR_104_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_105_DIRECT_IS_ASYNC(M_AXIS_SCALAR_105_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_106_DIRECT_IS_ASYNC(M_AXIS_SCALAR_106_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_107_DIRECT_IS_ASYNC(M_AXIS_SCALAR_107_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_108_DIRECT_IS_ASYNC(M_AXIS_SCALAR_108_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_109_DIRECT_IS_ASYNC(M_AXIS_SCALAR_109_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_110_DIRECT_IS_ASYNC(M_AXIS_SCALAR_110_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_111_DIRECT_IS_ASYNC(M_AXIS_SCALAR_111_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_112_DIRECT_IS_ASYNC(M_AXIS_SCALAR_112_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_113_DIRECT_IS_ASYNC(M_AXIS_SCALAR_113_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_114_DIRECT_IS_ASYNC(M_AXIS_SCALAR_114_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_115_DIRECT_IS_ASYNC(M_AXIS_SCALAR_115_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_116_DIRECT_IS_ASYNC(M_AXIS_SCALAR_116_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_117_DIRECT_IS_ASYNC(M_AXIS_SCALAR_117_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_118_DIRECT_IS_ASYNC(M_AXIS_SCALAR_118_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_119_DIRECT_IS_ASYNC(M_AXIS_SCALAR_119_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_120_DIRECT_IS_ASYNC(M_AXIS_SCALAR_120_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_121_DIRECT_IS_ASYNC(M_AXIS_SCALAR_121_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_122_DIRECT_IS_ASYNC(M_AXIS_SCALAR_122_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_123_DIRECT_IS_ASYNC(M_AXIS_SCALAR_123_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_124_DIRECT_IS_ASYNC(M_AXIS_SCALAR_124_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_125_DIRECT_IS_ASYNC(M_AXIS_SCALAR_125_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_126_DIRECT_IS_ASYNC(M_AXIS_SCALAR_126_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_127_DIRECT_IS_ASYNC(M_AXIS_SCALAR_127_DIRECT_IS_ASYNC),
        .M_AXIS_SCALAR_0_DIRECT_DEPTH(M_AXIS_SCALAR_0_DIRECT_DEPTH),
        .M_AXIS_SCALAR_1_DIRECT_DEPTH(M_AXIS_SCALAR_1_DIRECT_DEPTH),
        .M_AXIS_SCALAR_2_DIRECT_DEPTH(M_AXIS_SCALAR_2_DIRECT_DEPTH),
        .M_AXIS_SCALAR_3_DIRECT_DEPTH(M_AXIS_SCALAR_3_DIRECT_DEPTH),
        .M_AXIS_SCALAR_4_DIRECT_DEPTH(M_AXIS_SCALAR_4_DIRECT_DEPTH),
        .M_AXIS_SCALAR_5_DIRECT_DEPTH(M_AXIS_SCALAR_5_DIRECT_DEPTH),
        .M_AXIS_SCALAR_6_DIRECT_DEPTH(M_AXIS_SCALAR_6_DIRECT_DEPTH),
        .M_AXIS_SCALAR_7_DIRECT_DEPTH(M_AXIS_SCALAR_7_DIRECT_DEPTH),
        .M_AXIS_SCALAR_8_DIRECT_DEPTH(M_AXIS_SCALAR_8_DIRECT_DEPTH),
        .M_AXIS_SCALAR_9_DIRECT_DEPTH(M_AXIS_SCALAR_9_DIRECT_DEPTH),
        .M_AXIS_SCALAR_10_DIRECT_DEPTH(M_AXIS_SCALAR_10_DIRECT_DEPTH),
        .M_AXIS_SCALAR_11_DIRECT_DEPTH(M_AXIS_SCALAR_11_DIRECT_DEPTH),
        .M_AXIS_SCALAR_12_DIRECT_DEPTH(M_AXIS_SCALAR_12_DIRECT_DEPTH),
        .M_AXIS_SCALAR_13_DIRECT_DEPTH(M_AXIS_SCALAR_13_DIRECT_DEPTH),
        .M_AXIS_SCALAR_14_DIRECT_DEPTH(M_AXIS_SCALAR_14_DIRECT_DEPTH),
        .M_AXIS_SCALAR_15_DIRECT_DEPTH(M_AXIS_SCALAR_15_DIRECT_DEPTH),
        .M_AXIS_SCALAR_16_DIRECT_DEPTH(M_AXIS_SCALAR_16_DIRECT_DEPTH),
        .M_AXIS_SCALAR_17_DIRECT_DEPTH(M_AXIS_SCALAR_17_DIRECT_DEPTH),
        .M_AXIS_SCALAR_18_DIRECT_DEPTH(M_AXIS_SCALAR_18_DIRECT_DEPTH),
        .M_AXIS_SCALAR_19_DIRECT_DEPTH(M_AXIS_SCALAR_19_DIRECT_DEPTH),
        .M_AXIS_SCALAR_20_DIRECT_DEPTH(M_AXIS_SCALAR_20_DIRECT_DEPTH),
        .M_AXIS_SCALAR_21_DIRECT_DEPTH(M_AXIS_SCALAR_21_DIRECT_DEPTH),
        .M_AXIS_SCALAR_22_DIRECT_DEPTH(M_AXIS_SCALAR_22_DIRECT_DEPTH),
        .M_AXIS_SCALAR_23_DIRECT_DEPTH(M_AXIS_SCALAR_23_DIRECT_DEPTH),
        .M_AXIS_SCALAR_24_DIRECT_DEPTH(M_AXIS_SCALAR_24_DIRECT_DEPTH),
        .M_AXIS_SCALAR_25_DIRECT_DEPTH(M_AXIS_SCALAR_25_DIRECT_DEPTH),
        .M_AXIS_SCALAR_26_DIRECT_DEPTH(M_AXIS_SCALAR_26_DIRECT_DEPTH),
        .M_AXIS_SCALAR_27_DIRECT_DEPTH(M_AXIS_SCALAR_27_DIRECT_DEPTH),
        .M_AXIS_SCALAR_28_DIRECT_DEPTH(M_AXIS_SCALAR_28_DIRECT_DEPTH),
        .M_AXIS_SCALAR_29_DIRECT_DEPTH(M_AXIS_SCALAR_29_DIRECT_DEPTH),
        .M_AXIS_SCALAR_30_DIRECT_DEPTH(M_AXIS_SCALAR_30_DIRECT_DEPTH),
        .M_AXIS_SCALAR_31_DIRECT_DEPTH(M_AXIS_SCALAR_31_DIRECT_DEPTH),
        .M_AXIS_SCALAR_32_DIRECT_DEPTH(M_AXIS_SCALAR_32_DIRECT_DEPTH),
        .M_AXIS_SCALAR_33_DIRECT_DEPTH(M_AXIS_SCALAR_33_DIRECT_DEPTH),
        .M_AXIS_SCALAR_34_DIRECT_DEPTH(M_AXIS_SCALAR_34_DIRECT_DEPTH),
        .M_AXIS_SCALAR_35_DIRECT_DEPTH(M_AXIS_SCALAR_35_DIRECT_DEPTH),
        .M_AXIS_SCALAR_36_DIRECT_DEPTH(M_AXIS_SCALAR_36_DIRECT_DEPTH),
        .M_AXIS_SCALAR_37_DIRECT_DEPTH(M_AXIS_SCALAR_37_DIRECT_DEPTH),
        .M_AXIS_SCALAR_38_DIRECT_DEPTH(M_AXIS_SCALAR_38_DIRECT_DEPTH),
        .M_AXIS_SCALAR_39_DIRECT_DEPTH(M_AXIS_SCALAR_39_DIRECT_DEPTH),
        .M_AXIS_SCALAR_40_DIRECT_DEPTH(M_AXIS_SCALAR_40_DIRECT_DEPTH),
        .M_AXIS_SCALAR_41_DIRECT_DEPTH(M_AXIS_SCALAR_41_DIRECT_DEPTH),
        .M_AXIS_SCALAR_42_DIRECT_DEPTH(M_AXIS_SCALAR_42_DIRECT_DEPTH),
        .M_AXIS_SCALAR_43_DIRECT_DEPTH(M_AXIS_SCALAR_43_DIRECT_DEPTH),
        .M_AXIS_SCALAR_44_DIRECT_DEPTH(M_AXIS_SCALAR_44_DIRECT_DEPTH),
        .M_AXIS_SCALAR_45_DIRECT_DEPTH(M_AXIS_SCALAR_45_DIRECT_DEPTH),
        .M_AXIS_SCALAR_46_DIRECT_DEPTH(M_AXIS_SCALAR_46_DIRECT_DEPTH),
        .M_AXIS_SCALAR_47_DIRECT_DEPTH(M_AXIS_SCALAR_47_DIRECT_DEPTH),
        .M_AXIS_SCALAR_48_DIRECT_DEPTH(M_AXIS_SCALAR_48_DIRECT_DEPTH),
        .M_AXIS_SCALAR_49_DIRECT_DEPTH(M_AXIS_SCALAR_49_DIRECT_DEPTH),
        .M_AXIS_SCALAR_50_DIRECT_DEPTH(M_AXIS_SCALAR_50_DIRECT_DEPTH),
        .M_AXIS_SCALAR_51_DIRECT_DEPTH(M_AXIS_SCALAR_51_DIRECT_DEPTH),
        .M_AXIS_SCALAR_52_DIRECT_DEPTH(M_AXIS_SCALAR_52_DIRECT_DEPTH),
        .M_AXIS_SCALAR_53_DIRECT_DEPTH(M_AXIS_SCALAR_53_DIRECT_DEPTH),
        .M_AXIS_SCALAR_54_DIRECT_DEPTH(M_AXIS_SCALAR_54_DIRECT_DEPTH),
        .M_AXIS_SCALAR_55_DIRECT_DEPTH(M_AXIS_SCALAR_55_DIRECT_DEPTH),
        .M_AXIS_SCALAR_56_DIRECT_DEPTH(M_AXIS_SCALAR_56_DIRECT_DEPTH),
        .M_AXIS_SCALAR_57_DIRECT_DEPTH(M_AXIS_SCALAR_57_DIRECT_DEPTH),
        .M_AXIS_SCALAR_58_DIRECT_DEPTH(M_AXIS_SCALAR_58_DIRECT_DEPTH),
        .M_AXIS_SCALAR_59_DIRECT_DEPTH(M_AXIS_SCALAR_59_DIRECT_DEPTH),
        .M_AXIS_SCALAR_60_DIRECT_DEPTH(M_AXIS_SCALAR_60_DIRECT_DEPTH),
        .M_AXIS_SCALAR_61_DIRECT_DEPTH(M_AXIS_SCALAR_61_DIRECT_DEPTH),
        .M_AXIS_SCALAR_62_DIRECT_DEPTH(M_AXIS_SCALAR_62_DIRECT_DEPTH),
        .M_AXIS_SCALAR_63_DIRECT_DEPTH(M_AXIS_SCALAR_63_DIRECT_DEPTH),
        .M_AXIS_SCALAR_64_DIRECT_DEPTH(M_AXIS_SCALAR_64_DIRECT_DEPTH),
        .M_AXIS_SCALAR_65_DIRECT_DEPTH(M_AXIS_SCALAR_65_DIRECT_DEPTH),
        .M_AXIS_SCALAR_66_DIRECT_DEPTH(M_AXIS_SCALAR_66_DIRECT_DEPTH),
        .M_AXIS_SCALAR_67_DIRECT_DEPTH(M_AXIS_SCALAR_67_DIRECT_DEPTH),
        .M_AXIS_SCALAR_68_DIRECT_DEPTH(M_AXIS_SCALAR_68_DIRECT_DEPTH),
        .M_AXIS_SCALAR_69_DIRECT_DEPTH(M_AXIS_SCALAR_69_DIRECT_DEPTH),
        .M_AXIS_SCALAR_70_DIRECT_DEPTH(M_AXIS_SCALAR_70_DIRECT_DEPTH),
        .M_AXIS_SCALAR_71_DIRECT_DEPTH(M_AXIS_SCALAR_71_DIRECT_DEPTH),
        .M_AXIS_SCALAR_72_DIRECT_DEPTH(M_AXIS_SCALAR_72_DIRECT_DEPTH),
        .M_AXIS_SCALAR_73_DIRECT_DEPTH(M_AXIS_SCALAR_73_DIRECT_DEPTH),
        .M_AXIS_SCALAR_74_DIRECT_DEPTH(M_AXIS_SCALAR_74_DIRECT_DEPTH),
        .M_AXIS_SCALAR_75_DIRECT_DEPTH(M_AXIS_SCALAR_75_DIRECT_DEPTH),
        .M_AXIS_SCALAR_76_DIRECT_DEPTH(M_AXIS_SCALAR_76_DIRECT_DEPTH),
        .M_AXIS_SCALAR_77_DIRECT_DEPTH(M_AXIS_SCALAR_77_DIRECT_DEPTH),
        .M_AXIS_SCALAR_78_DIRECT_DEPTH(M_AXIS_SCALAR_78_DIRECT_DEPTH),
        .M_AXIS_SCALAR_79_DIRECT_DEPTH(M_AXIS_SCALAR_79_DIRECT_DEPTH),
        .M_AXIS_SCALAR_80_DIRECT_DEPTH(M_AXIS_SCALAR_80_DIRECT_DEPTH),
        .M_AXIS_SCALAR_81_DIRECT_DEPTH(M_AXIS_SCALAR_81_DIRECT_DEPTH),
        .M_AXIS_SCALAR_82_DIRECT_DEPTH(M_AXIS_SCALAR_82_DIRECT_DEPTH),
        .M_AXIS_SCALAR_83_DIRECT_DEPTH(M_AXIS_SCALAR_83_DIRECT_DEPTH),
        .M_AXIS_SCALAR_84_DIRECT_DEPTH(M_AXIS_SCALAR_84_DIRECT_DEPTH),
        .M_AXIS_SCALAR_85_DIRECT_DEPTH(M_AXIS_SCALAR_85_DIRECT_DEPTH),
        .M_AXIS_SCALAR_86_DIRECT_DEPTH(M_AXIS_SCALAR_86_DIRECT_DEPTH),
        .M_AXIS_SCALAR_87_DIRECT_DEPTH(M_AXIS_SCALAR_87_DIRECT_DEPTH),
        .M_AXIS_SCALAR_88_DIRECT_DEPTH(M_AXIS_SCALAR_88_DIRECT_DEPTH),
        .M_AXIS_SCALAR_89_DIRECT_DEPTH(M_AXIS_SCALAR_89_DIRECT_DEPTH),
        .M_AXIS_SCALAR_90_DIRECT_DEPTH(M_AXIS_SCALAR_90_DIRECT_DEPTH),
        .M_AXIS_SCALAR_91_DIRECT_DEPTH(M_AXIS_SCALAR_91_DIRECT_DEPTH),
        .M_AXIS_SCALAR_92_DIRECT_DEPTH(M_AXIS_SCALAR_92_DIRECT_DEPTH),
        .M_AXIS_SCALAR_93_DIRECT_DEPTH(M_AXIS_SCALAR_93_DIRECT_DEPTH),
        .M_AXIS_SCALAR_94_DIRECT_DEPTH(M_AXIS_SCALAR_94_DIRECT_DEPTH),
        .M_AXIS_SCALAR_95_DIRECT_DEPTH(M_AXIS_SCALAR_95_DIRECT_DEPTH),
        .M_AXIS_SCALAR_96_DIRECT_DEPTH(M_AXIS_SCALAR_96_DIRECT_DEPTH),
        .M_AXIS_SCALAR_97_DIRECT_DEPTH(M_AXIS_SCALAR_97_DIRECT_DEPTH),
        .M_AXIS_SCALAR_98_DIRECT_DEPTH(M_AXIS_SCALAR_98_DIRECT_DEPTH),
        .M_AXIS_SCALAR_99_DIRECT_DEPTH(M_AXIS_SCALAR_99_DIRECT_DEPTH),
        .M_AXIS_SCALAR_100_DIRECT_DEPTH(M_AXIS_SCALAR_100_DIRECT_DEPTH),
        .M_AXIS_SCALAR_101_DIRECT_DEPTH(M_AXIS_SCALAR_101_DIRECT_DEPTH),
        .M_AXIS_SCALAR_102_DIRECT_DEPTH(M_AXIS_SCALAR_102_DIRECT_DEPTH),
        .M_AXIS_SCALAR_103_DIRECT_DEPTH(M_AXIS_SCALAR_103_DIRECT_DEPTH),
        .M_AXIS_SCALAR_104_DIRECT_DEPTH(M_AXIS_SCALAR_104_DIRECT_DEPTH),
        .M_AXIS_SCALAR_105_DIRECT_DEPTH(M_AXIS_SCALAR_105_DIRECT_DEPTH),
        .M_AXIS_SCALAR_106_DIRECT_DEPTH(M_AXIS_SCALAR_106_DIRECT_DEPTH),
        .M_AXIS_SCALAR_107_DIRECT_DEPTH(M_AXIS_SCALAR_107_DIRECT_DEPTH),
        .M_AXIS_SCALAR_108_DIRECT_DEPTH(M_AXIS_SCALAR_108_DIRECT_DEPTH),
        .M_AXIS_SCALAR_109_DIRECT_DEPTH(M_AXIS_SCALAR_109_DIRECT_DEPTH),
        .M_AXIS_SCALAR_110_DIRECT_DEPTH(M_AXIS_SCALAR_110_DIRECT_DEPTH),
        .M_AXIS_SCALAR_111_DIRECT_DEPTH(M_AXIS_SCALAR_111_DIRECT_DEPTH),
        .M_AXIS_SCALAR_112_DIRECT_DEPTH(M_AXIS_SCALAR_112_DIRECT_DEPTH),
        .M_AXIS_SCALAR_113_DIRECT_DEPTH(M_AXIS_SCALAR_113_DIRECT_DEPTH),
        .M_AXIS_SCALAR_114_DIRECT_DEPTH(M_AXIS_SCALAR_114_DIRECT_DEPTH),
        .M_AXIS_SCALAR_115_DIRECT_DEPTH(M_AXIS_SCALAR_115_DIRECT_DEPTH),
        .M_AXIS_SCALAR_116_DIRECT_DEPTH(M_AXIS_SCALAR_116_DIRECT_DEPTH),
        .M_AXIS_SCALAR_117_DIRECT_DEPTH(M_AXIS_SCALAR_117_DIRECT_DEPTH),
        .M_AXIS_SCALAR_118_DIRECT_DEPTH(M_AXIS_SCALAR_118_DIRECT_DEPTH),
        .M_AXIS_SCALAR_119_DIRECT_DEPTH(M_AXIS_SCALAR_119_DIRECT_DEPTH),
        .M_AXIS_SCALAR_120_DIRECT_DEPTH(M_AXIS_SCALAR_120_DIRECT_DEPTH),
        .M_AXIS_SCALAR_121_DIRECT_DEPTH(M_AXIS_SCALAR_121_DIRECT_DEPTH),
        .M_AXIS_SCALAR_122_DIRECT_DEPTH(M_AXIS_SCALAR_122_DIRECT_DEPTH),
        .M_AXIS_SCALAR_123_DIRECT_DEPTH(M_AXIS_SCALAR_123_DIRECT_DEPTH),
        .M_AXIS_SCALAR_124_DIRECT_DEPTH(M_AXIS_SCALAR_124_DIRECT_DEPTH),
        .M_AXIS_SCALAR_125_DIRECT_DEPTH(M_AXIS_SCALAR_125_DIRECT_DEPTH),
        .M_AXIS_SCALAR_126_DIRECT_DEPTH(M_AXIS_SCALAR_126_DIRECT_DEPTH),
        .M_AXIS_SCALAR_127_DIRECT_DEPTH(M_AXIS_SCALAR_127_DIRECT_DEPTH)
    ) scalar_i (
        .clk(s_axi_aclk),
        .acc_clk(acc_aclk),
        //control interface
        .scalar_read_addr(scalar_read_addr),
        .scalar_re(scalar_re),
        .scalar_dout(scalar_dout),
        .scalar_we(scalar_we),
        .scalar_write_addr(scalar_write_addr),
        .scalar_din(scalar_din),
        .outscalar_capture(ap_done),
        .inscalar_next(inscalar_next),
        .inscalar_fifo_empty(inscalar_fifo_empty),
        .inscalar_fifo_full(inscalar_fifo_full),
        .outscalar_fifo_empty(outscalar_fifo_empty),
        .outscalar_fifo_full(outscalar_fifo_full),
        .outscalar_null_empty(outscalar_null_empty),
        .outscalar_null_dout(outscalar_null_dout),
        .outscalar_null_read(outscalar_null_read),
        .inscalar0(ap_iscalar_0_dout),
        .inscalar1(ap_iscalar_1_dout),
        .inscalar2(ap_iscalar_2_dout),
        .inscalar3(ap_iscalar_3_dout),
        .inscalar4(ap_iscalar_4_dout),
        .inscalar5(ap_iscalar_5_dout),
        .inscalar6(ap_iscalar_6_dout),
        .inscalar7(ap_iscalar_7_dout),
        .inscalar8(ap_iscalar_8_dout),
        .inscalar9(ap_iscalar_9_dout),
        .inscalar10(ap_iscalar_10_dout),
        .inscalar11(ap_iscalar_11_dout),
        .inscalar12(ap_iscalar_12_dout),
        .inscalar13(ap_iscalar_13_dout),
        .inscalar14(ap_iscalar_14_dout),
        .inscalar15(ap_iscalar_15_dout),
        .inscalar16(ap_iscalar_16_dout),
        .inscalar17(ap_iscalar_17_dout),
        .inscalar18(ap_iscalar_18_dout),
        .inscalar19(ap_iscalar_19_dout),
        .inscalar20(ap_iscalar_20_dout),
        .inscalar21(ap_iscalar_21_dout),
        .inscalar22(ap_iscalar_22_dout),
        .inscalar23(ap_iscalar_23_dout),
        .inscalar24(ap_iscalar_24_dout),
        .inscalar25(ap_iscalar_25_dout),
        .inscalar26(ap_iscalar_26_dout),
        .inscalar27(ap_iscalar_27_dout),
        .inscalar28(ap_iscalar_28_dout),
        .inscalar29(ap_iscalar_29_dout),
        .inscalar30(ap_iscalar_30_dout),
        .inscalar31(ap_iscalar_31_dout),
        .inscalar32(ap_iscalar_32_dout),
        .inscalar33(ap_iscalar_33_dout),
        .inscalar34(ap_iscalar_34_dout),
        .inscalar35(ap_iscalar_35_dout),
        .inscalar36(ap_iscalar_36_dout),
        .inscalar37(ap_iscalar_37_dout),
        .inscalar38(ap_iscalar_38_dout),
        .inscalar39(ap_iscalar_39_dout),
        .inscalar40(ap_iscalar_40_dout),
        .inscalar41(ap_iscalar_41_dout),
        .inscalar42(ap_iscalar_42_dout),
        .inscalar43(ap_iscalar_43_dout),
        .inscalar44(ap_iscalar_44_dout),
        .inscalar45(ap_iscalar_45_dout),
        .inscalar46(ap_iscalar_46_dout),
        .inscalar47(ap_iscalar_47_dout),
        .inscalar48(ap_iscalar_48_dout),
        .inscalar49(ap_iscalar_49_dout),
        .inscalar50(ap_iscalar_50_dout),
        .inscalar51(ap_iscalar_51_dout),
        .inscalar52(ap_iscalar_52_dout),
        .inscalar53(ap_iscalar_53_dout),
        .inscalar54(ap_iscalar_54_dout),
        .inscalar55(ap_iscalar_55_dout),
        .inscalar56(ap_iscalar_56_dout),
        .inscalar57(ap_iscalar_57_dout),
        .inscalar58(ap_iscalar_58_dout),
        .inscalar59(ap_iscalar_59_dout),
        .inscalar60(ap_iscalar_60_dout),
        .inscalar61(ap_iscalar_61_dout),
        .inscalar62(ap_iscalar_62_dout),
        .inscalar63(ap_iscalar_63_dout),
        .inscalar64(ap_iscalar_64_dout),
        .inscalar65(ap_iscalar_65_dout),
        .inscalar66(ap_iscalar_66_dout),
        .inscalar67(ap_iscalar_67_dout),
        .inscalar68(ap_iscalar_68_dout),
        .inscalar69(ap_iscalar_69_dout),
        .inscalar70(ap_iscalar_70_dout),
        .inscalar71(ap_iscalar_71_dout),
        .inscalar72(ap_iscalar_72_dout),
        .inscalar73(ap_iscalar_73_dout),
        .inscalar74(ap_iscalar_74_dout),
        .inscalar75(ap_iscalar_75_dout),
        .inscalar76(ap_iscalar_76_dout),
        .inscalar77(ap_iscalar_77_dout),
        .inscalar78(ap_iscalar_78_dout),
        .inscalar79(ap_iscalar_79_dout),
        .inscalar80(ap_iscalar_80_dout),
        .inscalar81(ap_iscalar_81_dout),
        .inscalar82(ap_iscalar_82_dout),
        .inscalar83(ap_iscalar_83_dout),
        .inscalar84(ap_iscalar_84_dout),
        .inscalar85(ap_iscalar_85_dout),
        .inscalar86(ap_iscalar_86_dout),
        .inscalar87(ap_iscalar_87_dout),
        .inscalar88(ap_iscalar_88_dout),
        .inscalar89(ap_iscalar_89_dout),
        .inscalar90(ap_iscalar_90_dout),
        .inscalar91(ap_iscalar_91_dout),
        .inscalar92(ap_iscalar_92_dout),
        .inscalar93(ap_iscalar_93_dout),
        .inscalar94(ap_iscalar_94_dout),
        .inscalar95(ap_iscalar_95_dout),
        .inscalar96(ap_iscalar_96_dout),
        .inscalar97(ap_iscalar_97_dout),
        .inscalar98(ap_iscalar_98_dout),
        .inscalar99(ap_iscalar_99_dout),
        .inscalar100(ap_iscalar_100_dout),
        .inscalar101(ap_iscalar_101_dout),
        .inscalar102(ap_iscalar_102_dout),
        .inscalar103(ap_iscalar_103_dout),
        .inscalar104(ap_iscalar_104_dout),
        .inscalar105(ap_iscalar_105_dout),
        .inscalar106(ap_iscalar_106_dout),
        .inscalar107(ap_iscalar_107_dout),
        .inscalar108(ap_iscalar_108_dout),
        .inscalar109(ap_iscalar_109_dout),
        .inscalar110(ap_iscalar_110_dout),
        .inscalar111(ap_iscalar_111_dout),
        .inscalar112(ap_iscalar_112_dout),
        .inscalar113(ap_iscalar_113_dout),
        .inscalar114(ap_iscalar_114_dout),
        .inscalar115(ap_iscalar_115_dout),
        .inscalar116(ap_iscalar_116_dout),
        .inscalar117(ap_iscalar_117_dout),
        .inscalar118(ap_iscalar_118_dout),
        .inscalar119(ap_iscalar_119_dout),
        .inscalar120(ap_iscalar_120_dout),
        .inscalar121(ap_iscalar_121_dout),
        .inscalar122(ap_iscalar_122_dout),
        .inscalar123(ap_iscalar_123_dout),
        .inscalar124(ap_iscalar_124_dout),
        .inscalar125(ap_iscalar_125_dout),
        .inscalar126(ap_iscalar_126_dout),
        .inscalar127(ap_iscalar_127_dout),
        .s_axis_scalar_0_aclk(s_axis_scalar_0_aclk),
        .s_axis_scalar_0_aresetn(s_axis_scalar_0_aresetn),
        .s_axis_scalar_0_tlast(s_axis_scalar_0_tlast),
        .s_axis_scalar_0_tvalid(s_axis_scalar_0_tvalid),
        .s_axis_scalar_0_tkeep(s_axis_scalar_0_tkeep),
        .s_axis_scalar_0_tstrb(s_axis_scalar_0_tstrb),
        .s_axis_scalar_0_tdata(s_axis_scalar_0_tdata),
        .s_axis_scalar_0_tready(s_axis_scalar_0_tready),
        .s_axis_scalar_1_aclk(s_axis_scalar_1_aclk),
        .s_axis_scalar_1_aresetn(s_axis_scalar_1_aresetn),
        .s_axis_scalar_1_tlast(s_axis_scalar_1_tlast),
        .s_axis_scalar_1_tvalid(s_axis_scalar_1_tvalid),
        .s_axis_scalar_1_tkeep(s_axis_scalar_1_tkeep),
        .s_axis_scalar_1_tstrb(s_axis_scalar_1_tstrb),
        .s_axis_scalar_1_tdata(s_axis_scalar_1_tdata),
        .s_axis_scalar_1_tready(s_axis_scalar_1_tready),
        .s_axis_scalar_2_aclk(s_axis_scalar_2_aclk),
        .s_axis_scalar_2_aresetn(s_axis_scalar_2_aresetn),
        .s_axis_scalar_2_tlast(s_axis_scalar_2_tlast),
        .s_axis_scalar_2_tvalid(s_axis_scalar_2_tvalid),
        .s_axis_scalar_2_tkeep(s_axis_scalar_2_tkeep),
        .s_axis_scalar_2_tstrb(s_axis_scalar_2_tstrb),
        .s_axis_scalar_2_tdata(s_axis_scalar_2_tdata),
        .s_axis_scalar_2_tready(s_axis_scalar_2_tready),
        .s_axis_scalar_3_aclk(s_axis_scalar_3_aclk),
        .s_axis_scalar_3_aresetn(s_axis_scalar_3_aresetn),
        .s_axis_scalar_3_tlast(s_axis_scalar_3_tlast),
        .s_axis_scalar_3_tvalid(s_axis_scalar_3_tvalid),
        .s_axis_scalar_3_tkeep(s_axis_scalar_3_tkeep),
        .s_axis_scalar_3_tstrb(s_axis_scalar_3_tstrb),
        .s_axis_scalar_3_tdata(s_axis_scalar_3_tdata),
        .s_axis_scalar_3_tready(s_axis_scalar_3_tready),
        .s_axis_scalar_4_aclk(s_axis_scalar_4_aclk),
        .s_axis_scalar_4_aresetn(s_axis_scalar_4_aresetn),
        .s_axis_scalar_4_tlast(s_axis_scalar_4_tlast),
        .s_axis_scalar_4_tvalid(s_axis_scalar_4_tvalid),
        .s_axis_scalar_4_tkeep(s_axis_scalar_4_tkeep),
        .s_axis_scalar_4_tstrb(s_axis_scalar_4_tstrb),
        .s_axis_scalar_4_tdata(s_axis_scalar_4_tdata),
        .s_axis_scalar_4_tready(s_axis_scalar_4_tready),
        .s_axis_scalar_5_aclk(s_axis_scalar_5_aclk),
        .s_axis_scalar_5_aresetn(s_axis_scalar_5_aresetn),
        .s_axis_scalar_5_tlast(s_axis_scalar_5_tlast),
        .s_axis_scalar_5_tvalid(s_axis_scalar_5_tvalid),
        .s_axis_scalar_5_tkeep(s_axis_scalar_5_tkeep),
        .s_axis_scalar_5_tstrb(s_axis_scalar_5_tstrb),
        .s_axis_scalar_5_tdata(s_axis_scalar_5_tdata),
        .s_axis_scalar_5_tready(s_axis_scalar_5_tready),
        .s_axis_scalar_6_aclk(s_axis_scalar_6_aclk),
        .s_axis_scalar_6_aresetn(s_axis_scalar_6_aresetn),
        .s_axis_scalar_6_tlast(s_axis_scalar_6_tlast),
        .s_axis_scalar_6_tvalid(s_axis_scalar_6_tvalid),
        .s_axis_scalar_6_tkeep(s_axis_scalar_6_tkeep),
        .s_axis_scalar_6_tstrb(s_axis_scalar_6_tstrb),
        .s_axis_scalar_6_tdata(s_axis_scalar_6_tdata),
        .s_axis_scalar_6_tready(s_axis_scalar_6_tready),
        .s_axis_scalar_7_aclk(s_axis_scalar_7_aclk),
        .s_axis_scalar_7_aresetn(s_axis_scalar_7_aresetn),
        .s_axis_scalar_7_tlast(s_axis_scalar_7_tlast),
        .s_axis_scalar_7_tvalid(s_axis_scalar_7_tvalid),
        .s_axis_scalar_7_tkeep(s_axis_scalar_7_tkeep),
        .s_axis_scalar_7_tstrb(s_axis_scalar_7_tstrb),
        .s_axis_scalar_7_tdata(s_axis_scalar_7_tdata),
        .s_axis_scalar_7_tready(s_axis_scalar_7_tready),
        .s_axis_scalar_8_aclk(s_axis_scalar_8_aclk),
        .s_axis_scalar_8_aresetn(s_axis_scalar_8_aresetn),
        .s_axis_scalar_8_tlast(s_axis_scalar_8_tlast),
        .s_axis_scalar_8_tvalid(s_axis_scalar_8_tvalid),
        .s_axis_scalar_8_tkeep(s_axis_scalar_8_tkeep),
        .s_axis_scalar_8_tstrb(s_axis_scalar_8_tstrb),
        .s_axis_scalar_8_tdata(s_axis_scalar_8_tdata),
        .s_axis_scalar_8_tready(s_axis_scalar_8_tready),
        .s_axis_scalar_9_aclk(s_axis_scalar_9_aclk),
        .s_axis_scalar_9_aresetn(s_axis_scalar_9_aresetn),
        .s_axis_scalar_9_tlast(s_axis_scalar_9_tlast),
        .s_axis_scalar_9_tvalid(s_axis_scalar_9_tvalid),
        .s_axis_scalar_9_tkeep(s_axis_scalar_9_tkeep),
        .s_axis_scalar_9_tstrb(s_axis_scalar_9_tstrb),
        .s_axis_scalar_9_tdata(s_axis_scalar_9_tdata),
        .s_axis_scalar_9_tready(s_axis_scalar_9_tready),
        .s_axis_scalar_10_aclk(s_axis_scalar_10_aclk),
        .s_axis_scalar_10_aresetn(s_axis_scalar_10_aresetn),
        .s_axis_scalar_10_tlast(s_axis_scalar_10_tlast),
        .s_axis_scalar_10_tvalid(s_axis_scalar_10_tvalid),
        .s_axis_scalar_10_tkeep(s_axis_scalar_10_tkeep),
        .s_axis_scalar_10_tstrb(s_axis_scalar_10_tstrb),
        .s_axis_scalar_10_tdata(s_axis_scalar_10_tdata),
        .s_axis_scalar_10_tready(s_axis_scalar_10_tready),
        .s_axis_scalar_11_aclk(s_axis_scalar_11_aclk),
        .s_axis_scalar_11_aresetn(s_axis_scalar_11_aresetn),
        .s_axis_scalar_11_tlast(s_axis_scalar_11_tlast),
        .s_axis_scalar_11_tvalid(s_axis_scalar_11_tvalid),
        .s_axis_scalar_11_tkeep(s_axis_scalar_11_tkeep),
        .s_axis_scalar_11_tstrb(s_axis_scalar_11_tstrb),
        .s_axis_scalar_11_tdata(s_axis_scalar_11_tdata),
        .s_axis_scalar_11_tready(s_axis_scalar_11_tready),
        .s_axis_scalar_12_aclk(s_axis_scalar_12_aclk),
        .s_axis_scalar_12_aresetn(s_axis_scalar_12_aresetn),
        .s_axis_scalar_12_tlast(s_axis_scalar_12_tlast),
        .s_axis_scalar_12_tvalid(s_axis_scalar_12_tvalid),
        .s_axis_scalar_12_tkeep(s_axis_scalar_12_tkeep),
        .s_axis_scalar_12_tstrb(s_axis_scalar_12_tstrb),
        .s_axis_scalar_12_tdata(s_axis_scalar_12_tdata),
        .s_axis_scalar_12_tready(s_axis_scalar_12_tready),
        .s_axis_scalar_13_aclk(s_axis_scalar_13_aclk),
        .s_axis_scalar_13_aresetn(s_axis_scalar_13_aresetn),
        .s_axis_scalar_13_tlast(s_axis_scalar_13_tlast),
        .s_axis_scalar_13_tvalid(s_axis_scalar_13_tvalid),
        .s_axis_scalar_13_tkeep(s_axis_scalar_13_tkeep),
        .s_axis_scalar_13_tstrb(s_axis_scalar_13_tstrb),
        .s_axis_scalar_13_tdata(s_axis_scalar_13_tdata),
        .s_axis_scalar_13_tready(s_axis_scalar_13_tready),
        .s_axis_scalar_14_aclk(s_axis_scalar_14_aclk),
        .s_axis_scalar_14_aresetn(s_axis_scalar_14_aresetn),
        .s_axis_scalar_14_tlast(s_axis_scalar_14_tlast),
        .s_axis_scalar_14_tvalid(s_axis_scalar_14_tvalid),
        .s_axis_scalar_14_tkeep(s_axis_scalar_14_tkeep),
        .s_axis_scalar_14_tstrb(s_axis_scalar_14_tstrb),
        .s_axis_scalar_14_tdata(s_axis_scalar_14_tdata),
        .s_axis_scalar_14_tready(s_axis_scalar_14_tready),
        .s_axis_scalar_15_aclk(s_axis_scalar_15_aclk),
        .s_axis_scalar_15_aresetn(s_axis_scalar_15_aresetn),
        .s_axis_scalar_15_tlast(s_axis_scalar_15_tlast),
        .s_axis_scalar_15_tvalid(s_axis_scalar_15_tvalid),
        .s_axis_scalar_15_tkeep(s_axis_scalar_15_tkeep),
        .s_axis_scalar_15_tstrb(s_axis_scalar_15_tstrb),
        .s_axis_scalar_15_tdata(s_axis_scalar_15_tdata),
        .s_axis_scalar_15_tready(s_axis_scalar_15_tready),
        .s_axis_scalar_16_aclk(s_axis_scalar_16_aclk),
        .s_axis_scalar_16_aresetn(s_axis_scalar_16_aresetn),
        .s_axis_scalar_16_tlast(s_axis_scalar_16_tlast),
        .s_axis_scalar_16_tvalid(s_axis_scalar_16_tvalid),
        .s_axis_scalar_16_tkeep(s_axis_scalar_16_tkeep),
        .s_axis_scalar_16_tstrb(s_axis_scalar_16_tstrb),
        .s_axis_scalar_16_tdata(s_axis_scalar_16_tdata),
        .s_axis_scalar_16_tready(s_axis_scalar_16_tready),
        .s_axis_scalar_17_aclk(s_axis_scalar_17_aclk),
        .s_axis_scalar_17_aresetn(s_axis_scalar_17_aresetn),
        .s_axis_scalar_17_tlast(s_axis_scalar_17_tlast),
        .s_axis_scalar_17_tvalid(s_axis_scalar_17_tvalid),
        .s_axis_scalar_17_tkeep(s_axis_scalar_17_tkeep),
        .s_axis_scalar_17_tstrb(s_axis_scalar_17_tstrb),
        .s_axis_scalar_17_tdata(s_axis_scalar_17_tdata),
        .s_axis_scalar_17_tready(s_axis_scalar_17_tready),
        .s_axis_scalar_18_aclk(s_axis_scalar_18_aclk),
        .s_axis_scalar_18_aresetn(s_axis_scalar_18_aresetn),
        .s_axis_scalar_18_tlast(s_axis_scalar_18_tlast),
        .s_axis_scalar_18_tvalid(s_axis_scalar_18_tvalid),
        .s_axis_scalar_18_tkeep(s_axis_scalar_18_tkeep),
        .s_axis_scalar_18_tstrb(s_axis_scalar_18_tstrb),
        .s_axis_scalar_18_tdata(s_axis_scalar_18_tdata),
        .s_axis_scalar_18_tready(s_axis_scalar_18_tready),
        .s_axis_scalar_19_aclk(s_axis_scalar_19_aclk),
        .s_axis_scalar_19_aresetn(s_axis_scalar_19_aresetn),
        .s_axis_scalar_19_tlast(s_axis_scalar_19_tlast),
        .s_axis_scalar_19_tvalid(s_axis_scalar_19_tvalid),
        .s_axis_scalar_19_tkeep(s_axis_scalar_19_tkeep),
        .s_axis_scalar_19_tstrb(s_axis_scalar_19_tstrb),
        .s_axis_scalar_19_tdata(s_axis_scalar_19_tdata),
        .s_axis_scalar_19_tready(s_axis_scalar_19_tready),
        .s_axis_scalar_20_aclk(s_axis_scalar_20_aclk),
        .s_axis_scalar_20_aresetn(s_axis_scalar_20_aresetn),
        .s_axis_scalar_20_tlast(s_axis_scalar_20_tlast),
        .s_axis_scalar_20_tvalid(s_axis_scalar_20_tvalid),
        .s_axis_scalar_20_tkeep(s_axis_scalar_20_tkeep),
        .s_axis_scalar_20_tstrb(s_axis_scalar_20_tstrb),
        .s_axis_scalar_20_tdata(s_axis_scalar_20_tdata),
        .s_axis_scalar_20_tready(s_axis_scalar_20_tready),
        .s_axis_scalar_21_aclk(s_axis_scalar_21_aclk),
        .s_axis_scalar_21_aresetn(s_axis_scalar_21_aresetn),
        .s_axis_scalar_21_tlast(s_axis_scalar_21_tlast),
        .s_axis_scalar_21_tvalid(s_axis_scalar_21_tvalid),
        .s_axis_scalar_21_tkeep(s_axis_scalar_21_tkeep),
        .s_axis_scalar_21_tstrb(s_axis_scalar_21_tstrb),
        .s_axis_scalar_21_tdata(s_axis_scalar_21_tdata),
        .s_axis_scalar_21_tready(s_axis_scalar_21_tready),
        .s_axis_scalar_22_aclk(s_axis_scalar_22_aclk),
        .s_axis_scalar_22_aresetn(s_axis_scalar_22_aresetn),
        .s_axis_scalar_22_tlast(s_axis_scalar_22_tlast),
        .s_axis_scalar_22_tvalid(s_axis_scalar_22_tvalid),
        .s_axis_scalar_22_tkeep(s_axis_scalar_22_tkeep),
        .s_axis_scalar_22_tstrb(s_axis_scalar_22_tstrb),
        .s_axis_scalar_22_tdata(s_axis_scalar_22_tdata),
        .s_axis_scalar_22_tready(s_axis_scalar_22_tready),
        .s_axis_scalar_23_aclk(s_axis_scalar_23_aclk),
        .s_axis_scalar_23_aresetn(s_axis_scalar_23_aresetn),
        .s_axis_scalar_23_tlast(s_axis_scalar_23_tlast),
        .s_axis_scalar_23_tvalid(s_axis_scalar_23_tvalid),
        .s_axis_scalar_23_tkeep(s_axis_scalar_23_tkeep),
        .s_axis_scalar_23_tstrb(s_axis_scalar_23_tstrb),
        .s_axis_scalar_23_tdata(s_axis_scalar_23_tdata),
        .s_axis_scalar_23_tready(s_axis_scalar_23_tready),
        .s_axis_scalar_24_aclk(s_axis_scalar_24_aclk),
        .s_axis_scalar_24_aresetn(s_axis_scalar_24_aresetn),
        .s_axis_scalar_24_tlast(s_axis_scalar_24_tlast),
        .s_axis_scalar_24_tvalid(s_axis_scalar_24_tvalid),
        .s_axis_scalar_24_tkeep(s_axis_scalar_24_tkeep),
        .s_axis_scalar_24_tstrb(s_axis_scalar_24_tstrb),
        .s_axis_scalar_24_tdata(s_axis_scalar_24_tdata),
        .s_axis_scalar_24_tready(s_axis_scalar_24_tready),
        .s_axis_scalar_25_aclk(s_axis_scalar_25_aclk),
        .s_axis_scalar_25_aresetn(s_axis_scalar_25_aresetn),
        .s_axis_scalar_25_tlast(s_axis_scalar_25_tlast),
        .s_axis_scalar_25_tvalid(s_axis_scalar_25_tvalid),
        .s_axis_scalar_25_tkeep(s_axis_scalar_25_tkeep),
        .s_axis_scalar_25_tstrb(s_axis_scalar_25_tstrb),
        .s_axis_scalar_25_tdata(s_axis_scalar_25_tdata),
        .s_axis_scalar_25_tready(s_axis_scalar_25_tready),
        .s_axis_scalar_26_aclk(s_axis_scalar_26_aclk),
        .s_axis_scalar_26_aresetn(s_axis_scalar_26_aresetn),
        .s_axis_scalar_26_tlast(s_axis_scalar_26_tlast),
        .s_axis_scalar_26_tvalid(s_axis_scalar_26_tvalid),
        .s_axis_scalar_26_tkeep(s_axis_scalar_26_tkeep),
        .s_axis_scalar_26_tstrb(s_axis_scalar_26_tstrb),
        .s_axis_scalar_26_tdata(s_axis_scalar_26_tdata),
        .s_axis_scalar_26_tready(s_axis_scalar_26_tready),
        .s_axis_scalar_27_aclk(s_axis_scalar_27_aclk),
        .s_axis_scalar_27_aresetn(s_axis_scalar_27_aresetn),
        .s_axis_scalar_27_tlast(s_axis_scalar_27_tlast),
        .s_axis_scalar_27_tvalid(s_axis_scalar_27_tvalid),
        .s_axis_scalar_27_tkeep(s_axis_scalar_27_tkeep),
        .s_axis_scalar_27_tstrb(s_axis_scalar_27_tstrb),
        .s_axis_scalar_27_tdata(s_axis_scalar_27_tdata),
        .s_axis_scalar_27_tready(s_axis_scalar_27_tready),
        .s_axis_scalar_28_aclk(s_axis_scalar_28_aclk),
        .s_axis_scalar_28_aresetn(s_axis_scalar_28_aresetn),
        .s_axis_scalar_28_tlast(s_axis_scalar_28_tlast),
        .s_axis_scalar_28_tvalid(s_axis_scalar_28_tvalid),
        .s_axis_scalar_28_tkeep(s_axis_scalar_28_tkeep),
        .s_axis_scalar_28_tstrb(s_axis_scalar_28_tstrb),
        .s_axis_scalar_28_tdata(s_axis_scalar_28_tdata),
        .s_axis_scalar_28_tready(s_axis_scalar_28_tready),
        .s_axis_scalar_29_aclk(s_axis_scalar_29_aclk),
        .s_axis_scalar_29_aresetn(s_axis_scalar_29_aresetn),
        .s_axis_scalar_29_tlast(s_axis_scalar_29_tlast),
        .s_axis_scalar_29_tvalid(s_axis_scalar_29_tvalid),
        .s_axis_scalar_29_tkeep(s_axis_scalar_29_tkeep),
        .s_axis_scalar_29_tstrb(s_axis_scalar_29_tstrb),
        .s_axis_scalar_29_tdata(s_axis_scalar_29_tdata),
        .s_axis_scalar_29_tready(s_axis_scalar_29_tready),
        .s_axis_scalar_30_aclk(s_axis_scalar_30_aclk),
        .s_axis_scalar_30_aresetn(s_axis_scalar_30_aresetn),
        .s_axis_scalar_30_tlast(s_axis_scalar_30_tlast),
        .s_axis_scalar_30_tvalid(s_axis_scalar_30_tvalid),
        .s_axis_scalar_30_tkeep(s_axis_scalar_30_tkeep),
        .s_axis_scalar_30_tstrb(s_axis_scalar_30_tstrb),
        .s_axis_scalar_30_tdata(s_axis_scalar_30_tdata),
        .s_axis_scalar_30_tready(s_axis_scalar_30_tready),
        .s_axis_scalar_31_aclk(s_axis_scalar_31_aclk),
        .s_axis_scalar_31_aresetn(s_axis_scalar_31_aresetn),
        .s_axis_scalar_31_tlast(s_axis_scalar_31_tlast),
        .s_axis_scalar_31_tvalid(s_axis_scalar_31_tvalid),
        .s_axis_scalar_31_tkeep(s_axis_scalar_31_tkeep),
        .s_axis_scalar_31_tstrb(s_axis_scalar_31_tstrb),
        .s_axis_scalar_31_tdata(s_axis_scalar_31_tdata),
        .s_axis_scalar_31_tready(s_axis_scalar_31_tready),
        .s_axis_scalar_32_aclk(s_axis_scalar_32_aclk),
        .s_axis_scalar_32_aresetn(s_axis_scalar_32_aresetn),
        .s_axis_scalar_32_tlast(s_axis_scalar_32_tlast),
        .s_axis_scalar_32_tvalid(s_axis_scalar_32_tvalid),
        .s_axis_scalar_32_tkeep(s_axis_scalar_32_tkeep),
        .s_axis_scalar_32_tstrb(s_axis_scalar_32_tstrb),
        .s_axis_scalar_32_tdata(s_axis_scalar_32_tdata),
        .s_axis_scalar_32_tready(s_axis_scalar_32_tready),
        .s_axis_scalar_33_aclk(s_axis_scalar_33_aclk),
        .s_axis_scalar_33_aresetn(s_axis_scalar_33_aresetn),
        .s_axis_scalar_33_tlast(s_axis_scalar_33_tlast),
        .s_axis_scalar_33_tvalid(s_axis_scalar_33_tvalid),
        .s_axis_scalar_33_tkeep(s_axis_scalar_33_tkeep),
        .s_axis_scalar_33_tstrb(s_axis_scalar_33_tstrb),
        .s_axis_scalar_33_tdata(s_axis_scalar_33_tdata),
        .s_axis_scalar_33_tready(s_axis_scalar_33_tready),
        .s_axis_scalar_34_aclk(s_axis_scalar_34_aclk),
        .s_axis_scalar_34_aresetn(s_axis_scalar_34_aresetn),
        .s_axis_scalar_34_tlast(s_axis_scalar_34_tlast),
        .s_axis_scalar_34_tvalid(s_axis_scalar_34_tvalid),
        .s_axis_scalar_34_tkeep(s_axis_scalar_34_tkeep),
        .s_axis_scalar_34_tstrb(s_axis_scalar_34_tstrb),
        .s_axis_scalar_34_tdata(s_axis_scalar_34_tdata),
        .s_axis_scalar_34_tready(s_axis_scalar_34_tready),
        .s_axis_scalar_35_aclk(s_axis_scalar_35_aclk),
        .s_axis_scalar_35_aresetn(s_axis_scalar_35_aresetn),
        .s_axis_scalar_35_tlast(s_axis_scalar_35_tlast),
        .s_axis_scalar_35_tvalid(s_axis_scalar_35_tvalid),
        .s_axis_scalar_35_tkeep(s_axis_scalar_35_tkeep),
        .s_axis_scalar_35_tstrb(s_axis_scalar_35_tstrb),
        .s_axis_scalar_35_tdata(s_axis_scalar_35_tdata),
        .s_axis_scalar_35_tready(s_axis_scalar_35_tready),
        .s_axis_scalar_36_aclk(s_axis_scalar_36_aclk),
        .s_axis_scalar_36_aresetn(s_axis_scalar_36_aresetn),
        .s_axis_scalar_36_tlast(s_axis_scalar_36_tlast),
        .s_axis_scalar_36_tvalid(s_axis_scalar_36_tvalid),
        .s_axis_scalar_36_tkeep(s_axis_scalar_36_tkeep),
        .s_axis_scalar_36_tstrb(s_axis_scalar_36_tstrb),
        .s_axis_scalar_36_tdata(s_axis_scalar_36_tdata),
        .s_axis_scalar_36_tready(s_axis_scalar_36_tready),
        .s_axis_scalar_37_aclk(s_axis_scalar_37_aclk),
        .s_axis_scalar_37_aresetn(s_axis_scalar_37_aresetn),
        .s_axis_scalar_37_tlast(s_axis_scalar_37_tlast),
        .s_axis_scalar_37_tvalid(s_axis_scalar_37_tvalid),
        .s_axis_scalar_37_tkeep(s_axis_scalar_37_tkeep),
        .s_axis_scalar_37_tstrb(s_axis_scalar_37_tstrb),
        .s_axis_scalar_37_tdata(s_axis_scalar_37_tdata),
        .s_axis_scalar_37_tready(s_axis_scalar_37_tready),
        .s_axis_scalar_38_aclk(s_axis_scalar_38_aclk),
        .s_axis_scalar_38_aresetn(s_axis_scalar_38_aresetn),
        .s_axis_scalar_38_tlast(s_axis_scalar_38_tlast),
        .s_axis_scalar_38_tvalid(s_axis_scalar_38_tvalid),
        .s_axis_scalar_38_tkeep(s_axis_scalar_38_tkeep),
        .s_axis_scalar_38_tstrb(s_axis_scalar_38_tstrb),
        .s_axis_scalar_38_tdata(s_axis_scalar_38_tdata),
        .s_axis_scalar_38_tready(s_axis_scalar_38_tready),
        .s_axis_scalar_39_aclk(s_axis_scalar_39_aclk),
        .s_axis_scalar_39_aresetn(s_axis_scalar_39_aresetn),
        .s_axis_scalar_39_tlast(s_axis_scalar_39_tlast),
        .s_axis_scalar_39_tvalid(s_axis_scalar_39_tvalid),
        .s_axis_scalar_39_tkeep(s_axis_scalar_39_tkeep),
        .s_axis_scalar_39_tstrb(s_axis_scalar_39_tstrb),
        .s_axis_scalar_39_tdata(s_axis_scalar_39_tdata),
        .s_axis_scalar_39_tready(s_axis_scalar_39_tready),
        .s_axis_scalar_40_aclk(s_axis_scalar_40_aclk),
        .s_axis_scalar_40_aresetn(s_axis_scalar_40_aresetn),
        .s_axis_scalar_40_tlast(s_axis_scalar_40_tlast),
        .s_axis_scalar_40_tvalid(s_axis_scalar_40_tvalid),
        .s_axis_scalar_40_tkeep(s_axis_scalar_40_tkeep),
        .s_axis_scalar_40_tstrb(s_axis_scalar_40_tstrb),
        .s_axis_scalar_40_tdata(s_axis_scalar_40_tdata),
        .s_axis_scalar_40_tready(s_axis_scalar_40_tready),
        .s_axis_scalar_41_aclk(s_axis_scalar_41_aclk),
        .s_axis_scalar_41_aresetn(s_axis_scalar_41_aresetn),
        .s_axis_scalar_41_tlast(s_axis_scalar_41_tlast),
        .s_axis_scalar_41_tvalid(s_axis_scalar_41_tvalid),
        .s_axis_scalar_41_tkeep(s_axis_scalar_41_tkeep),
        .s_axis_scalar_41_tstrb(s_axis_scalar_41_tstrb),
        .s_axis_scalar_41_tdata(s_axis_scalar_41_tdata),
        .s_axis_scalar_41_tready(s_axis_scalar_41_tready),
        .s_axis_scalar_42_aclk(s_axis_scalar_42_aclk),
        .s_axis_scalar_42_aresetn(s_axis_scalar_42_aresetn),
        .s_axis_scalar_42_tlast(s_axis_scalar_42_tlast),
        .s_axis_scalar_42_tvalid(s_axis_scalar_42_tvalid),
        .s_axis_scalar_42_tkeep(s_axis_scalar_42_tkeep),
        .s_axis_scalar_42_tstrb(s_axis_scalar_42_tstrb),
        .s_axis_scalar_42_tdata(s_axis_scalar_42_tdata),
        .s_axis_scalar_42_tready(s_axis_scalar_42_tready),
        .s_axis_scalar_43_aclk(s_axis_scalar_43_aclk),
        .s_axis_scalar_43_aresetn(s_axis_scalar_43_aresetn),
        .s_axis_scalar_43_tlast(s_axis_scalar_43_tlast),
        .s_axis_scalar_43_tvalid(s_axis_scalar_43_tvalid),
        .s_axis_scalar_43_tkeep(s_axis_scalar_43_tkeep),
        .s_axis_scalar_43_tstrb(s_axis_scalar_43_tstrb),
        .s_axis_scalar_43_tdata(s_axis_scalar_43_tdata),
        .s_axis_scalar_43_tready(s_axis_scalar_43_tready),
        .s_axis_scalar_44_aclk(s_axis_scalar_44_aclk),
        .s_axis_scalar_44_aresetn(s_axis_scalar_44_aresetn),
        .s_axis_scalar_44_tlast(s_axis_scalar_44_tlast),
        .s_axis_scalar_44_tvalid(s_axis_scalar_44_tvalid),
        .s_axis_scalar_44_tkeep(s_axis_scalar_44_tkeep),
        .s_axis_scalar_44_tstrb(s_axis_scalar_44_tstrb),
        .s_axis_scalar_44_tdata(s_axis_scalar_44_tdata),
        .s_axis_scalar_44_tready(s_axis_scalar_44_tready),
        .s_axis_scalar_45_aclk(s_axis_scalar_45_aclk),
        .s_axis_scalar_45_aresetn(s_axis_scalar_45_aresetn),
        .s_axis_scalar_45_tlast(s_axis_scalar_45_tlast),
        .s_axis_scalar_45_tvalid(s_axis_scalar_45_tvalid),
        .s_axis_scalar_45_tkeep(s_axis_scalar_45_tkeep),
        .s_axis_scalar_45_tstrb(s_axis_scalar_45_tstrb),
        .s_axis_scalar_45_tdata(s_axis_scalar_45_tdata),
        .s_axis_scalar_45_tready(s_axis_scalar_45_tready),
        .s_axis_scalar_46_aclk(s_axis_scalar_46_aclk),
        .s_axis_scalar_46_aresetn(s_axis_scalar_46_aresetn),
        .s_axis_scalar_46_tlast(s_axis_scalar_46_tlast),
        .s_axis_scalar_46_tvalid(s_axis_scalar_46_tvalid),
        .s_axis_scalar_46_tkeep(s_axis_scalar_46_tkeep),
        .s_axis_scalar_46_tstrb(s_axis_scalar_46_tstrb),
        .s_axis_scalar_46_tdata(s_axis_scalar_46_tdata),
        .s_axis_scalar_46_tready(s_axis_scalar_46_tready),
        .s_axis_scalar_47_aclk(s_axis_scalar_47_aclk),
        .s_axis_scalar_47_aresetn(s_axis_scalar_47_aresetn),
        .s_axis_scalar_47_tlast(s_axis_scalar_47_tlast),
        .s_axis_scalar_47_tvalid(s_axis_scalar_47_tvalid),
        .s_axis_scalar_47_tkeep(s_axis_scalar_47_tkeep),
        .s_axis_scalar_47_tstrb(s_axis_scalar_47_tstrb),
        .s_axis_scalar_47_tdata(s_axis_scalar_47_tdata),
        .s_axis_scalar_47_tready(s_axis_scalar_47_tready),
        .s_axis_scalar_48_aclk(s_axis_scalar_48_aclk),
        .s_axis_scalar_48_aresetn(s_axis_scalar_48_aresetn),
        .s_axis_scalar_48_tlast(s_axis_scalar_48_tlast),
        .s_axis_scalar_48_tvalid(s_axis_scalar_48_tvalid),
        .s_axis_scalar_48_tkeep(s_axis_scalar_48_tkeep),
        .s_axis_scalar_48_tstrb(s_axis_scalar_48_tstrb),
        .s_axis_scalar_48_tdata(s_axis_scalar_48_tdata),
        .s_axis_scalar_48_tready(s_axis_scalar_48_tready),
        .s_axis_scalar_49_aclk(s_axis_scalar_49_aclk),
        .s_axis_scalar_49_aresetn(s_axis_scalar_49_aresetn),
        .s_axis_scalar_49_tlast(s_axis_scalar_49_tlast),
        .s_axis_scalar_49_tvalid(s_axis_scalar_49_tvalid),
        .s_axis_scalar_49_tkeep(s_axis_scalar_49_tkeep),
        .s_axis_scalar_49_tstrb(s_axis_scalar_49_tstrb),
        .s_axis_scalar_49_tdata(s_axis_scalar_49_tdata),
        .s_axis_scalar_49_tready(s_axis_scalar_49_tready),
        .s_axis_scalar_50_aclk(s_axis_scalar_50_aclk),
        .s_axis_scalar_50_aresetn(s_axis_scalar_50_aresetn),
        .s_axis_scalar_50_tlast(s_axis_scalar_50_tlast),
        .s_axis_scalar_50_tvalid(s_axis_scalar_50_tvalid),
        .s_axis_scalar_50_tkeep(s_axis_scalar_50_tkeep),
        .s_axis_scalar_50_tstrb(s_axis_scalar_50_tstrb),
        .s_axis_scalar_50_tdata(s_axis_scalar_50_tdata),
        .s_axis_scalar_50_tready(s_axis_scalar_50_tready),
        .s_axis_scalar_51_aclk(s_axis_scalar_51_aclk),
        .s_axis_scalar_51_aresetn(s_axis_scalar_51_aresetn),
        .s_axis_scalar_51_tlast(s_axis_scalar_51_tlast),
        .s_axis_scalar_51_tvalid(s_axis_scalar_51_tvalid),
        .s_axis_scalar_51_tkeep(s_axis_scalar_51_tkeep),
        .s_axis_scalar_51_tstrb(s_axis_scalar_51_tstrb),
        .s_axis_scalar_51_tdata(s_axis_scalar_51_tdata),
        .s_axis_scalar_51_tready(s_axis_scalar_51_tready),
        .s_axis_scalar_52_aclk(s_axis_scalar_52_aclk),
        .s_axis_scalar_52_aresetn(s_axis_scalar_52_aresetn),
        .s_axis_scalar_52_tlast(s_axis_scalar_52_tlast),
        .s_axis_scalar_52_tvalid(s_axis_scalar_52_tvalid),
        .s_axis_scalar_52_tkeep(s_axis_scalar_52_tkeep),
        .s_axis_scalar_52_tstrb(s_axis_scalar_52_tstrb),
        .s_axis_scalar_52_tdata(s_axis_scalar_52_tdata),
        .s_axis_scalar_52_tready(s_axis_scalar_52_tready),
        .s_axis_scalar_53_aclk(s_axis_scalar_53_aclk),
        .s_axis_scalar_53_aresetn(s_axis_scalar_53_aresetn),
        .s_axis_scalar_53_tlast(s_axis_scalar_53_tlast),
        .s_axis_scalar_53_tvalid(s_axis_scalar_53_tvalid),
        .s_axis_scalar_53_tkeep(s_axis_scalar_53_tkeep),
        .s_axis_scalar_53_tstrb(s_axis_scalar_53_tstrb),
        .s_axis_scalar_53_tdata(s_axis_scalar_53_tdata),
        .s_axis_scalar_53_tready(s_axis_scalar_53_tready),
        .s_axis_scalar_54_aclk(s_axis_scalar_54_aclk),
        .s_axis_scalar_54_aresetn(s_axis_scalar_54_aresetn),
        .s_axis_scalar_54_tlast(s_axis_scalar_54_tlast),
        .s_axis_scalar_54_tvalid(s_axis_scalar_54_tvalid),
        .s_axis_scalar_54_tkeep(s_axis_scalar_54_tkeep),
        .s_axis_scalar_54_tstrb(s_axis_scalar_54_tstrb),
        .s_axis_scalar_54_tdata(s_axis_scalar_54_tdata),
        .s_axis_scalar_54_tready(s_axis_scalar_54_tready),
        .s_axis_scalar_55_aclk(s_axis_scalar_55_aclk),
        .s_axis_scalar_55_aresetn(s_axis_scalar_55_aresetn),
        .s_axis_scalar_55_tlast(s_axis_scalar_55_tlast),
        .s_axis_scalar_55_tvalid(s_axis_scalar_55_tvalid),
        .s_axis_scalar_55_tkeep(s_axis_scalar_55_tkeep),
        .s_axis_scalar_55_tstrb(s_axis_scalar_55_tstrb),
        .s_axis_scalar_55_tdata(s_axis_scalar_55_tdata),
        .s_axis_scalar_55_tready(s_axis_scalar_55_tready),
        .s_axis_scalar_56_aclk(s_axis_scalar_56_aclk),
        .s_axis_scalar_56_aresetn(s_axis_scalar_56_aresetn),
        .s_axis_scalar_56_tlast(s_axis_scalar_56_tlast),
        .s_axis_scalar_56_tvalid(s_axis_scalar_56_tvalid),
        .s_axis_scalar_56_tkeep(s_axis_scalar_56_tkeep),
        .s_axis_scalar_56_tstrb(s_axis_scalar_56_tstrb),
        .s_axis_scalar_56_tdata(s_axis_scalar_56_tdata),
        .s_axis_scalar_56_tready(s_axis_scalar_56_tready),
        .s_axis_scalar_57_aclk(s_axis_scalar_57_aclk),
        .s_axis_scalar_57_aresetn(s_axis_scalar_57_aresetn),
        .s_axis_scalar_57_tlast(s_axis_scalar_57_tlast),
        .s_axis_scalar_57_tvalid(s_axis_scalar_57_tvalid),
        .s_axis_scalar_57_tkeep(s_axis_scalar_57_tkeep),
        .s_axis_scalar_57_tstrb(s_axis_scalar_57_tstrb),
        .s_axis_scalar_57_tdata(s_axis_scalar_57_tdata),
        .s_axis_scalar_57_tready(s_axis_scalar_57_tready),
        .s_axis_scalar_58_aclk(s_axis_scalar_58_aclk),
        .s_axis_scalar_58_aresetn(s_axis_scalar_58_aresetn),
        .s_axis_scalar_58_tlast(s_axis_scalar_58_tlast),
        .s_axis_scalar_58_tvalid(s_axis_scalar_58_tvalid),
        .s_axis_scalar_58_tkeep(s_axis_scalar_58_tkeep),
        .s_axis_scalar_58_tstrb(s_axis_scalar_58_tstrb),
        .s_axis_scalar_58_tdata(s_axis_scalar_58_tdata),
        .s_axis_scalar_58_tready(s_axis_scalar_58_tready),
        .s_axis_scalar_59_aclk(s_axis_scalar_59_aclk),
        .s_axis_scalar_59_aresetn(s_axis_scalar_59_aresetn),
        .s_axis_scalar_59_tlast(s_axis_scalar_59_tlast),
        .s_axis_scalar_59_tvalid(s_axis_scalar_59_tvalid),
        .s_axis_scalar_59_tkeep(s_axis_scalar_59_tkeep),
        .s_axis_scalar_59_tstrb(s_axis_scalar_59_tstrb),
        .s_axis_scalar_59_tdata(s_axis_scalar_59_tdata),
        .s_axis_scalar_59_tready(s_axis_scalar_59_tready),
        .s_axis_scalar_60_aclk(s_axis_scalar_60_aclk),
        .s_axis_scalar_60_aresetn(s_axis_scalar_60_aresetn),
        .s_axis_scalar_60_tlast(s_axis_scalar_60_tlast),
        .s_axis_scalar_60_tvalid(s_axis_scalar_60_tvalid),
        .s_axis_scalar_60_tkeep(s_axis_scalar_60_tkeep),
        .s_axis_scalar_60_tstrb(s_axis_scalar_60_tstrb),
        .s_axis_scalar_60_tdata(s_axis_scalar_60_tdata),
        .s_axis_scalar_60_tready(s_axis_scalar_60_tready),
        .s_axis_scalar_61_aclk(s_axis_scalar_61_aclk),
        .s_axis_scalar_61_aresetn(s_axis_scalar_61_aresetn),
        .s_axis_scalar_61_tlast(s_axis_scalar_61_tlast),
        .s_axis_scalar_61_tvalid(s_axis_scalar_61_tvalid),
        .s_axis_scalar_61_tkeep(s_axis_scalar_61_tkeep),
        .s_axis_scalar_61_tstrb(s_axis_scalar_61_tstrb),
        .s_axis_scalar_61_tdata(s_axis_scalar_61_tdata),
        .s_axis_scalar_61_tready(s_axis_scalar_61_tready),
        .s_axis_scalar_62_aclk(s_axis_scalar_62_aclk),
        .s_axis_scalar_62_aresetn(s_axis_scalar_62_aresetn),
        .s_axis_scalar_62_tlast(s_axis_scalar_62_tlast),
        .s_axis_scalar_62_tvalid(s_axis_scalar_62_tvalid),
        .s_axis_scalar_62_tkeep(s_axis_scalar_62_tkeep),
        .s_axis_scalar_62_tstrb(s_axis_scalar_62_tstrb),
        .s_axis_scalar_62_tdata(s_axis_scalar_62_tdata),
        .s_axis_scalar_62_tready(s_axis_scalar_62_tready),
        .s_axis_scalar_63_aclk(s_axis_scalar_63_aclk),
        .s_axis_scalar_63_aresetn(s_axis_scalar_63_aresetn),
        .s_axis_scalar_63_tlast(s_axis_scalar_63_tlast),
        .s_axis_scalar_63_tvalid(s_axis_scalar_63_tvalid),
        .s_axis_scalar_63_tkeep(s_axis_scalar_63_tkeep),
        .s_axis_scalar_63_tstrb(s_axis_scalar_63_tstrb),
        .s_axis_scalar_63_tdata(s_axis_scalar_63_tdata),
        .s_axis_scalar_63_tready(s_axis_scalar_63_tready),
        .s_axis_scalar_64_aclk(s_axis_scalar_64_aclk),
        .s_axis_scalar_64_aresetn(s_axis_scalar_64_aresetn),
        .s_axis_scalar_64_tlast(s_axis_scalar_64_tlast),
        .s_axis_scalar_64_tvalid(s_axis_scalar_64_tvalid),
        .s_axis_scalar_64_tkeep(s_axis_scalar_64_tkeep),
        .s_axis_scalar_64_tstrb(s_axis_scalar_64_tstrb),
        .s_axis_scalar_64_tdata(s_axis_scalar_64_tdata),
        .s_axis_scalar_64_tready(s_axis_scalar_64_tready),
        .s_axis_scalar_65_aclk(s_axis_scalar_65_aclk),
        .s_axis_scalar_65_aresetn(s_axis_scalar_65_aresetn),
        .s_axis_scalar_65_tlast(s_axis_scalar_65_tlast),
        .s_axis_scalar_65_tvalid(s_axis_scalar_65_tvalid),
        .s_axis_scalar_65_tkeep(s_axis_scalar_65_tkeep),
        .s_axis_scalar_65_tstrb(s_axis_scalar_65_tstrb),
        .s_axis_scalar_65_tdata(s_axis_scalar_65_tdata),
        .s_axis_scalar_65_tready(s_axis_scalar_65_tready),
        .s_axis_scalar_66_aclk(s_axis_scalar_66_aclk),
        .s_axis_scalar_66_aresetn(s_axis_scalar_66_aresetn),
        .s_axis_scalar_66_tlast(s_axis_scalar_66_tlast),
        .s_axis_scalar_66_tvalid(s_axis_scalar_66_tvalid),
        .s_axis_scalar_66_tkeep(s_axis_scalar_66_tkeep),
        .s_axis_scalar_66_tstrb(s_axis_scalar_66_tstrb),
        .s_axis_scalar_66_tdata(s_axis_scalar_66_tdata),
        .s_axis_scalar_66_tready(s_axis_scalar_66_tready),
        .s_axis_scalar_67_aclk(s_axis_scalar_67_aclk),
        .s_axis_scalar_67_aresetn(s_axis_scalar_67_aresetn),
        .s_axis_scalar_67_tlast(s_axis_scalar_67_tlast),
        .s_axis_scalar_67_tvalid(s_axis_scalar_67_tvalid),
        .s_axis_scalar_67_tkeep(s_axis_scalar_67_tkeep),
        .s_axis_scalar_67_tstrb(s_axis_scalar_67_tstrb),
        .s_axis_scalar_67_tdata(s_axis_scalar_67_tdata),
        .s_axis_scalar_67_tready(s_axis_scalar_67_tready),
        .s_axis_scalar_68_aclk(s_axis_scalar_68_aclk),
        .s_axis_scalar_68_aresetn(s_axis_scalar_68_aresetn),
        .s_axis_scalar_68_tlast(s_axis_scalar_68_tlast),
        .s_axis_scalar_68_tvalid(s_axis_scalar_68_tvalid),
        .s_axis_scalar_68_tkeep(s_axis_scalar_68_tkeep),
        .s_axis_scalar_68_tstrb(s_axis_scalar_68_tstrb),
        .s_axis_scalar_68_tdata(s_axis_scalar_68_tdata),
        .s_axis_scalar_68_tready(s_axis_scalar_68_tready),
        .s_axis_scalar_69_aclk(s_axis_scalar_69_aclk),
        .s_axis_scalar_69_aresetn(s_axis_scalar_69_aresetn),
        .s_axis_scalar_69_tlast(s_axis_scalar_69_tlast),
        .s_axis_scalar_69_tvalid(s_axis_scalar_69_tvalid),
        .s_axis_scalar_69_tkeep(s_axis_scalar_69_tkeep),
        .s_axis_scalar_69_tstrb(s_axis_scalar_69_tstrb),
        .s_axis_scalar_69_tdata(s_axis_scalar_69_tdata),
        .s_axis_scalar_69_tready(s_axis_scalar_69_tready),
        .s_axis_scalar_70_aclk(s_axis_scalar_70_aclk),
        .s_axis_scalar_70_aresetn(s_axis_scalar_70_aresetn),
        .s_axis_scalar_70_tlast(s_axis_scalar_70_tlast),
        .s_axis_scalar_70_tvalid(s_axis_scalar_70_tvalid),
        .s_axis_scalar_70_tkeep(s_axis_scalar_70_tkeep),
        .s_axis_scalar_70_tstrb(s_axis_scalar_70_tstrb),
        .s_axis_scalar_70_tdata(s_axis_scalar_70_tdata),
        .s_axis_scalar_70_tready(s_axis_scalar_70_tready),
        .s_axis_scalar_71_aclk(s_axis_scalar_71_aclk),
        .s_axis_scalar_71_aresetn(s_axis_scalar_71_aresetn),
        .s_axis_scalar_71_tlast(s_axis_scalar_71_tlast),
        .s_axis_scalar_71_tvalid(s_axis_scalar_71_tvalid),
        .s_axis_scalar_71_tkeep(s_axis_scalar_71_tkeep),
        .s_axis_scalar_71_tstrb(s_axis_scalar_71_tstrb),
        .s_axis_scalar_71_tdata(s_axis_scalar_71_tdata),
        .s_axis_scalar_71_tready(s_axis_scalar_71_tready),
        .s_axis_scalar_72_aclk(s_axis_scalar_72_aclk),
        .s_axis_scalar_72_aresetn(s_axis_scalar_72_aresetn),
        .s_axis_scalar_72_tlast(s_axis_scalar_72_tlast),
        .s_axis_scalar_72_tvalid(s_axis_scalar_72_tvalid),
        .s_axis_scalar_72_tkeep(s_axis_scalar_72_tkeep),
        .s_axis_scalar_72_tstrb(s_axis_scalar_72_tstrb),
        .s_axis_scalar_72_tdata(s_axis_scalar_72_tdata),
        .s_axis_scalar_72_tready(s_axis_scalar_72_tready),
        .s_axis_scalar_73_aclk(s_axis_scalar_73_aclk),
        .s_axis_scalar_73_aresetn(s_axis_scalar_73_aresetn),
        .s_axis_scalar_73_tlast(s_axis_scalar_73_tlast),
        .s_axis_scalar_73_tvalid(s_axis_scalar_73_tvalid),
        .s_axis_scalar_73_tkeep(s_axis_scalar_73_tkeep),
        .s_axis_scalar_73_tstrb(s_axis_scalar_73_tstrb),
        .s_axis_scalar_73_tdata(s_axis_scalar_73_tdata),
        .s_axis_scalar_73_tready(s_axis_scalar_73_tready),
        .s_axis_scalar_74_aclk(s_axis_scalar_74_aclk),
        .s_axis_scalar_74_aresetn(s_axis_scalar_74_aresetn),
        .s_axis_scalar_74_tlast(s_axis_scalar_74_tlast),
        .s_axis_scalar_74_tvalid(s_axis_scalar_74_tvalid),
        .s_axis_scalar_74_tkeep(s_axis_scalar_74_tkeep),
        .s_axis_scalar_74_tstrb(s_axis_scalar_74_tstrb),
        .s_axis_scalar_74_tdata(s_axis_scalar_74_tdata),
        .s_axis_scalar_74_tready(s_axis_scalar_74_tready),
        .s_axis_scalar_75_aclk(s_axis_scalar_75_aclk),
        .s_axis_scalar_75_aresetn(s_axis_scalar_75_aresetn),
        .s_axis_scalar_75_tlast(s_axis_scalar_75_tlast),
        .s_axis_scalar_75_tvalid(s_axis_scalar_75_tvalid),
        .s_axis_scalar_75_tkeep(s_axis_scalar_75_tkeep),
        .s_axis_scalar_75_tstrb(s_axis_scalar_75_tstrb),
        .s_axis_scalar_75_tdata(s_axis_scalar_75_tdata),
        .s_axis_scalar_75_tready(s_axis_scalar_75_tready),
        .s_axis_scalar_76_aclk(s_axis_scalar_76_aclk),
        .s_axis_scalar_76_aresetn(s_axis_scalar_76_aresetn),
        .s_axis_scalar_76_tlast(s_axis_scalar_76_tlast),
        .s_axis_scalar_76_tvalid(s_axis_scalar_76_tvalid),
        .s_axis_scalar_76_tkeep(s_axis_scalar_76_tkeep),
        .s_axis_scalar_76_tstrb(s_axis_scalar_76_tstrb),
        .s_axis_scalar_76_tdata(s_axis_scalar_76_tdata),
        .s_axis_scalar_76_tready(s_axis_scalar_76_tready),
        .s_axis_scalar_77_aclk(s_axis_scalar_77_aclk),
        .s_axis_scalar_77_aresetn(s_axis_scalar_77_aresetn),
        .s_axis_scalar_77_tlast(s_axis_scalar_77_tlast),
        .s_axis_scalar_77_tvalid(s_axis_scalar_77_tvalid),
        .s_axis_scalar_77_tkeep(s_axis_scalar_77_tkeep),
        .s_axis_scalar_77_tstrb(s_axis_scalar_77_tstrb),
        .s_axis_scalar_77_tdata(s_axis_scalar_77_tdata),
        .s_axis_scalar_77_tready(s_axis_scalar_77_tready),
        .s_axis_scalar_78_aclk(s_axis_scalar_78_aclk),
        .s_axis_scalar_78_aresetn(s_axis_scalar_78_aresetn),
        .s_axis_scalar_78_tlast(s_axis_scalar_78_tlast),
        .s_axis_scalar_78_tvalid(s_axis_scalar_78_tvalid),
        .s_axis_scalar_78_tkeep(s_axis_scalar_78_tkeep),
        .s_axis_scalar_78_tstrb(s_axis_scalar_78_tstrb),
        .s_axis_scalar_78_tdata(s_axis_scalar_78_tdata),
        .s_axis_scalar_78_tready(s_axis_scalar_78_tready),
        .s_axis_scalar_79_aclk(s_axis_scalar_79_aclk),
        .s_axis_scalar_79_aresetn(s_axis_scalar_79_aresetn),
        .s_axis_scalar_79_tlast(s_axis_scalar_79_tlast),
        .s_axis_scalar_79_tvalid(s_axis_scalar_79_tvalid),
        .s_axis_scalar_79_tkeep(s_axis_scalar_79_tkeep),
        .s_axis_scalar_79_tstrb(s_axis_scalar_79_tstrb),
        .s_axis_scalar_79_tdata(s_axis_scalar_79_tdata),
        .s_axis_scalar_79_tready(s_axis_scalar_79_tready),
        .s_axis_scalar_80_aclk(s_axis_scalar_80_aclk),
        .s_axis_scalar_80_aresetn(s_axis_scalar_80_aresetn),
        .s_axis_scalar_80_tlast(s_axis_scalar_80_tlast),
        .s_axis_scalar_80_tvalid(s_axis_scalar_80_tvalid),
        .s_axis_scalar_80_tkeep(s_axis_scalar_80_tkeep),
        .s_axis_scalar_80_tstrb(s_axis_scalar_80_tstrb),
        .s_axis_scalar_80_tdata(s_axis_scalar_80_tdata),
        .s_axis_scalar_80_tready(s_axis_scalar_80_tready),
        .s_axis_scalar_81_aclk(s_axis_scalar_81_aclk),
        .s_axis_scalar_81_aresetn(s_axis_scalar_81_aresetn),
        .s_axis_scalar_81_tlast(s_axis_scalar_81_tlast),
        .s_axis_scalar_81_tvalid(s_axis_scalar_81_tvalid),
        .s_axis_scalar_81_tkeep(s_axis_scalar_81_tkeep),
        .s_axis_scalar_81_tstrb(s_axis_scalar_81_tstrb),
        .s_axis_scalar_81_tdata(s_axis_scalar_81_tdata),
        .s_axis_scalar_81_tready(s_axis_scalar_81_tready),
        .s_axis_scalar_82_aclk(s_axis_scalar_82_aclk),
        .s_axis_scalar_82_aresetn(s_axis_scalar_82_aresetn),
        .s_axis_scalar_82_tlast(s_axis_scalar_82_tlast),
        .s_axis_scalar_82_tvalid(s_axis_scalar_82_tvalid),
        .s_axis_scalar_82_tkeep(s_axis_scalar_82_tkeep),
        .s_axis_scalar_82_tstrb(s_axis_scalar_82_tstrb),
        .s_axis_scalar_82_tdata(s_axis_scalar_82_tdata),
        .s_axis_scalar_82_tready(s_axis_scalar_82_tready),
        .s_axis_scalar_83_aclk(s_axis_scalar_83_aclk),
        .s_axis_scalar_83_aresetn(s_axis_scalar_83_aresetn),
        .s_axis_scalar_83_tlast(s_axis_scalar_83_tlast),
        .s_axis_scalar_83_tvalid(s_axis_scalar_83_tvalid),
        .s_axis_scalar_83_tkeep(s_axis_scalar_83_tkeep),
        .s_axis_scalar_83_tstrb(s_axis_scalar_83_tstrb),
        .s_axis_scalar_83_tdata(s_axis_scalar_83_tdata),
        .s_axis_scalar_83_tready(s_axis_scalar_83_tready),
        .s_axis_scalar_84_aclk(s_axis_scalar_84_aclk),
        .s_axis_scalar_84_aresetn(s_axis_scalar_84_aresetn),
        .s_axis_scalar_84_tlast(s_axis_scalar_84_tlast),
        .s_axis_scalar_84_tvalid(s_axis_scalar_84_tvalid),
        .s_axis_scalar_84_tkeep(s_axis_scalar_84_tkeep),
        .s_axis_scalar_84_tstrb(s_axis_scalar_84_tstrb),
        .s_axis_scalar_84_tdata(s_axis_scalar_84_tdata),
        .s_axis_scalar_84_tready(s_axis_scalar_84_tready),
        .s_axis_scalar_85_aclk(s_axis_scalar_85_aclk),
        .s_axis_scalar_85_aresetn(s_axis_scalar_85_aresetn),
        .s_axis_scalar_85_tlast(s_axis_scalar_85_tlast),
        .s_axis_scalar_85_tvalid(s_axis_scalar_85_tvalid),
        .s_axis_scalar_85_tkeep(s_axis_scalar_85_tkeep),
        .s_axis_scalar_85_tstrb(s_axis_scalar_85_tstrb),
        .s_axis_scalar_85_tdata(s_axis_scalar_85_tdata),
        .s_axis_scalar_85_tready(s_axis_scalar_85_tready),
        .s_axis_scalar_86_aclk(s_axis_scalar_86_aclk),
        .s_axis_scalar_86_aresetn(s_axis_scalar_86_aresetn),
        .s_axis_scalar_86_tlast(s_axis_scalar_86_tlast),
        .s_axis_scalar_86_tvalid(s_axis_scalar_86_tvalid),
        .s_axis_scalar_86_tkeep(s_axis_scalar_86_tkeep),
        .s_axis_scalar_86_tstrb(s_axis_scalar_86_tstrb),
        .s_axis_scalar_86_tdata(s_axis_scalar_86_tdata),
        .s_axis_scalar_86_tready(s_axis_scalar_86_tready),
        .s_axis_scalar_87_aclk(s_axis_scalar_87_aclk),
        .s_axis_scalar_87_aresetn(s_axis_scalar_87_aresetn),
        .s_axis_scalar_87_tlast(s_axis_scalar_87_tlast),
        .s_axis_scalar_87_tvalid(s_axis_scalar_87_tvalid),
        .s_axis_scalar_87_tkeep(s_axis_scalar_87_tkeep),
        .s_axis_scalar_87_tstrb(s_axis_scalar_87_tstrb),
        .s_axis_scalar_87_tdata(s_axis_scalar_87_tdata),
        .s_axis_scalar_87_tready(s_axis_scalar_87_tready),
        .s_axis_scalar_88_aclk(s_axis_scalar_88_aclk),
        .s_axis_scalar_88_aresetn(s_axis_scalar_88_aresetn),
        .s_axis_scalar_88_tlast(s_axis_scalar_88_tlast),
        .s_axis_scalar_88_tvalid(s_axis_scalar_88_tvalid),
        .s_axis_scalar_88_tkeep(s_axis_scalar_88_tkeep),
        .s_axis_scalar_88_tstrb(s_axis_scalar_88_tstrb),
        .s_axis_scalar_88_tdata(s_axis_scalar_88_tdata),
        .s_axis_scalar_88_tready(s_axis_scalar_88_tready),
        .s_axis_scalar_89_aclk(s_axis_scalar_89_aclk),
        .s_axis_scalar_89_aresetn(s_axis_scalar_89_aresetn),
        .s_axis_scalar_89_tlast(s_axis_scalar_89_tlast),
        .s_axis_scalar_89_tvalid(s_axis_scalar_89_tvalid),
        .s_axis_scalar_89_tkeep(s_axis_scalar_89_tkeep),
        .s_axis_scalar_89_tstrb(s_axis_scalar_89_tstrb),
        .s_axis_scalar_89_tdata(s_axis_scalar_89_tdata),
        .s_axis_scalar_89_tready(s_axis_scalar_89_tready),
        .s_axis_scalar_90_aclk(s_axis_scalar_90_aclk),
        .s_axis_scalar_90_aresetn(s_axis_scalar_90_aresetn),
        .s_axis_scalar_90_tlast(s_axis_scalar_90_tlast),
        .s_axis_scalar_90_tvalid(s_axis_scalar_90_tvalid),
        .s_axis_scalar_90_tkeep(s_axis_scalar_90_tkeep),
        .s_axis_scalar_90_tstrb(s_axis_scalar_90_tstrb),
        .s_axis_scalar_90_tdata(s_axis_scalar_90_tdata),
        .s_axis_scalar_90_tready(s_axis_scalar_90_tready),
        .s_axis_scalar_91_aclk(s_axis_scalar_91_aclk),
        .s_axis_scalar_91_aresetn(s_axis_scalar_91_aresetn),
        .s_axis_scalar_91_tlast(s_axis_scalar_91_tlast),
        .s_axis_scalar_91_tvalid(s_axis_scalar_91_tvalid),
        .s_axis_scalar_91_tkeep(s_axis_scalar_91_tkeep),
        .s_axis_scalar_91_tstrb(s_axis_scalar_91_tstrb),
        .s_axis_scalar_91_tdata(s_axis_scalar_91_tdata),
        .s_axis_scalar_91_tready(s_axis_scalar_91_tready),
        .s_axis_scalar_92_aclk(s_axis_scalar_92_aclk),
        .s_axis_scalar_92_aresetn(s_axis_scalar_92_aresetn),
        .s_axis_scalar_92_tlast(s_axis_scalar_92_tlast),
        .s_axis_scalar_92_tvalid(s_axis_scalar_92_tvalid),
        .s_axis_scalar_92_tkeep(s_axis_scalar_92_tkeep),
        .s_axis_scalar_92_tstrb(s_axis_scalar_92_tstrb),
        .s_axis_scalar_92_tdata(s_axis_scalar_92_tdata),
        .s_axis_scalar_92_tready(s_axis_scalar_92_tready),
        .s_axis_scalar_93_aclk(s_axis_scalar_93_aclk),
        .s_axis_scalar_93_aresetn(s_axis_scalar_93_aresetn),
        .s_axis_scalar_93_tlast(s_axis_scalar_93_tlast),
        .s_axis_scalar_93_tvalid(s_axis_scalar_93_tvalid),
        .s_axis_scalar_93_tkeep(s_axis_scalar_93_tkeep),
        .s_axis_scalar_93_tstrb(s_axis_scalar_93_tstrb),
        .s_axis_scalar_93_tdata(s_axis_scalar_93_tdata),
        .s_axis_scalar_93_tready(s_axis_scalar_93_tready),
        .s_axis_scalar_94_aclk(s_axis_scalar_94_aclk),
        .s_axis_scalar_94_aresetn(s_axis_scalar_94_aresetn),
        .s_axis_scalar_94_tlast(s_axis_scalar_94_tlast),
        .s_axis_scalar_94_tvalid(s_axis_scalar_94_tvalid),
        .s_axis_scalar_94_tkeep(s_axis_scalar_94_tkeep),
        .s_axis_scalar_94_tstrb(s_axis_scalar_94_tstrb),
        .s_axis_scalar_94_tdata(s_axis_scalar_94_tdata),
        .s_axis_scalar_94_tready(s_axis_scalar_94_tready),
        .s_axis_scalar_95_aclk(s_axis_scalar_95_aclk),
        .s_axis_scalar_95_aresetn(s_axis_scalar_95_aresetn),
        .s_axis_scalar_95_tlast(s_axis_scalar_95_tlast),
        .s_axis_scalar_95_tvalid(s_axis_scalar_95_tvalid),
        .s_axis_scalar_95_tkeep(s_axis_scalar_95_tkeep),
        .s_axis_scalar_95_tstrb(s_axis_scalar_95_tstrb),
        .s_axis_scalar_95_tdata(s_axis_scalar_95_tdata),
        .s_axis_scalar_95_tready(s_axis_scalar_95_tready),
        .s_axis_scalar_96_aclk(s_axis_scalar_96_aclk),
        .s_axis_scalar_96_aresetn(s_axis_scalar_96_aresetn),
        .s_axis_scalar_96_tlast(s_axis_scalar_96_tlast),
        .s_axis_scalar_96_tvalid(s_axis_scalar_96_tvalid),
        .s_axis_scalar_96_tkeep(s_axis_scalar_96_tkeep),
        .s_axis_scalar_96_tstrb(s_axis_scalar_96_tstrb),
        .s_axis_scalar_96_tdata(s_axis_scalar_96_tdata),
        .s_axis_scalar_96_tready(s_axis_scalar_96_tready),
        .s_axis_scalar_97_aclk(s_axis_scalar_97_aclk),
        .s_axis_scalar_97_aresetn(s_axis_scalar_97_aresetn),
        .s_axis_scalar_97_tlast(s_axis_scalar_97_tlast),
        .s_axis_scalar_97_tvalid(s_axis_scalar_97_tvalid),
        .s_axis_scalar_97_tkeep(s_axis_scalar_97_tkeep),
        .s_axis_scalar_97_tstrb(s_axis_scalar_97_tstrb),
        .s_axis_scalar_97_tdata(s_axis_scalar_97_tdata),
        .s_axis_scalar_97_tready(s_axis_scalar_97_tready),
        .s_axis_scalar_98_aclk(s_axis_scalar_98_aclk),
        .s_axis_scalar_98_aresetn(s_axis_scalar_98_aresetn),
        .s_axis_scalar_98_tlast(s_axis_scalar_98_tlast),
        .s_axis_scalar_98_tvalid(s_axis_scalar_98_tvalid),
        .s_axis_scalar_98_tkeep(s_axis_scalar_98_tkeep),
        .s_axis_scalar_98_tstrb(s_axis_scalar_98_tstrb),
        .s_axis_scalar_98_tdata(s_axis_scalar_98_tdata),
        .s_axis_scalar_98_tready(s_axis_scalar_98_tready),
        .s_axis_scalar_99_aclk(s_axis_scalar_99_aclk),
        .s_axis_scalar_99_aresetn(s_axis_scalar_99_aresetn),
        .s_axis_scalar_99_tlast(s_axis_scalar_99_tlast),
        .s_axis_scalar_99_tvalid(s_axis_scalar_99_tvalid),
        .s_axis_scalar_99_tkeep(s_axis_scalar_99_tkeep),
        .s_axis_scalar_99_tstrb(s_axis_scalar_99_tstrb),
        .s_axis_scalar_99_tdata(s_axis_scalar_99_tdata),
        .s_axis_scalar_99_tready(s_axis_scalar_99_tready),
        .s_axis_scalar_100_aclk(s_axis_scalar_100_aclk),
        .s_axis_scalar_100_aresetn(s_axis_scalar_100_aresetn),
        .s_axis_scalar_100_tlast(s_axis_scalar_100_tlast),
        .s_axis_scalar_100_tvalid(s_axis_scalar_100_tvalid),
        .s_axis_scalar_100_tkeep(s_axis_scalar_100_tkeep),
        .s_axis_scalar_100_tstrb(s_axis_scalar_100_tstrb),
        .s_axis_scalar_100_tdata(s_axis_scalar_100_tdata),
        .s_axis_scalar_100_tready(s_axis_scalar_100_tready),
        .s_axis_scalar_101_aclk(s_axis_scalar_101_aclk),
        .s_axis_scalar_101_aresetn(s_axis_scalar_101_aresetn),
        .s_axis_scalar_101_tlast(s_axis_scalar_101_tlast),
        .s_axis_scalar_101_tvalid(s_axis_scalar_101_tvalid),
        .s_axis_scalar_101_tkeep(s_axis_scalar_101_tkeep),
        .s_axis_scalar_101_tstrb(s_axis_scalar_101_tstrb),
        .s_axis_scalar_101_tdata(s_axis_scalar_101_tdata),
        .s_axis_scalar_101_tready(s_axis_scalar_101_tready),
        .s_axis_scalar_102_aclk(s_axis_scalar_102_aclk),
        .s_axis_scalar_102_aresetn(s_axis_scalar_102_aresetn),
        .s_axis_scalar_102_tlast(s_axis_scalar_102_tlast),
        .s_axis_scalar_102_tvalid(s_axis_scalar_102_tvalid),
        .s_axis_scalar_102_tkeep(s_axis_scalar_102_tkeep),
        .s_axis_scalar_102_tstrb(s_axis_scalar_102_tstrb),
        .s_axis_scalar_102_tdata(s_axis_scalar_102_tdata),
        .s_axis_scalar_102_tready(s_axis_scalar_102_tready),
        .s_axis_scalar_103_aclk(s_axis_scalar_103_aclk),
        .s_axis_scalar_103_aresetn(s_axis_scalar_103_aresetn),
        .s_axis_scalar_103_tlast(s_axis_scalar_103_tlast),
        .s_axis_scalar_103_tvalid(s_axis_scalar_103_tvalid),
        .s_axis_scalar_103_tkeep(s_axis_scalar_103_tkeep),
        .s_axis_scalar_103_tstrb(s_axis_scalar_103_tstrb),
        .s_axis_scalar_103_tdata(s_axis_scalar_103_tdata),
        .s_axis_scalar_103_tready(s_axis_scalar_103_tready),
        .s_axis_scalar_104_aclk(s_axis_scalar_104_aclk),
        .s_axis_scalar_104_aresetn(s_axis_scalar_104_aresetn),
        .s_axis_scalar_104_tlast(s_axis_scalar_104_tlast),
        .s_axis_scalar_104_tvalid(s_axis_scalar_104_tvalid),
        .s_axis_scalar_104_tkeep(s_axis_scalar_104_tkeep),
        .s_axis_scalar_104_tstrb(s_axis_scalar_104_tstrb),
        .s_axis_scalar_104_tdata(s_axis_scalar_104_tdata),
        .s_axis_scalar_104_tready(s_axis_scalar_104_tready),
        .s_axis_scalar_105_aclk(s_axis_scalar_105_aclk),
        .s_axis_scalar_105_aresetn(s_axis_scalar_105_aresetn),
        .s_axis_scalar_105_tlast(s_axis_scalar_105_tlast),
        .s_axis_scalar_105_tvalid(s_axis_scalar_105_tvalid),
        .s_axis_scalar_105_tkeep(s_axis_scalar_105_tkeep),
        .s_axis_scalar_105_tstrb(s_axis_scalar_105_tstrb),
        .s_axis_scalar_105_tdata(s_axis_scalar_105_tdata),
        .s_axis_scalar_105_tready(s_axis_scalar_105_tready),
        .s_axis_scalar_106_aclk(s_axis_scalar_106_aclk),
        .s_axis_scalar_106_aresetn(s_axis_scalar_106_aresetn),
        .s_axis_scalar_106_tlast(s_axis_scalar_106_tlast),
        .s_axis_scalar_106_tvalid(s_axis_scalar_106_tvalid),
        .s_axis_scalar_106_tkeep(s_axis_scalar_106_tkeep),
        .s_axis_scalar_106_tstrb(s_axis_scalar_106_tstrb),
        .s_axis_scalar_106_tdata(s_axis_scalar_106_tdata),
        .s_axis_scalar_106_tready(s_axis_scalar_106_tready),
        .s_axis_scalar_107_aclk(s_axis_scalar_107_aclk),
        .s_axis_scalar_107_aresetn(s_axis_scalar_107_aresetn),
        .s_axis_scalar_107_tlast(s_axis_scalar_107_tlast),
        .s_axis_scalar_107_tvalid(s_axis_scalar_107_tvalid),
        .s_axis_scalar_107_tkeep(s_axis_scalar_107_tkeep),
        .s_axis_scalar_107_tstrb(s_axis_scalar_107_tstrb),
        .s_axis_scalar_107_tdata(s_axis_scalar_107_tdata),
        .s_axis_scalar_107_tready(s_axis_scalar_107_tready),
        .s_axis_scalar_108_aclk(s_axis_scalar_108_aclk),
        .s_axis_scalar_108_aresetn(s_axis_scalar_108_aresetn),
        .s_axis_scalar_108_tlast(s_axis_scalar_108_tlast),
        .s_axis_scalar_108_tvalid(s_axis_scalar_108_tvalid),
        .s_axis_scalar_108_tkeep(s_axis_scalar_108_tkeep),
        .s_axis_scalar_108_tstrb(s_axis_scalar_108_tstrb),
        .s_axis_scalar_108_tdata(s_axis_scalar_108_tdata),
        .s_axis_scalar_108_tready(s_axis_scalar_108_tready),
        .s_axis_scalar_109_aclk(s_axis_scalar_109_aclk),
        .s_axis_scalar_109_aresetn(s_axis_scalar_109_aresetn),
        .s_axis_scalar_109_tlast(s_axis_scalar_109_tlast),
        .s_axis_scalar_109_tvalid(s_axis_scalar_109_tvalid),
        .s_axis_scalar_109_tkeep(s_axis_scalar_109_tkeep),
        .s_axis_scalar_109_tstrb(s_axis_scalar_109_tstrb),
        .s_axis_scalar_109_tdata(s_axis_scalar_109_tdata),
        .s_axis_scalar_109_tready(s_axis_scalar_109_tready),
        .s_axis_scalar_110_aclk(s_axis_scalar_110_aclk),
        .s_axis_scalar_110_aresetn(s_axis_scalar_110_aresetn),
        .s_axis_scalar_110_tlast(s_axis_scalar_110_tlast),
        .s_axis_scalar_110_tvalid(s_axis_scalar_110_tvalid),
        .s_axis_scalar_110_tkeep(s_axis_scalar_110_tkeep),
        .s_axis_scalar_110_tstrb(s_axis_scalar_110_tstrb),
        .s_axis_scalar_110_tdata(s_axis_scalar_110_tdata),
        .s_axis_scalar_110_tready(s_axis_scalar_110_tready),
        .s_axis_scalar_111_aclk(s_axis_scalar_111_aclk),
        .s_axis_scalar_111_aresetn(s_axis_scalar_111_aresetn),
        .s_axis_scalar_111_tlast(s_axis_scalar_111_tlast),
        .s_axis_scalar_111_tvalid(s_axis_scalar_111_tvalid),
        .s_axis_scalar_111_tkeep(s_axis_scalar_111_tkeep),
        .s_axis_scalar_111_tstrb(s_axis_scalar_111_tstrb),
        .s_axis_scalar_111_tdata(s_axis_scalar_111_tdata),
        .s_axis_scalar_111_tready(s_axis_scalar_111_tready),
        .s_axis_scalar_112_aclk(s_axis_scalar_112_aclk),
        .s_axis_scalar_112_aresetn(s_axis_scalar_112_aresetn),
        .s_axis_scalar_112_tlast(s_axis_scalar_112_tlast),
        .s_axis_scalar_112_tvalid(s_axis_scalar_112_tvalid),
        .s_axis_scalar_112_tkeep(s_axis_scalar_112_tkeep),
        .s_axis_scalar_112_tstrb(s_axis_scalar_112_tstrb),
        .s_axis_scalar_112_tdata(s_axis_scalar_112_tdata),
        .s_axis_scalar_112_tready(s_axis_scalar_112_tready),
        .s_axis_scalar_113_aclk(s_axis_scalar_113_aclk),
        .s_axis_scalar_113_aresetn(s_axis_scalar_113_aresetn),
        .s_axis_scalar_113_tlast(s_axis_scalar_113_tlast),
        .s_axis_scalar_113_tvalid(s_axis_scalar_113_tvalid),
        .s_axis_scalar_113_tkeep(s_axis_scalar_113_tkeep),
        .s_axis_scalar_113_tstrb(s_axis_scalar_113_tstrb),
        .s_axis_scalar_113_tdata(s_axis_scalar_113_tdata),
        .s_axis_scalar_113_tready(s_axis_scalar_113_tready),
        .s_axis_scalar_114_aclk(s_axis_scalar_114_aclk),
        .s_axis_scalar_114_aresetn(s_axis_scalar_114_aresetn),
        .s_axis_scalar_114_tlast(s_axis_scalar_114_tlast),
        .s_axis_scalar_114_tvalid(s_axis_scalar_114_tvalid),
        .s_axis_scalar_114_tkeep(s_axis_scalar_114_tkeep),
        .s_axis_scalar_114_tstrb(s_axis_scalar_114_tstrb),
        .s_axis_scalar_114_tdata(s_axis_scalar_114_tdata),
        .s_axis_scalar_114_tready(s_axis_scalar_114_tready),
        .s_axis_scalar_115_aclk(s_axis_scalar_115_aclk),
        .s_axis_scalar_115_aresetn(s_axis_scalar_115_aresetn),
        .s_axis_scalar_115_tlast(s_axis_scalar_115_tlast),
        .s_axis_scalar_115_tvalid(s_axis_scalar_115_tvalid),
        .s_axis_scalar_115_tkeep(s_axis_scalar_115_tkeep),
        .s_axis_scalar_115_tstrb(s_axis_scalar_115_tstrb),
        .s_axis_scalar_115_tdata(s_axis_scalar_115_tdata),
        .s_axis_scalar_115_tready(s_axis_scalar_115_tready),
        .s_axis_scalar_116_aclk(s_axis_scalar_116_aclk),
        .s_axis_scalar_116_aresetn(s_axis_scalar_116_aresetn),
        .s_axis_scalar_116_tlast(s_axis_scalar_116_tlast),
        .s_axis_scalar_116_tvalid(s_axis_scalar_116_tvalid),
        .s_axis_scalar_116_tkeep(s_axis_scalar_116_tkeep),
        .s_axis_scalar_116_tstrb(s_axis_scalar_116_tstrb),
        .s_axis_scalar_116_tdata(s_axis_scalar_116_tdata),
        .s_axis_scalar_116_tready(s_axis_scalar_116_tready),
        .s_axis_scalar_117_aclk(s_axis_scalar_117_aclk),
        .s_axis_scalar_117_aresetn(s_axis_scalar_117_aresetn),
        .s_axis_scalar_117_tlast(s_axis_scalar_117_tlast),
        .s_axis_scalar_117_tvalid(s_axis_scalar_117_tvalid),
        .s_axis_scalar_117_tkeep(s_axis_scalar_117_tkeep),
        .s_axis_scalar_117_tstrb(s_axis_scalar_117_tstrb),
        .s_axis_scalar_117_tdata(s_axis_scalar_117_tdata),
        .s_axis_scalar_117_tready(s_axis_scalar_117_tready),
        .s_axis_scalar_118_aclk(s_axis_scalar_118_aclk),
        .s_axis_scalar_118_aresetn(s_axis_scalar_118_aresetn),
        .s_axis_scalar_118_tlast(s_axis_scalar_118_tlast),
        .s_axis_scalar_118_tvalid(s_axis_scalar_118_tvalid),
        .s_axis_scalar_118_tkeep(s_axis_scalar_118_tkeep),
        .s_axis_scalar_118_tstrb(s_axis_scalar_118_tstrb),
        .s_axis_scalar_118_tdata(s_axis_scalar_118_tdata),
        .s_axis_scalar_118_tready(s_axis_scalar_118_tready),
        .s_axis_scalar_119_aclk(s_axis_scalar_119_aclk),
        .s_axis_scalar_119_aresetn(s_axis_scalar_119_aresetn),
        .s_axis_scalar_119_tlast(s_axis_scalar_119_tlast),
        .s_axis_scalar_119_tvalid(s_axis_scalar_119_tvalid),
        .s_axis_scalar_119_tkeep(s_axis_scalar_119_tkeep),
        .s_axis_scalar_119_tstrb(s_axis_scalar_119_tstrb),
        .s_axis_scalar_119_tdata(s_axis_scalar_119_tdata),
        .s_axis_scalar_119_tready(s_axis_scalar_119_tready),
        .s_axis_scalar_120_aclk(s_axis_scalar_120_aclk),
        .s_axis_scalar_120_aresetn(s_axis_scalar_120_aresetn),
        .s_axis_scalar_120_tlast(s_axis_scalar_120_tlast),
        .s_axis_scalar_120_tvalid(s_axis_scalar_120_tvalid),
        .s_axis_scalar_120_tkeep(s_axis_scalar_120_tkeep),
        .s_axis_scalar_120_tstrb(s_axis_scalar_120_tstrb),
        .s_axis_scalar_120_tdata(s_axis_scalar_120_tdata),
        .s_axis_scalar_120_tready(s_axis_scalar_120_tready),
        .s_axis_scalar_121_aclk(s_axis_scalar_121_aclk),
        .s_axis_scalar_121_aresetn(s_axis_scalar_121_aresetn),
        .s_axis_scalar_121_tlast(s_axis_scalar_121_tlast),
        .s_axis_scalar_121_tvalid(s_axis_scalar_121_tvalid),
        .s_axis_scalar_121_tkeep(s_axis_scalar_121_tkeep),
        .s_axis_scalar_121_tstrb(s_axis_scalar_121_tstrb),
        .s_axis_scalar_121_tdata(s_axis_scalar_121_tdata),
        .s_axis_scalar_121_tready(s_axis_scalar_121_tready),
        .s_axis_scalar_122_aclk(s_axis_scalar_122_aclk),
        .s_axis_scalar_122_aresetn(s_axis_scalar_122_aresetn),
        .s_axis_scalar_122_tlast(s_axis_scalar_122_tlast),
        .s_axis_scalar_122_tvalid(s_axis_scalar_122_tvalid),
        .s_axis_scalar_122_tkeep(s_axis_scalar_122_tkeep),
        .s_axis_scalar_122_tstrb(s_axis_scalar_122_tstrb),
        .s_axis_scalar_122_tdata(s_axis_scalar_122_tdata),
        .s_axis_scalar_122_tready(s_axis_scalar_122_tready),
        .s_axis_scalar_123_aclk(s_axis_scalar_123_aclk),
        .s_axis_scalar_123_aresetn(s_axis_scalar_123_aresetn),
        .s_axis_scalar_123_tlast(s_axis_scalar_123_tlast),
        .s_axis_scalar_123_tvalid(s_axis_scalar_123_tvalid),
        .s_axis_scalar_123_tkeep(s_axis_scalar_123_tkeep),
        .s_axis_scalar_123_tstrb(s_axis_scalar_123_tstrb),
        .s_axis_scalar_123_tdata(s_axis_scalar_123_tdata),
        .s_axis_scalar_123_tready(s_axis_scalar_123_tready),
        .s_axis_scalar_124_aclk(s_axis_scalar_124_aclk),
        .s_axis_scalar_124_aresetn(s_axis_scalar_124_aresetn),
        .s_axis_scalar_124_tlast(s_axis_scalar_124_tlast),
        .s_axis_scalar_124_tvalid(s_axis_scalar_124_tvalid),
        .s_axis_scalar_124_tkeep(s_axis_scalar_124_tkeep),
        .s_axis_scalar_124_tstrb(s_axis_scalar_124_tstrb),
        .s_axis_scalar_124_tdata(s_axis_scalar_124_tdata),
        .s_axis_scalar_124_tready(s_axis_scalar_124_tready),
        .s_axis_scalar_125_aclk(s_axis_scalar_125_aclk),
        .s_axis_scalar_125_aresetn(s_axis_scalar_125_aresetn),
        .s_axis_scalar_125_tlast(s_axis_scalar_125_tlast),
        .s_axis_scalar_125_tvalid(s_axis_scalar_125_tvalid),
        .s_axis_scalar_125_tkeep(s_axis_scalar_125_tkeep),
        .s_axis_scalar_125_tstrb(s_axis_scalar_125_tstrb),
        .s_axis_scalar_125_tdata(s_axis_scalar_125_tdata),
        .s_axis_scalar_125_tready(s_axis_scalar_125_tready),
        .s_axis_scalar_126_aclk(s_axis_scalar_126_aclk),
        .s_axis_scalar_126_aresetn(s_axis_scalar_126_aresetn),
        .s_axis_scalar_126_tlast(s_axis_scalar_126_tlast),
        .s_axis_scalar_126_tvalid(s_axis_scalar_126_tvalid),
        .s_axis_scalar_126_tkeep(s_axis_scalar_126_tkeep),
        .s_axis_scalar_126_tstrb(s_axis_scalar_126_tstrb),
        .s_axis_scalar_126_tdata(s_axis_scalar_126_tdata),
        .s_axis_scalar_126_tready(s_axis_scalar_126_tready),
        .s_axis_scalar_127_aclk(s_axis_scalar_127_aclk),
        .s_axis_scalar_127_aresetn(s_axis_scalar_127_aresetn),
        .s_axis_scalar_127_tlast(s_axis_scalar_127_tlast),
        .s_axis_scalar_127_tvalid(s_axis_scalar_127_tvalid),
        .s_axis_scalar_127_tkeep(s_axis_scalar_127_tkeep),
        .s_axis_scalar_127_tstrb(s_axis_scalar_127_tstrb),
        .s_axis_scalar_127_tdata(s_axis_scalar_127_tdata),
        .s_axis_scalar_127_tready(s_axis_scalar_127_tready),
        //.scalar ports
        .outscalar0(ap_oscalar_0_din),
        .outscalar1(ap_oscalar_1_din),
        .outscalar2(ap_oscalar_2_din),
        .outscalar3(ap_oscalar_3_din),
        .outscalar4(ap_oscalar_4_din),
        .outscalar5(ap_oscalar_5_din),
        .outscalar6(ap_oscalar_6_din),
        .outscalar7(ap_oscalar_7_din),
        .outscalar8(ap_oscalar_8_din),
        .outscalar9(ap_oscalar_9_din),
        .outscalar10(ap_oscalar_10_din),
        .outscalar11(ap_oscalar_11_din),
        .outscalar12(ap_oscalar_12_din),
        .outscalar13(ap_oscalar_13_din),
        .outscalar14(ap_oscalar_14_din),
        .outscalar15(ap_oscalar_15_din),
        .outscalar16(ap_oscalar_16_din),
        .outscalar17(ap_oscalar_17_din),
        .outscalar18(ap_oscalar_18_din),
        .outscalar19(ap_oscalar_19_din),
        .outscalar20(ap_oscalar_20_din),
        .outscalar21(ap_oscalar_21_din),
        .outscalar22(ap_oscalar_22_din),
        .outscalar23(ap_oscalar_23_din),
        .outscalar24(ap_oscalar_24_din),
        .outscalar25(ap_oscalar_25_din),
        .outscalar26(ap_oscalar_26_din),
        .outscalar27(ap_oscalar_27_din),
        .outscalar28(ap_oscalar_28_din),
        .outscalar29(ap_oscalar_29_din),
        .outscalar30(ap_oscalar_30_din),
        .outscalar31(ap_oscalar_31_din),
        .outscalar32(ap_oscalar_32_din),
        .outscalar33(ap_oscalar_33_din),
        .outscalar34(ap_oscalar_34_din),
        .outscalar35(ap_oscalar_35_din),
        .outscalar36(ap_oscalar_36_din),
        .outscalar37(ap_oscalar_37_din),
        .outscalar38(ap_oscalar_38_din),
        .outscalar39(ap_oscalar_39_din),
        .outscalar40(ap_oscalar_40_din),
        .outscalar41(ap_oscalar_41_din),
        .outscalar42(ap_oscalar_42_din),
        .outscalar43(ap_oscalar_43_din),
        .outscalar44(ap_oscalar_44_din),
        .outscalar45(ap_oscalar_45_din),
        .outscalar46(ap_oscalar_46_din),
        .outscalar47(ap_oscalar_47_din),
        .outscalar48(ap_oscalar_48_din),
        .outscalar49(ap_oscalar_49_din),
        .outscalar50(ap_oscalar_50_din),
        .outscalar51(ap_oscalar_51_din),
        .outscalar52(ap_oscalar_52_din),
        .outscalar53(ap_oscalar_53_din),
        .outscalar54(ap_oscalar_54_din),
        .outscalar55(ap_oscalar_55_din),
        .outscalar56(ap_oscalar_56_din),
        .outscalar57(ap_oscalar_57_din),
        .outscalar58(ap_oscalar_58_din),
        .outscalar59(ap_oscalar_59_din),
        .outscalar60(ap_oscalar_60_din),
        .outscalar61(ap_oscalar_61_din),
        .outscalar62(ap_oscalar_62_din),
        .outscalar63(ap_oscalar_63_din),
        .outscalar64(ap_oscalar_64_din),
        .outscalar65(ap_oscalar_65_din),
        .outscalar66(ap_oscalar_66_din),
        .outscalar67(ap_oscalar_67_din),
        .outscalar68(ap_oscalar_68_din),
        .outscalar69(ap_oscalar_69_din),
        .outscalar70(ap_oscalar_70_din),
        .outscalar71(ap_oscalar_71_din),
        .outscalar72(ap_oscalar_72_din),
        .outscalar73(ap_oscalar_73_din),
        .outscalar74(ap_oscalar_74_din),
        .outscalar75(ap_oscalar_75_din),
        .outscalar76(ap_oscalar_76_din),
        .outscalar77(ap_oscalar_77_din),
        .outscalar78(ap_oscalar_78_din),
        .outscalar79(ap_oscalar_79_din),
        .outscalar80(ap_oscalar_80_din),
        .outscalar81(ap_oscalar_81_din),
        .outscalar82(ap_oscalar_82_din),
        .outscalar83(ap_oscalar_83_din),
        .outscalar84(ap_oscalar_84_din),
        .outscalar85(ap_oscalar_85_din),
        .outscalar86(ap_oscalar_86_din),
        .outscalar87(ap_oscalar_87_din),
        .outscalar88(ap_oscalar_88_din),
        .outscalar89(ap_oscalar_89_din),
        .outscalar90(ap_oscalar_90_din),
        .outscalar91(ap_oscalar_91_din),
        .outscalar92(ap_oscalar_92_din),
        .outscalar93(ap_oscalar_93_din),
        .outscalar94(ap_oscalar_94_din),
        .outscalar95(ap_oscalar_95_din),
        .outscalar96(ap_oscalar_96_din),
        .outscalar97(ap_oscalar_97_din),
        .outscalar98(ap_oscalar_98_din),
        .outscalar99(ap_oscalar_99_din),
        .outscalar100(ap_oscalar_100_din),
        .outscalar101(ap_oscalar_101_din),
        .outscalar102(ap_oscalar_102_din),
        .outscalar103(ap_oscalar_103_din),
        .outscalar104(ap_oscalar_104_din),
        .outscalar105(ap_oscalar_105_din),
        .outscalar106(ap_oscalar_106_din),
        .outscalar107(ap_oscalar_107_din),
        .outscalar108(ap_oscalar_108_din),
        .outscalar109(ap_oscalar_109_din),
        .outscalar110(ap_oscalar_110_din),
        .outscalar111(ap_oscalar_111_din),
        .outscalar112(ap_oscalar_112_din),
        .outscalar113(ap_oscalar_113_din),
        .outscalar114(ap_oscalar_114_din),
        .outscalar115(ap_oscalar_115_din),
        .outscalar116(ap_oscalar_116_din),
        .outscalar117(ap_oscalar_117_din),
        .outscalar118(ap_oscalar_118_din),
        .outscalar119(ap_oscalar_119_din),
        .outscalar120(ap_oscalar_120_din),
        .outscalar121(ap_oscalar_121_din),
        .outscalar122(ap_oscalar_122_din),
        .outscalar123(ap_oscalar_123_din),
        .outscalar124(ap_oscalar_124_din),
        .outscalar125(ap_oscalar_125_din),
        .outscalar126(ap_oscalar_126_din),
        .outscalar127(ap_oscalar_127_din),
        //.scalar valid ports
        .outscalar0_vld(ap_oscalar_0_vld),
        .outscalar1_vld(ap_oscalar_1_vld),
        .outscalar2_vld(ap_oscalar_2_vld),
        .outscalar3_vld(ap_oscalar_3_vld),
        .outscalar4_vld(ap_oscalar_4_vld),
        .outscalar5_vld(ap_oscalar_5_vld),
        .outscalar6_vld(ap_oscalar_6_vld),
        .outscalar7_vld(ap_oscalar_7_vld),
        .outscalar8_vld(ap_oscalar_8_vld),
        .outscalar9_vld(ap_oscalar_9_vld),
        .outscalar10_vld(ap_oscalar_10_vld),
        .outscalar11_vld(ap_oscalar_11_vld),
        .outscalar12_vld(ap_oscalar_12_vld),
        .outscalar13_vld(ap_oscalar_13_vld),
        .outscalar14_vld(ap_oscalar_14_vld),
        .outscalar15_vld(ap_oscalar_15_vld),
        .outscalar16_vld(ap_oscalar_16_vld),
        .outscalar17_vld(ap_oscalar_17_vld),
        .outscalar18_vld(ap_oscalar_18_vld),
        .outscalar19_vld(ap_oscalar_19_vld),
        .outscalar20_vld(ap_oscalar_20_vld),
        .outscalar21_vld(ap_oscalar_21_vld),
        .outscalar22_vld(ap_oscalar_22_vld),
        .outscalar23_vld(ap_oscalar_23_vld),
        .outscalar24_vld(ap_oscalar_24_vld),
        .outscalar25_vld(ap_oscalar_25_vld),
        .outscalar26_vld(ap_oscalar_26_vld),
        .outscalar27_vld(ap_oscalar_27_vld),
        .outscalar28_vld(ap_oscalar_28_vld),
        .outscalar29_vld(ap_oscalar_29_vld),
        .outscalar30_vld(ap_oscalar_30_vld),
        .outscalar31_vld(ap_oscalar_31_vld),
        .outscalar32_vld(ap_oscalar_32_vld),
        .outscalar33_vld(ap_oscalar_33_vld),
        .outscalar34_vld(ap_oscalar_34_vld),
        .outscalar35_vld(ap_oscalar_35_vld),
        .outscalar36_vld(ap_oscalar_36_vld),
        .outscalar37_vld(ap_oscalar_37_vld),
        .outscalar38_vld(ap_oscalar_38_vld),
        .outscalar39_vld(ap_oscalar_39_vld),
        .outscalar40_vld(ap_oscalar_40_vld),
        .outscalar41_vld(ap_oscalar_41_vld),
        .outscalar42_vld(ap_oscalar_42_vld),
        .outscalar43_vld(ap_oscalar_43_vld),
        .outscalar44_vld(ap_oscalar_44_vld),
        .outscalar45_vld(ap_oscalar_45_vld),
        .outscalar46_vld(ap_oscalar_46_vld),
        .outscalar47_vld(ap_oscalar_47_vld),
        .outscalar48_vld(ap_oscalar_48_vld),
        .outscalar49_vld(ap_oscalar_49_vld),
        .outscalar50_vld(ap_oscalar_50_vld),
        .outscalar51_vld(ap_oscalar_51_vld),
        .outscalar52_vld(ap_oscalar_52_vld),
        .outscalar53_vld(ap_oscalar_53_vld),
        .outscalar54_vld(ap_oscalar_54_vld),
        .outscalar55_vld(ap_oscalar_55_vld),
        .outscalar56_vld(ap_oscalar_56_vld),
        .outscalar57_vld(ap_oscalar_57_vld),
        .outscalar58_vld(ap_oscalar_58_vld),
        .outscalar59_vld(ap_oscalar_59_vld),
        .outscalar60_vld(ap_oscalar_60_vld),
        .outscalar61_vld(ap_oscalar_61_vld),
        .outscalar62_vld(ap_oscalar_62_vld),
        .outscalar63_vld(ap_oscalar_63_vld),
        .outscalar64_vld(ap_oscalar_64_vld),
        .outscalar65_vld(ap_oscalar_65_vld),
        .outscalar66_vld(ap_oscalar_66_vld),
        .outscalar67_vld(ap_oscalar_67_vld),
        .outscalar68_vld(ap_oscalar_68_vld),
        .outscalar69_vld(ap_oscalar_69_vld),
        .outscalar70_vld(ap_oscalar_70_vld),
        .outscalar71_vld(ap_oscalar_71_vld),
        .outscalar72_vld(ap_oscalar_72_vld),
        .outscalar73_vld(ap_oscalar_73_vld),
        .outscalar74_vld(ap_oscalar_74_vld),
        .outscalar75_vld(ap_oscalar_75_vld),
        .outscalar76_vld(ap_oscalar_76_vld),
        .outscalar77_vld(ap_oscalar_77_vld),
        .outscalar78_vld(ap_oscalar_78_vld),
        .outscalar79_vld(ap_oscalar_79_vld),
        .outscalar80_vld(ap_oscalar_80_vld),
        .outscalar81_vld(ap_oscalar_81_vld),
        .outscalar82_vld(ap_oscalar_82_vld),
        .outscalar83_vld(ap_oscalar_83_vld),
        .outscalar84_vld(ap_oscalar_84_vld),
        .outscalar85_vld(ap_oscalar_85_vld),
        .outscalar86_vld(ap_oscalar_86_vld),
        .outscalar87_vld(ap_oscalar_87_vld),
        .outscalar88_vld(ap_oscalar_88_vld),
        .outscalar89_vld(ap_oscalar_89_vld),
        .outscalar90_vld(ap_oscalar_90_vld),
        .outscalar91_vld(ap_oscalar_91_vld),
        .outscalar92_vld(ap_oscalar_92_vld),
        .outscalar93_vld(ap_oscalar_93_vld),
        .outscalar94_vld(ap_oscalar_94_vld),
        .outscalar95_vld(ap_oscalar_95_vld),
        .outscalar96_vld(ap_oscalar_96_vld),
        .outscalar97_vld(ap_oscalar_97_vld),
        .outscalar98_vld(ap_oscalar_98_vld),
        .outscalar99_vld(ap_oscalar_99_vld),
        .outscalar100_vld(ap_oscalar_100_vld),
        .outscalar101_vld(ap_oscalar_101_vld),
        .outscalar102_vld(ap_oscalar_102_vld),
        .outscalar103_vld(ap_oscalar_103_vld),
        .outscalar104_vld(ap_oscalar_104_vld),
        .outscalar105_vld(ap_oscalar_105_vld),
        .outscalar106_vld(ap_oscalar_106_vld),
        .outscalar107_vld(ap_oscalar_107_vld),
        .outscalar108_vld(ap_oscalar_108_vld),
        .outscalar109_vld(ap_oscalar_109_vld),
        .outscalar110_vld(ap_oscalar_110_vld),
        .outscalar111_vld(ap_oscalar_111_vld),
        .outscalar112_vld(ap_oscalar_112_vld),
        .outscalar113_vld(ap_oscalar_113_vld),
        .outscalar114_vld(ap_oscalar_114_vld),
        .outscalar115_vld(ap_oscalar_115_vld),
        .outscalar116_vld(ap_oscalar_116_vld),
        .outscalar117_vld(ap_oscalar_117_vld),
        .outscalar118_vld(ap_oscalar_118_vld),
        .outscalar119_vld(ap_oscalar_119_vld),
        .outscalar120_vld(ap_oscalar_120_vld),
        .outscalar121_vld(ap_oscalar_121_vld),
        .outscalar122_vld(ap_oscalar_122_vld),
        .outscalar123_vld(ap_oscalar_123_vld),
        .outscalar124_vld(ap_oscalar_124_vld),
        .outscalar125_vld(ap_oscalar_125_vld),
        .outscalar126_vld(ap_oscalar_126_vld),
        .outscalar127_vld(ap_oscalar_127_vld),
        .m_axis_scalar_0_aclk(m_axis_scalar_0_aclk),
        .m_axis_scalar_0_aresetn(m_axis_scalar_0_aresetn),
        .m_axis_scalar_0_tlast(m_axis_scalar_0_tlast),
        .m_axis_scalar_0_tvalid(m_axis_scalar_0_tvalid),
        .m_axis_scalar_0_tkeep(m_axis_scalar_0_tkeep),
        .m_axis_scalar_0_tstrb(m_axis_scalar_0_tstrb),
        .m_axis_scalar_0_tdata(m_axis_scalar_0_tdata),
        .m_axis_scalar_0_tready(m_axis_scalar_0_tready),
        .m_axis_scalar_1_aclk(m_axis_scalar_1_aclk),
        .m_axis_scalar_1_aresetn(m_axis_scalar_1_aresetn),
        .m_axis_scalar_1_tlast(m_axis_scalar_1_tlast),
        .m_axis_scalar_1_tvalid(m_axis_scalar_1_tvalid),
        .m_axis_scalar_1_tkeep(m_axis_scalar_1_tkeep),
        .m_axis_scalar_1_tstrb(m_axis_scalar_1_tstrb),
        .m_axis_scalar_1_tdata(m_axis_scalar_1_tdata),
        .m_axis_scalar_1_tready(m_axis_scalar_1_tready),
        .m_axis_scalar_2_aclk(m_axis_scalar_2_aclk),
        .m_axis_scalar_2_aresetn(m_axis_scalar_2_aresetn),
        .m_axis_scalar_2_tlast(m_axis_scalar_2_tlast),
        .m_axis_scalar_2_tvalid(m_axis_scalar_2_tvalid),
        .m_axis_scalar_2_tkeep(m_axis_scalar_2_tkeep),
        .m_axis_scalar_2_tstrb(m_axis_scalar_2_tstrb),
        .m_axis_scalar_2_tdata(m_axis_scalar_2_tdata),
        .m_axis_scalar_2_tready(m_axis_scalar_2_tready),
        .m_axis_scalar_3_aclk(m_axis_scalar_3_aclk),
        .m_axis_scalar_3_aresetn(m_axis_scalar_3_aresetn),
        .m_axis_scalar_3_tlast(m_axis_scalar_3_tlast),
        .m_axis_scalar_3_tvalid(m_axis_scalar_3_tvalid),
        .m_axis_scalar_3_tkeep(m_axis_scalar_3_tkeep),
        .m_axis_scalar_3_tstrb(m_axis_scalar_3_tstrb),
        .m_axis_scalar_3_tdata(m_axis_scalar_3_tdata),
        .m_axis_scalar_3_tready(m_axis_scalar_3_tready),
        .m_axis_scalar_4_aclk(m_axis_scalar_4_aclk),
        .m_axis_scalar_4_aresetn(m_axis_scalar_4_aresetn),
        .m_axis_scalar_4_tlast(m_axis_scalar_4_tlast),
        .m_axis_scalar_4_tvalid(m_axis_scalar_4_tvalid),
        .m_axis_scalar_4_tkeep(m_axis_scalar_4_tkeep),
        .m_axis_scalar_4_tstrb(m_axis_scalar_4_tstrb),
        .m_axis_scalar_4_tdata(m_axis_scalar_4_tdata),
        .m_axis_scalar_4_tready(m_axis_scalar_4_tready),
        .m_axis_scalar_5_aclk(m_axis_scalar_5_aclk),
        .m_axis_scalar_5_aresetn(m_axis_scalar_5_aresetn),
        .m_axis_scalar_5_tlast(m_axis_scalar_5_tlast),
        .m_axis_scalar_5_tvalid(m_axis_scalar_5_tvalid),
        .m_axis_scalar_5_tkeep(m_axis_scalar_5_tkeep),
        .m_axis_scalar_5_tstrb(m_axis_scalar_5_tstrb),
        .m_axis_scalar_5_tdata(m_axis_scalar_5_tdata),
        .m_axis_scalar_5_tready(m_axis_scalar_5_tready),
        .m_axis_scalar_6_aclk(m_axis_scalar_6_aclk),
        .m_axis_scalar_6_aresetn(m_axis_scalar_6_aresetn),
        .m_axis_scalar_6_tlast(m_axis_scalar_6_tlast),
        .m_axis_scalar_6_tvalid(m_axis_scalar_6_tvalid),
        .m_axis_scalar_6_tkeep(m_axis_scalar_6_tkeep),
        .m_axis_scalar_6_tstrb(m_axis_scalar_6_tstrb),
        .m_axis_scalar_6_tdata(m_axis_scalar_6_tdata),
        .m_axis_scalar_6_tready(m_axis_scalar_6_tready),
        .m_axis_scalar_7_aclk(m_axis_scalar_7_aclk),
        .m_axis_scalar_7_aresetn(m_axis_scalar_7_aresetn),
        .m_axis_scalar_7_tlast(m_axis_scalar_7_tlast),
        .m_axis_scalar_7_tvalid(m_axis_scalar_7_tvalid),
        .m_axis_scalar_7_tkeep(m_axis_scalar_7_tkeep),
        .m_axis_scalar_7_tstrb(m_axis_scalar_7_tstrb),
        .m_axis_scalar_7_tdata(m_axis_scalar_7_tdata),
        .m_axis_scalar_7_tready(m_axis_scalar_7_tready),
        .m_axis_scalar_8_aclk(m_axis_scalar_8_aclk),
        .m_axis_scalar_8_aresetn(m_axis_scalar_8_aresetn),
        .m_axis_scalar_8_tlast(m_axis_scalar_8_tlast),
        .m_axis_scalar_8_tvalid(m_axis_scalar_8_tvalid),
        .m_axis_scalar_8_tkeep(m_axis_scalar_8_tkeep),
        .m_axis_scalar_8_tstrb(m_axis_scalar_8_tstrb),
        .m_axis_scalar_8_tdata(m_axis_scalar_8_tdata),
        .m_axis_scalar_8_tready(m_axis_scalar_8_tready),
        .m_axis_scalar_9_aclk(m_axis_scalar_9_aclk),
        .m_axis_scalar_9_aresetn(m_axis_scalar_9_aresetn),
        .m_axis_scalar_9_tlast(m_axis_scalar_9_tlast),
        .m_axis_scalar_9_tvalid(m_axis_scalar_9_tvalid),
        .m_axis_scalar_9_tkeep(m_axis_scalar_9_tkeep),
        .m_axis_scalar_9_tstrb(m_axis_scalar_9_tstrb),
        .m_axis_scalar_9_tdata(m_axis_scalar_9_tdata),
        .m_axis_scalar_9_tready(m_axis_scalar_9_tready),
        .m_axis_scalar_10_aclk(m_axis_scalar_10_aclk),
        .m_axis_scalar_10_aresetn(m_axis_scalar_10_aresetn),
        .m_axis_scalar_10_tlast(m_axis_scalar_10_tlast),
        .m_axis_scalar_10_tvalid(m_axis_scalar_10_tvalid),
        .m_axis_scalar_10_tkeep(m_axis_scalar_10_tkeep),
        .m_axis_scalar_10_tstrb(m_axis_scalar_10_tstrb),
        .m_axis_scalar_10_tdata(m_axis_scalar_10_tdata),
        .m_axis_scalar_10_tready(m_axis_scalar_10_tready),
        .m_axis_scalar_11_aclk(m_axis_scalar_11_aclk),
        .m_axis_scalar_11_aresetn(m_axis_scalar_11_aresetn),
        .m_axis_scalar_11_tlast(m_axis_scalar_11_tlast),
        .m_axis_scalar_11_tvalid(m_axis_scalar_11_tvalid),
        .m_axis_scalar_11_tkeep(m_axis_scalar_11_tkeep),
        .m_axis_scalar_11_tstrb(m_axis_scalar_11_tstrb),
        .m_axis_scalar_11_tdata(m_axis_scalar_11_tdata),
        .m_axis_scalar_11_tready(m_axis_scalar_11_tready),
        .m_axis_scalar_12_aclk(m_axis_scalar_12_aclk),
        .m_axis_scalar_12_aresetn(m_axis_scalar_12_aresetn),
        .m_axis_scalar_12_tlast(m_axis_scalar_12_tlast),
        .m_axis_scalar_12_tvalid(m_axis_scalar_12_tvalid),
        .m_axis_scalar_12_tkeep(m_axis_scalar_12_tkeep),
        .m_axis_scalar_12_tstrb(m_axis_scalar_12_tstrb),
        .m_axis_scalar_12_tdata(m_axis_scalar_12_tdata),
        .m_axis_scalar_12_tready(m_axis_scalar_12_tready),
        .m_axis_scalar_13_aclk(m_axis_scalar_13_aclk),
        .m_axis_scalar_13_aresetn(m_axis_scalar_13_aresetn),
        .m_axis_scalar_13_tlast(m_axis_scalar_13_tlast),
        .m_axis_scalar_13_tvalid(m_axis_scalar_13_tvalid),
        .m_axis_scalar_13_tkeep(m_axis_scalar_13_tkeep),
        .m_axis_scalar_13_tstrb(m_axis_scalar_13_tstrb),
        .m_axis_scalar_13_tdata(m_axis_scalar_13_tdata),
        .m_axis_scalar_13_tready(m_axis_scalar_13_tready),
        .m_axis_scalar_14_aclk(m_axis_scalar_14_aclk),
        .m_axis_scalar_14_aresetn(m_axis_scalar_14_aresetn),
        .m_axis_scalar_14_tlast(m_axis_scalar_14_tlast),
        .m_axis_scalar_14_tvalid(m_axis_scalar_14_tvalid),
        .m_axis_scalar_14_tkeep(m_axis_scalar_14_tkeep),
        .m_axis_scalar_14_tstrb(m_axis_scalar_14_tstrb),
        .m_axis_scalar_14_tdata(m_axis_scalar_14_tdata),
        .m_axis_scalar_14_tready(m_axis_scalar_14_tready),
        .m_axis_scalar_15_aclk(m_axis_scalar_15_aclk),
        .m_axis_scalar_15_aresetn(m_axis_scalar_15_aresetn),
        .m_axis_scalar_15_tlast(m_axis_scalar_15_tlast),
        .m_axis_scalar_15_tvalid(m_axis_scalar_15_tvalid),
        .m_axis_scalar_15_tkeep(m_axis_scalar_15_tkeep),
        .m_axis_scalar_15_tstrb(m_axis_scalar_15_tstrb),
        .m_axis_scalar_15_tdata(m_axis_scalar_15_tdata),
        .m_axis_scalar_15_tready(m_axis_scalar_15_tready),
        .m_axis_scalar_16_aclk(m_axis_scalar_16_aclk),
        .m_axis_scalar_16_aresetn(m_axis_scalar_16_aresetn),
        .m_axis_scalar_16_tlast(m_axis_scalar_16_tlast),
        .m_axis_scalar_16_tvalid(m_axis_scalar_16_tvalid),
        .m_axis_scalar_16_tkeep(m_axis_scalar_16_tkeep),
        .m_axis_scalar_16_tstrb(m_axis_scalar_16_tstrb),
        .m_axis_scalar_16_tdata(m_axis_scalar_16_tdata),
        .m_axis_scalar_16_tready(m_axis_scalar_16_tready),
        .m_axis_scalar_17_aclk(m_axis_scalar_17_aclk),
        .m_axis_scalar_17_aresetn(m_axis_scalar_17_aresetn),
        .m_axis_scalar_17_tlast(m_axis_scalar_17_tlast),
        .m_axis_scalar_17_tvalid(m_axis_scalar_17_tvalid),
        .m_axis_scalar_17_tkeep(m_axis_scalar_17_tkeep),
        .m_axis_scalar_17_tstrb(m_axis_scalar_17_tstrb),
        .m_axis_scalar_17_tdata(m_axis_scalar_17_tdata),
        .m_axis_scalar_17_tready(m_axis_scalar_17_tready),
        .m_axis_scalar_18_aclk(m_axis_scalar_18_aclk),
        .m_axis_scalar_18_aresetn(m_axis_scalar_18_aresetn),
        .m_axis_scalar_18_tlast(m_axis_scalar_18_tlast),
        .m_axis_scalar_18_tvalid(m_axis_scalar_18_tvalid),
        .m_axis_scalar_18_tkeep(m_axis_scalar_18_tkeep),
        .m_axis_scalar_18_tstrb(m_axis_scalar_18_tstrb),
        .m_axis_scalar_18_tdata(m_axis_scalar_18_tdata),
        .m_axis_scalar_18_tready(m_axis_scalar_18_tready),
        .m_axis_scalar_19_aclk(m_axis_scalar_19_aclk),
        .m_axis_scalar_19_aresetn(m_axis_scalar_19_aresetn),
        .m_axis_scalar_19_tlast(m_axis_scalar_19_tlast),
        .m_axis_scalar_19_tvalid(m_axis_scalar_19_tvalid),
        .m_axis_scalar_19_tkeep(m_axis_scalar_19_tkeep),
        .m_axis_scalar_19_tstrb(m_axis_scalar_19_tstrb),
        .m_axis_scalar_19_tdata(m_axis_scalar_19_tdata),
        .m_axis_scalar_19_tready(m_axis_scalar_19_tready),
        .m_axis_scalar_20_aclk(m_axis_scalar_20_aclk),
        .m_axis_scalar_20_aresetn(m_axis_scalar_20_aresetn),
        .m_axis_scalar_20_tlast(m_axis_scalar_20_tlast),
        .m_axis_scalar_20_tvalid(m_axis_scalar_20_tvalid),
        .m_axis_scalar_20_tkeep(m_axis_scalar_20_tkeep),
        .m_axis_scalar_20_tstrb(m_axis_scalar_20_tstrb),
        .m_axis_scalar_20_tdata(m_axis_scalar_20_tdata),
        .m_axis_scalar_20_tready(m_axis_scalar_20_tready),
        .m_axis_scalar_21_aclk(m_axis_scalar_21_aclk),
        .m_axis_scalar_21_aresetn(m_axis_scalar_21_aresetn),
        .m_axis_scalar_21_tlast(m_axis_scalar_21_tlast),
        .m_axis_scalar_21_tvalid(m_axis_scalar_21_tvalid),
        .m_axis_scalar_21_tkeep(m_axis_scalar_21_tkeep),
        .m_axis_scalar_21_tstrb(m_axis_scalar_21_tstrb),
        .m_axis_scalar_21_tdata(m_axis_scalar_21_tdata),
        .m_axis_scalar_21_tready(m_axis_scalar_21_tready),
        .m_axis_scalar_22_aclk(m_axis_scalar_22_aclk),
        .m_axis_scalar_22_aresetn(m_axis_scalar_22_aresetn),
        .m_axis_scalar_22_tlast(m_axis_scalar_22_tlast),
        .m_axis_scalar_22_tvalid(m_axis_scalar_22_tvalid),
        .m_axis_scalar_22_tkeep(m_axis_scalar_22_tkeep),
        .m_axis_scalar_22_tstrb(m_axis_scalar_22_tstrb),
        .m_axis_scalar_22_tdata(m_axis_scalar_22_tdata),
        .m_axis_scalar_22_tready(m_axis_scalar_22_tready),
        .m_axis_scalar_23_aclk(m_axis_scalar_23_aclk),
        .m_axis_scalar_23_aresetn(m_axis_scalar_23_aresetn),
        .m_axis_scalar_23_tlast(m_axis_scalar_23_tlast),
        .m_axis_scalar_23_tvalid(m_axis_scalar_23_tvalid),
        .m_axis_scalar_23_tkeep(m_axis_scalar_23_tkeep),
        .m_axis_scalar_23_tstrb(m_axis_scalar_23_tstrb),
        .m_axis_scalar_23_tdata(m_axis_scalar_23_tdata),
        .m_axis_scalar_23_tready(m_axis_scalar_23_tready),
        .m_axis_scalar_24_aclk(m_axis_scalar_24_aclk),
        .m_axis_scalar_24_aresetn(m_axis_scalar_24_aresetn),
        .m_axis_scalar_24_tlast(m_axis_scalar_24_tlast),
        .m_axis_scalar_24_tvalid(m_axis_scalar_24_tvalid),
        .m_axis_scalar_24_tkeep(m_axis_scalar_24_tkeep),
        .m_axis_scalar_24_tstrb(m_axis_scalar_24_tstrb),
        .m_axis_scalar_24_tdata(m_axis_scalar_24_tdata),
        .m_axis_scalar_24_tready(m_axis_scalar_24_tready),
        .m_axis_scalar_25_aclk(m_axis_scalar_25_aclk),
        .m_axis_scalar_25_aresetn(m_axis_scalar_25_aresetn),
        .m_axis_scalar_25_tlast(m_axis_scalar_25_tlast),
        .m_axis_scalar_25_tvalid(m_axis_scalar_25_tvalid),
        .m_axis_scalar_25_tkeep(m_axis_scalar_25_tkeep),
        .m_axis_scalar_25_tstrb(m_axis_scalar_25_tstrb),
        .m_axis_scalar_25_tdata(m_axis_scalar_25_tdata),
        .m_axis_scalar_25_tready(m_axis_scalar_25_tready),
        .m_axis_scalar_26_aclk(m_axis_scalar_26_aclk),
        .m_axis_scalar_26_aresetn(m_axis_scalar_26_aresetn),
        .m_axis_scalar_26_tlast(m_axis_scalar_26_tlast),
        .m_axis_scalar_26_tvalid(m_axis_scalar_26_tvalid),
        .m_axis_scalar_26_tkeep(m_axis_scalar_26_tkeep),
        .m_axis_scalar_26_tstrb(m_axis_scalar_26_tstrb),
        .m_axis_scalar_26_tdata(m_axis_scalar_26_tdata),
        .m_axis_scalar_26_tready(m_axis_scalar_26_tready),
        .m_axis_scalar_27_aclk(m_axis_scalar_27_aclk),
        .m_axis_scalar_27_aresetn(m_axis_scalar_27_aresetn),
        .m_axis_scalar_27_tlast(m_axis_scalar_27_tlast),
        .m_axis_scalar_27_tvalid(m_axis_scalar_27_tvalid),
        .m_axis_scalar_27_tkeep(m_axis_scalar_27_tkeep),
        .m_axis_scalar_27_tstrb(m_axis_scalar_27_tstrb),
        .m_axis_scalar_27_tdata(m_axis_scalar_27_tdata),
        .m_axis_scalar_27_tready(m_axis_scalar_27_tready),
        .m_axis_scalar_28_aclk(m_axis_scalar_28_aclk),
        .m_axis_scalar_28_aresetn(m_axis_scalar_28_aresetn),
        .m_axis_scalar_28_tlast(m_axis_scalar_28_tlast),
        .m_axis_scalar_28_tvalid(m_axis_scalar_28_tvalid),
        .m_axis_scalar_28_tkeep(m_axis_scalar_28_tkeep),
        .m_axis_scalar_28_tstrb(m_axis_scalar_28_tstrb),
        .m_axis_scalar_28_tdata(m_axis_scalar_28_tdata),
        .m_axis_scalar_28_tready(m_axis_scalar_28_tready),
        .m_axis_scalar_29_aclk(m_axis_scalar_29_aclk),
        .m_axis_scalar_29_aresetn(m_axis_scalar_29_aresetn),
        .m_axis_scalar_29_tlast(m_axis_scalar_29_tlast),
        .m_axis_scalar_29_tvalid(m_axis_scalar_29_tvalid),
        .m_axis_scalar_29_tkeep(m_axis_scalar_29_tkeep),
        .m_axis_scalar_29_tstrb(m_axis_scalar_29_tstrb),
        .m_axis_scalar_29_tdata(m_axis_scalar_29_tdata),
        .m_axis_scalar_29_tready(m_axis_scalar_29_tready),
        .m_axis_scalar_30_aclk(m_axis_scalar_30_aclk),
        .m_axis_scalar_30_aresetn(m_axis_scalar_30_aresetn),
        .m_axis_scalar_30_tlast(m_axis_scalar_30_tlast),
        .m_axis_scalar_30_tvalid(m_axis_scalar_30_tvalid),
        .m_axis_scalar_30_tkeep(m_axis_scalar_30_tkeep),
        .m_axis_scalar_30_tstrb(m_axis_scalar_30_tstrb),
        .m_axis_scalar_30_tdata(m_axis_scalar_30_tdata),
        .m_axis_scalar_30_tready(m_axis_scalar_30_tready),
        .m_axis_scalar_31_aclk(m_axis_scalar_31_aclk),
        .m_axis_scalar_31_aresetn(m_axis_scalar_31_aresetn),
        .m_axis_scalar_31_tlast(m_axis_scalar_31_tlast),
        .m_axis_scalar_31_tvalid(m_axis_scalar_31_tvalid),
        .m_axis_scalar_31_tkeep(m_axis_scalar_31_tkeep),
        .m_axis_scalar_31_tstrb(m_axis_scalar_31_tstrb),
        .m_axis_scalar_31_tdata(m_axis_scalar_31_tdata),
        .m_axis_scalar_31_tready(m_axis_scalar_31_tready),
        .m_axis_scalar_32_aclk(m_axis_scalar_32_aclk),
        .m_axis_scalar_32_aresetn(m_axis_scalar_32_aresetn),
        .m_axis_scalar_32_tlast(m_axis_scalar_32_tlast),
        .m_axis_scalar_32_tvalid(m_axis_scalar_32_tvalid),
        .m_axis_scalar_32_tkeep(m_axis_scalar_32_tkeep),
        .m_axis_scalar_32_tstrb(m_axis_scalar_32_tstrb),
        .m_axis_scalar_32_tdata(m_axis_scalar_32_tdata),
        .m_axis_scalar_32_tready(m_axis_scalar_32_tready),
        .m_axis_scalar_33_aclk(m_axis_scalar_33_aclk),
        .m_axis_scalar_33_aresetn(m_axis_scalar_33_aresetn),
        .m_axis_scalar_33_tlast(m_axis_scalar_33_tlast),
        .m_axis_scalar_33_tvalid(m_axis_scalar_33_tvalid),
        .m_axis_scalar_33_tkeep(m_axis_scalar_33_tkeep),
        .m_axis_scalar_33_tstrb(m_axis_scalar_33_tstrb),
        .m_axis_scalar_33_tdata(m_axis_scalar_33_tdata),
        .m_axis_scalar_33_tready(m_axis_scalar_33_tready),
        .m_axis_scalar_34_aclk(m_axis_scalar_34_aclk),
        .m_axis_scalar_34_aresetn(m_axis_scalar_34_aresetn),
        .m_axis_scalar_34_tlast(m_axis_scalar_34_tlast),
        .m_axis_scalar_34_tvalid(m_axis_scalar_34_tvalid),
        .m_axis_scalar_34_tkeep(m_axis_scalar_34_tkeep),
        .m_axis_scalar_34_tstrb(m_axis_scalar_34_tstrb),
        .m_axis_scalar_34_tdata(m_axis_scalar_34_tdata),
        .m_axis_scalar_34_tready(m_axis_scalar_34_tready),
        .m_axis_scalar_35_aclk(m_axis_scalar_35_aclk),
        .m_axis_scalar_35_aresetn(m_axis_scalar_35_aresetn),
        .m_axis_scalar_35_tlast(m_axis_scalar_35_tlast),
        .m_axis_scalar_35_tvalid(m_axis_scalar_35_tvalid),
        .m_axis_scalar_35_tkeep(m_axis_scalar_35_tkeep),
        .m_axis_scalar_35_tstrb(m_axis_scalar_35_tstrb),
        .m_axis_scalar_35_tdata(m_axis_scalar_35_tdata),
        .m_axis_scalar_35_tready(m_axis_scalar_35_tready),
        .m_axis_scalar_36_aclk(m_axis_scalar_36_aclk),
        .m_axis_scalar_36_aresetn(m_axis_scalar_36_aresetn),
        .m_axis_scalar_36_tlast(m_axis_scalar_36_tlast),
        .m_axis_scalar_36_tvalid(m_axis_scalar_36_tvalid),
        .m_axis_scalar_36_tkeep(m_axis_scalar_36_tkeep),
        .m_axis_scalar_36_tstrb(m_axis_scalar_36_tstrb),
        .m_axis_scalar_36_tdata(m_axis_scalar_36_tdata),
        .m_axis_scalar_36_tready(m_axis_scalar_36_tready),
        .m_axis_scalar_37_aclk(m_axis_scalar_37_aclk),
        .m_axis_scalar_37_aresetn(m_axis_scalar_37_aresetn),
        .m_axis_scalar_37_tlast(m_axis_scalar_37_tlast),
        .m_axis_scalar_37_tvalid(m_axis_scalar_37_tvalid),
        .m_axis_scalar_37_tkeep(m_axis_scalar_37_tkeep),
        .m_axis_scalar_37_tstrb(m_axis_scalar_37_tstrb),
        .m_axis_scalar_37_tdata(m_axis_scalar_37_tdata),
        .m_axis_scalar_37_tready(m_axis_scalar_37_tready),
        .m_axis_scalar_38_aclk(m_axis_scalar_38_aclk),
        .m_axis_scalar_38_aresetn(m_axis_scalar_38_aresetn),
        .m_axis_scalar_38_tlast(m_axis_scalar_38_tlast),
        .m_axis_scalar_38_tvalid(m_axis_scalar_38_tvalid),
        .m_axis_scalar_38_tkeep(m_axis_scalar_38_tkeep),
        .m_axis_scalar_38_tstrb(m_axis_scalar_38_tstrb),
        .m_axis_scalar_38_tdata(m_axis_scalar_38_tdata),
        .m_axis_scalar_38_tready(m_axis_scalar_38_tready),
        .m_axis_scalar_39_aclk(m_axis_scalar_39_aclk),
        .m_axis_scalar_39_aresetn(m_axis_scalar_39_aresetn),
        .m_axis_scalar_39_tlast(m_axis_scalar_39_tlast),
        .m_axis_scalar_39_tvalid(m_axis_scalar_39_tvalid),
        .m_axis_scalar_39_tkeep(m_axis_scalar_39_tkeep),
        .m_axis_scalar_39_tstrb(m_axis_scalar_39_tstrb),
        .m_axis_scalar_39_tdata(m_axis_scalar_39_tdata),
        .m_axis_scalar_39_tready(m_axis_scalar_39_tready),
        .m_axis_scalar_40_aclk(m_axis_scalar_40_aclk),
        .m_axis_scalar_40_aresetn(m_axis_scalar_40_aresetn),
        .m_axis_scalar_40_tlast(m_axis_scalar_40_tlast),
        .m_axis_scalar_40_tvalid(m_axis_scalar_40_tvalid),
        .m_axis_scalar_40_tkeep(m_axis_scalar_40_tkeep),
        .m_axis_scalar_40_tstrb(m_axis_scalar_40_tstrb),
        .m_axis_scalar_40_tdata(m_axis_scalar_40_tdata),
        .m_axis_scalar_40_tready(m_axis_scalar_40_tready),
        .m_axis_scalar_41_aclk(m_axis_scalar_41_aclk),
        .m_axis_scalar_41_aresetn(m_axis_scalar_41_aresetn),
        .m_axis_scalar_41_tlast(m_axis_scalar_41_tlast),
        .m_axis_scalar_41_tvalid(m_axis_scalar_41_tvalid),
        .m_axis_scalar_41_tkeep(m_axis_scalar_41_tkeep),
        .m_axis_scalar_41_tstrb(m_axis_scalar_41_tstrb),
        .m_axis_scalar_41_tdata(m_axis_scalar_41_tdata),
        .m_axis_scalar_41_tready(m_axis_scalar_41_tready),
        .m_axis_scalar_42_aclk(m_axis_scalar_42_aclk),
        .m_axis_scalar_42_aresetn(m_axis_scalar_42_aresetn),
        .m_axis_scalar_42_tlast(m_axis_scalar_42_tlast),
        .m_axis_scalar_42_tvalid(m_axis_scalar_42_tvalid),
        .m_axis_scalar_42_tkeep(m_axis_scalar_42_tkeep),
        .m_axis_scalar_42_tstrb(m_axis_scalar_42_tstrb),
        .m_axis_scalar_42_tdata(m_axis_scalar_42_tdata),
        .m_axis_scalar_42_tready(m_axis_scalar_42_tready),
        .m_axis_scalar_43_aclk(m_axis_scalar_43_aclk),
        .m_axis_scalar_43_aresetn(m_axis_scalar_43_aresetn),
        .m_axis_scalar_43_tlast(m_axis_scalar_43_tlast),
        .m_axis_scalar_43_tvalid(m_axis_scalar_43_tvalid),
        .m_axis_scalar_43_tkeep(m_axis_scalar_43_tkeep),
        .m_axis_scalar_43_tstrb(m_axis_scalar_43_tstrb),
        .m_axis_scalar_43_tdata(m_axis_scalar_43_tdata),
        .m_axis_scalar_43_tready(m_axis_scalar_43_tready),
        .m_axis_scalar_44_aclk(m_axis_scalar_44_aclk),
        .m_axis_scalar_44_aresetn(m_axis_scalar_44_aresetn),
        .m_axis_scalar_44_tlast(m_axis_scalar_44_tlast),
        .m_axis_scalar_44_tvalid(m_axis_scalar_44_tvalid),
        .m_axis_scalar_44_tkeep(m_axis_scalar_44_tkeep),
        .m_axis_scalar_44_tstrb(m_axis_scalar_44_tstrb),
        .m_axis_scalar_44_tdata(m_axis_scalar_44_tdata),
        .m_axis_scalar_44_tready(m_axis_scalar_44_tready),
        .m_axis_scalar_45_aclk(m_axis_scalar_45_aclk),
        .m_axis_scalar_45_aresetn(m_axis_scalar_45_aresetn),
        .m_axis_scalar_45_tlast(m_axis_scalar_45_tlast),
        .m_axis_scalar_45_tvalid(m_axis_scalar_45_tvalid),
        .m_axis_scalar_45_tkeep(m_axis_scalar_45_tkeep),
        .m_axis_scalar_45_tstrb(m_axis_scalar_45_tstrb),
        .m_axis_scalar_45_tdata(m_axis_scalar_45_tdata),
        .m_axis_scalar_45_tready(m_axis_scalar_45_tready),
        .m_axis_scalar_46_aclk(m_axis_scalar_46_aclk),
        .m_axis_scalar_46_aresetn(m_axis_scalar_46_aresetn),
        .m_axis_scalar_46_tlast(m_axis_scalar_46_tlast),
        .m_axis_scalar_46_tvalid(m_axis_scalar_46_tvalid),
        .m_axis_scalar_46_tkeep(m_axis_scalar_46_tkeep),
        .m_axis_scalar_46_tstrb(m_axis_scalar_46_tstrb),
        .m_axis_scalar_46_tdata(m_axis_scalar_46_tdata),
        .m_axis_scalar_46_tready(m_axis_scalar_46_tready),
        .m_axis_scalar_47_aclk(m_axis_scalar_47_aclk),
        .m_axis_scalar_47_aresetn(m_axis_scalar_47_aresetn),
        .m_axis_scalar_47_tlast(m_axis_scalar_47_tlast),
        .m_axis_scalar_47_tvalid(m_axis_scalar_47_tvalid),
        .m_axis_scalar_47_tkeep(m_axis_scalar_47_tkeep),
        .m_axis_scalar_47_tstrb(m_axis_scalar_47_tstrb),
        .m_axis_scalar_47_tdata(m_axis_scalar_47_tdata),
        .m_axis_scalar_47_tready(m_axis_scalar_47_tready),
        .m_axis_scalar_48_aclk(m_axis_scalar_48_aclk),
        .m_axis_scalar_48_aresetn(m_axis_scalar_48_aresetn),
        .m_axis_scalar_48_tlast(m_axis_scalar_48_tlast),
        .m_axis_scalar_48_tvalid(m_axis_scalar_48_tvalid),
        .m_axis_scalar_48_tkeep(m_axis_scalar_48_tkeep),
        .m_axis_scalar_48_tstrb(m_axis_scalar_48_tstrb),
        .m_axis_scalar_48_tdata(m_axis_scalar_48_tdata),
        .m_axis_scalar_48_tready(m_axis_scalar_48_tready),
        .m_axis_scalar_49_aclk(m_axis_scalar_49_aclk),
        .m_axis_scalar_49_aresetn(m_axis_scalar_49_aresetn),
        .m_axis_scalar_49_tlast(m_axis_scalar_49_tlast),
        .m_axis_scalar_49_tvalid(m_axis_scalar_49_tvalid),
        .m_axis_scalar_49_tkeep(m_axis_scalar_49_tkeep),
        .m_axis_scalar_49_tstrb(m_axis_scalar_49_tstrb),
        .m_axis_scalar_49_tdata(m_axis_scalar_49_tdata),
        .m_axis_scalar_49_tready(m_axis_scalar_49_tready),
        .m_axis_scalar_50_aclk(m_axis_scalar_50_aclk),
        .m_axis_scalar_50_aresetn(m_axis_scalar_50_aresetn),
        .m_axis_scalar_50_tlast(m_axis_scalar_50_tlast),
        .m_axis_scalar_50_tvalid(m_axis_scalar_50_tvalid),
        .m_axis_scalar_50_tkeep(m_axis_scalar_50_tkeep),
        .m_axis_scalar_50_tstrb(m_axis_scalar_50_tstrb),
        .m_axis_scalar_50_tdata(m_axis_scalar_50_tdata),
        .m_axis_scalar_50_tready(m_axis_scalar_50_tready),
        .m_axis_scalar_51_aclk(m_axis_scalar_51_aclk),
        .m_axis_scalar_51_aresetn(m_axis_scalar_51_aresetn),
        .m_axis_scalar_51_tlast(m_axis_scalar_51_tlast),
        .m_axis_scalar_51_tvalid(m_axis_scalar_51_tvalid),
        .m_axis_scalar_51_tkeep(m_axis_scalar_51_tkeep),
        .m_axis_scalar_51_tstrb(m_axis_scalar_51_tstrb),
        .m_axis_scalar_51_tdata(m_axis_scalar_51_tdata),
        .m_axis_scalar_51_tready(m_axis_scalar_51_tready),
        .m_axis_scalar_52_aclk(m_axis_scalar_52_aclk),
        .m_axis_scalar_52_aresetn(m_axis_scalar_52_aresetn),
        .m_axis_scalar_52_tlast(m_axis_scalar_52_tlast),
        .m_axis_scalar_52_tvalid(m_axis_scalar_52_tvalid),
        .m_axis_scalar_52_tkeep(m_axis_scalar_52_tkeep),
        .m_axis_scalar_52_tstrb(m_axis_scalar_52_tstrb),
        .m_axis_scalar_52_tdata(m_axis_scalar_52_tdata),
        .m_axis_scalar_52_tready(m_axis_scalar_52_tready),
        .m_axis_scalar_53_aclk(m_axis_scalar_53_aclk),
        .m_axis_scalar_53_aresetn(m_axis_scalar_53_aresetn),
        .m_axis_scalar_53_tlast(m_axis_scalar_53_tlast),
        .m_axis_scalar_53_tvalid(m_axis_scalar_53_tvalid),
        .m_axis_scalar_53_tkeep(m_axis_scalar_53_tkeep),
        .m_axis_scalar_53_tstrb(m_axis_scalar_53_tstrb),
        .m_axis_scalar_53_tdata(m_axis_scalar_53_tdata),
        .m_axis_scalar_53_tready(m_axis_scalar_53_tready),
        .m_axis_scalar_54_aclk(m_axis_scalar_54_aclk),
        .m_axis_scalar_54_aresetn(m_axis_scalar_54_aresetn),
        .m_axis_scalar_54_tlast(m_axis_scalar_54_tlast),
        .m_axis_scalar_54_tvalid(m_axis_scalar_54_tvalid),
        .m_axis_scalar_54_tkeep(m_axis_scalar_54_tkeep),
        .m_axis_scalar_54_tstrb(m_axis_scalar_54_tstrb),
        .m_axis_scalar_54_tdata(m_axis_scalar_54_tdata),
        .m_axis_scalar_54_tready(m_axis_scalar_54_tready),
        .m_axis_scalar_55_aclk(m_axis_scalar_55_aclk),
        .m_axis_scalar_55_aresetn(m_axis_scalar_55_aresetn),
        .m_axis_scalar_55_tlast(m_axis_scalar_55_tlast),
        .m_axis_scalar_55_tvalid(m_axis_scalar_55_tvalid),
        .m_axis_scalar_55_tkeep(m_axis_scalar_55_tkeep),
        .m_axis_scalar_55_tstrb(m_axis_scalar_55_tstrb),
        .m_axis_scalar_55_tdata(m_axis_scalar_55_tdata),
        .m_axis_scalar_55_tready(m_axis_scalar_55_tready),
        .m_axis_scalar_56_aclk(m_axis_scalar_56_aclk),
        .m_axis_scalar_56_aresetn(m_axis_scalar_56_aresetn),
        .m_axis_scalar_56_tlast(m_axis_scalar_56_tlast),
        .m_axis_scalar_56_tvalid(m_axis_scalar_56_tvalid),
        .m_axis_scalar_56_tkeep(m_axis_scalar_56_tkeep),
        .m_axis_scalar_56_tstrb(m_axis_scalar_56_tstrb),
        .m_axis_scalar_56_tdata(m_axis_scalar_56_tdata),
        .m_axis_scalar_56_tready(m_axis_scalar_56_tready),
        .m_axis_scalar_57_aclk(m_axis_scalar_57_aclk),
        .m_axis_scalar_57_aresetn(m_axis_scalar_57_aresetn),
        .m_axis_scalar_57_tlast(m_axis_scalar_57_tlast),
        .m_axis_scalar_57_tvalid(m_axis_scalar_57_tvalid),
        .m_axis_scalar_57_tkeep(m_axis_scalar_57_tkeep),
        .m_axis_scalar_57_tstrb(m_axis_scalar_57_tstrb),
        .m_axis_scalar_57_tdata(m_axis_scalar_57_tdata),
        .m_axis_scalar_57_tready(m_axis_scalar_57_tready),
        .m_axis_scalar_58_aclk(m_axis_scalar_58_aclk),
        .m_axis_scalar_58_aresetn(m_axis_scalar_58_aresetn),
        .m_axis_scalar_58_tlast(m_axis_scalar_58_tlast),
        .m_axis_scalar_58_tvalid(m_axis_scalar_58_tvalid),
        .m_axis_scalar_58_tkeep(m_axis_scalar_58_tkeep),
        .m_axis_scalar_58_tstrb(m_axis_scalar_58_tstrb),
        .m_axis_scalar_58_tdata(m_axis_scalar_58_tdata),
        .m_axis_scalar_58_tready(m_axis_scalar_58_tready),
        .m_axis_scalar_59_aclk(m_axis_scalar_59_aclk),
        .m_axis_scalar_59_aresetn(m_axis_scalar_59_aresetn),
        .m_axis_scalar_59_tlast(m_axis_scalar_59_tlast),
        .m_axis_scalar_59_tvalid(m_axis_scalar_59_tvalid),
        .m_axis_scalar_59_tkeep(m_axis_scalar_59_tkeep),
        .m_axis_scalar_59_tstrb(m_axis_scalar_59_tstrb),
        .m_axis_scalar_59_tdata(m_axis_scalar_59_tdata),
        .m_axis_scalar_59_tready(m_axis_scalar_59_tready),
        .m_axis_scalar_60_aclk(m_axis_scalar_60_aclk),
        .m_axis_scalar_60_aresetn(m_axis_scalar_60_aresetn),
        .m_axis_scalar_60_tlast(m_axis_scalar_60_tlast),
        .m_axis_scalar_60_tvalid(m_axis_scalar_60_tvalid),
        .m_axis_scalar_60_tkeep(m_axis_scalar_60_tkeep),
        .m_axis_scalar_60_tstrb(m_axis_scalar_60_tstrb),
        .m_axis_scalar_60_tdata(m_axis_scalar_60_tdata),
        .m_axis_scalar_60_tready(m_axis_scalar_60_tready),
        .m_axis_scalar_61_aclk(m_axis_scalar_61_aclk),
        .m_axis_scalar_61_aresetn(m_axis_scalar_61_aresetn),
        .m_axis_scalar_61_tlast(m_axis_scalar_61_tlast),
        .m_axis_scalar_61_tvalid(m_axis_scalar_61_tvalid),
        .m_axis_scalar_61_tkeep(m_axis_scalar_61_tkeep),
        .m_axis_scalar_61_tstrb(m_axis_scalar_61_tstrb),
        .m_axis_scalar_61_tdata(m_axis_scalar_61_tdata),
        .m_axis_scalar_61_tready(m_axis_scalar_61_tready),
        .m_axis_scalar_62_aclk(m_axis_scalar_62_aclk),
        .m_axis_scalar_62_aresetn(m_axis_scalar_62_aresetn),
        .m_axis_scalar_62_tlast(m_axis_scalar_62_tlast),
        .m_axis_scalar_62_tvalid(m_axis_scalar_62_tvalid),
        .m_axis_scalar_62_tkeep(m_axis_scalar_62_tkeep),
        .m_axis_scalar_62_tstrb(m_axis_scalar_62_tstrb),
        .m_axis_scalar_62_tdata(m_axis_scalar_62_tdata),
        .m_axis_scalar_62_tready(m_axis_scalar_62_tready),
        .m_axis_scalar_63_aclk(m_axis_scalar_63_aclk),
        .m_axis_scalar_63_aresetn(m_axis_scalar_63_aresetn),
        .m_axis_scalar_63_tlast(m_axis_scalar_63_tlast),
        .m_axis_scalar_63_tvalid(m_axis_scalar_63_tvalid),
        .m_axis_scalar_63_tkeep(m_axis_scalar_63_tkeep),
        .m_axis_scalar_63_tstrb(m_axis_scalar_63_tstrb),
        .m_axis_scalar_63_tdata(m_axis_scalar_63_tdata),
        .m_axis_scalar_63_tready(m_axis_scalar_63_tready),
        .m_axis_scalar_64_aclk(m_axis_scalar_64_aclk),
        .m_axis_scalar_64_aresetn(m_axis_scalar_64_aresetn),
        .m_axis_scalar_64_tlast(m_axis_scalar_64_tlast),
        .m_axis_scalar_64_tvalid(m_axis_scalar_64_tvalid),
        .m_axis_scalar_64_tkeep(m_axis_scalar_64_tkeep),
        .m_axis_scalar_64_tstrb(m_axis_scalar_64_tstrb),
        .m_axis_scalar_64_tdata(m_axis_scalar_64_tdata),
        .m_axis_scalar_64_tready(m_axis_scalar_64_tready),
        .m_axis_scalar_65_aclk(m_axis_scalar_65_aclk),
        .m_axis_scalar_65_aresetn(m_axis_scalar_65_aresetn),
        .m_axis_scalar_65_tlast(m_axis_scalar_65_tlast),
        .m_axis_scalar_65_tvalid(m_axis_scalar_65_tvalid),
        .m_axis_scalar_65_tkeep(m_axis_scalar_65_tkeep),
        .m_axis_scalar_65_tstrb(m_axis_scalar_65_tstrb),
        .m_axis_scalar_65_tdata(m_axis_scalar_65_tdata),
        .m_axis_scalar_65_tready(m_axis_scalar_65_tready),
        .m_axis_scalar_66_aclk(m_axis_scalar_66_aclk),
        .m_axis_scalar_66_aresetn(m_axis_scalar_66_aresetn),
        .m_axis_scalar_66_tlast(m_axis_scalar_66_tlast),
        .m_axis_scalar_66_tvalid(m_axis_scalar_66_tvalid),
        .m_axis_scalar_66_tkeep(m_axis_scalar_66_tkeep),
        .m_axis_scalar_66_tstrb(m_axis_scalar_66_tstrb),
        .m_axis_scalar_66_tdata(m_axis_scalar_66_tdata),
        .m_axis_scalar_66_tready(m_axis_scalar_66_tready),
        .m_axis_scalar_67_aclk(m_axis_scalar_67_aclk),
        .m_axis_scalar_67_aresetn(m_axis_scalar_67_aresetn),
        .m_axis_scalar_67_tlast(m_axis_scalar_67_tlast),
        .m_axis_scalar_67_tvalid(m_axis_scalar_67_tvalid),
        .m_axis_scalar_67_tkeep(m_axis_scalar_67_tkeep),
        .m_axis_scalar_67_tstrb(m_axis_scalar_67_tstrb),
        .m_axis_scalar_67_tdata(m_axis_scalar_67_tdata),
        .m_axis_scalar_67_tready(m_axis_scalar_67_tready),
        .m_axis_scalar_68_aclk(m_axis_scalar_68_aclk),
        .m_axis_scalar_68_aresetn(m_axis_scalar_68_aresetn),
        .m_axis_scalar_68_tlast(m_axis_scalar_68_tlast),
        .m_axis_scalar_68_tvalid(m_axis_scalar_68_tvalid),
        .m_axis_scalar_68_tkeep(m_axis_scalar_68_tkeep),
        .m_axis_scalar_68_tstrb(m_axis_scalar_68_tstrb),
        .m_axis_scalar_68_tdata(m_axis_scalar_68_tdata),
        .m_axis_scalar_68_tready(m_axis_scalar_68_tready),
        .m_axis_scalar_69_aclk(m_axis_scalar_69_aclk),
        .m_axis_scalar_69_aresetn(m_axis_scalar_69_aresetn),
        .m_axis_scalar_69_tlast(m_axis_scalar_69_tlast),
        .m_axis_scalar_69_tvalid(m_axis_scalar_69_tvalid),
        .m_axis_scalar_69_tkeep(m_axis_scalar_69_tkeep),
        .m_axis_scalar_69_tstrb(m_axis_scalar_69_tstrb),
        .m_axis_scalar_69_tdata(m_axis_scalar_69_tdata),
        .m_axis_scalar_69_tready(m_axis_scalar_69_tready),
        .m_axis_scalar_70_aclk(m_axis_scalar_70_aclk),
        .m_axis_scalar_70_aresetn(m_axis_scalar_70_aresetn),
        .m_axis_scalar_70_tlast(m_axis_scalar_70_tlast),
        .m_axis_scalar_70_tvalid(m_axis_scalar_70_tvalid),
        .m_axis_scalar_70_tkeep(m_axis_scalar_70_tkeep),
        .m_axis_scalar_70_tstrb(m_axis_scalar_70_tstrb),
        .m_axis_scalar_70_tdata(m_axis_scalar_70_tdata),
        .m_axis_scalar_70_tready(m_axis_scalar_70_tready),
        .m_axis_scalar_71_aclk(m_axis_scalar_71_aclk),
        .m_axis_scalar_71_aresetn(m_axis_scalar_71_aresetn),
        .m_axis_scalar_71_tlast(m_axis_scalar_71_tlast),
        .m_axis_scalar_71_tvalid(m_axis_scalar_71_tvalid),
        .m_axis_scalar_71_tkeep(m_axis_scalar_71_tkeep),
        .m_axis_scalar_71_tstrb(m_axis_scalar_71_tstrb),
        .m_axis_scalar_71_tdata(m_axis_scalar_71_tdata),
        .m_axis_scalar_71_tready(m_axis_scalar_71_tready),
        .m_axis_scalar_72_aclk(m_axis_scalar_72_aclk),
        .m_axis_scalar_72_aresetn(m_axis_scalar_72_aresetn),
        .m_axis_scalar_72_tlast(m_axis_scalar_72_tlast),
        .m_axis_scalar_72_tvalid(m_axis_scalar_72_tvalid),
        .m_axis_scalar_72_tkeep(m_axis_scalar_72_tkeep),
        .m_axis_scalar_72_tstrb(m_axis_scalar_72_tstrb),
        .m_axis_scalar_72_tdata(m_axis_scalar_72_tdata),
        .m_axis_scalar_72_tready(m_axis_scalar_72_tready),
        .m_axis_scalar_73_aclk(m_axis_scalar_73_aclk),
        .m_axis_scalar_73_aresetn(m_axis_scalar_73_aresetn),
        .m_axis_scalar_73_tlast(m_axis_scalar_73_tlast),
        .m_axis_scalar_73_tvalid(m_axis_scalar_73_tvalid),
        .m_axis_scalar_73_tkeep(m_axis_scalar_73_tkeep),
        .m_axis_scalar_73_tstrb(m_axis_scalar_73_tstrb),
        .m_axis_scalar_73_tdata(m_axis_scalar_73_tdata),
        .m_axis_scalar_73_tready(m_axis_scalar_73_tready),
        .m_axis_scalar_74_aclk(m_axis_scalar_74_aclk),
        .m_axis_scalar_74_aresetn(m_axis_scalar_74_aresetn),
        .m_axis_scalar_74_tlast(m_axis_scalar_74_tlast),
        .m_axis_scalar_74_tvalid(m_axis_scalar_74_tvalid),
        .m_axis_scalar_74_tkeep(m_axis_scalar_74_tkeep),
        .m_axis_scalar_74_tstrb(m_axis_scalar_74_tstrb),
        .m_axis_scalar_74_tdata(m_axis_scalar_74_tdata),
        .m_axis_scalar_74_tready(m_axis_scalar_74_tready),
        .m_axis_scalar_75_aclk(m_axis_scalar_75_aclk),
        .m_axis_scalar_75_aresetn(m_axis_scalar_75_aresetn),
        .m_axis_scalar_75_tlast(m_axis_scalar_75_tlast),
        .m_axis_scalar_75_tvalid(m_axis_scalar_75_tvalid),
        .m_axis_scalar_75_tkeep(m_axis_scalar_75_tkeep),
        .m_axis_scalar_75_tstrb(m_axis_scalar_75_tstrb),
        .m_axis_scalar_75_tdata(m_axis_scalar_75_tdata),
        .m_axis_scalar_75_tready(m_axis_scalar_75_tready),
        .m_axis_scalar_76_aclk(m_axis_scalar_76_aclk),
        .m_axis_scalar_76_aresetn(m_axis_scalar_76_aresetn),
        .m_axis_scalar_76_tlast(m_axis_scalar_76_tlast),
        .m_axis_scalar_76_tvalid(m_axis_scalar_76_tvalid),
        .m_axis_scalar_76_tkeep(m_axis_scalar_76_tkeep),
        .m_axis_scalar_76_tstrb(m_axis_scalar_76_tstrb),
        .m_axis_scalar_76_tdata(m_axis_scalar_76_tdata),
        .m_axis_scalar_76_tready(m_axis_scalar_76_tready),
        .m_axis_scalar_77_aclk(m_axis_scalar_77_aclk),
        .m_axis_scalar_77_aresetn(m_axis_scalar_77_aresetn),
        .m_axis_scalar_77_tlast(m_axis_scalar_77_tlast),
        .m_axis_scalar_77_tvalid(m_axis_scalar_77_tvalid),
        .m_axis_scalar_77_tkeep(m_axis_scalar_77_tkeep),
        .m_axis_scalar_77_tstrb(m_axis_scalar_77_tstrb),
        .m_axis_scalar_77_tdata(m_axis_scalar_77_tdata),
        .m_axis_scalar_77_tready(m_axis_scalar_77_tready),
        .m_axis_scalar_78_aclk(m_axis_scalar_78_aclk),
        .m_axis_scalar_78_aresetn(m_axis_scalar_78_aresetn),
        .m_axis_scalar_78_tlast(m_axis_scalar_78_tlast),
        .m_axis_scalar_78_tvalid(m_axis_scalar_78_tvalid),
        .m_axis_scalar_78_tkeep(m_axis_scalar_78_tkeep),
        .m_axis_scalar_78_tstrb(m_axis_scalar_78_tstrb),
        .m_axis_scalar_78_tdata(m_axis_scalar_78_tdata),
        .m_axis_scalar_78_tready(m_axis_scalar_78_tready),
        .m_axis_scalar_79_aclk(m_axis_scalar_79_aclk),
        .m_axis_scalar_79_aresetn(m_axis_scalar_79_aresetn),
        .m_axis_scalar_79_tlast(m_axis_scalar_79_tlast),
        .m_axis_scalar_79_tvalid(m_axis_scalar_79_tvalid),
        .m_axis_scalar_79_tkeep(m_axis_scalar_79_tkeep),
        .m_axis_scalar_79_tstrb(m_axis_scalar_79_tstrb),
        .m_axis_scalar_79_tdata(m_axis_scalar_79_tdata),
        .m_axis_scalar_79_tready(m_axis_scalar_79_tready),
        .m_axis_scalar_80_aclk(m_axis_scalar_80_aclk),
        .m_axis_scalar_80_aresetn(m_axis_scalar_80_aresetn),
        .m_axis_scalar_80_tlast(m_axis_scalar_80_tlast),
        .m_axis_scalar_80_tvalid(m_axis_scalar_80_tvalid),
        .m_axis_scalar_80_tkeep(m_axis_scalar_80_tkeep),
        .m_axis_scalar_80_tstrb(m_axis_scalar_80_tstrb),
        .m_axis_scalar_80_tdata(m_axis_scalar_80_tdata),
        .m_axis_scalar_80_tready(m_axis_scalar_80_tready),
        .m_axis_scalar_81_aclk(m_axis_scalar_81_aclk),
        .m_axis_scalar_81_aresetn(m_axis_scalar_81_aresetn),
        .m_axis_scalar_81_tlast(m_axis_scalar_81_tlast),
        .m_axis_scalar_81_tvalid(m_axis_scalar_81_tvalid),
        .m_axis_scalar_81_tkeep(m_axis_scalar_81_tkeep),
        .m_axis_scalar_81_tstrb(m_axis_scalar_81_tstrb),
        .m_axis_scalar_81_tdata(m_axis_scalar_81_tdata),
        .m_axis_scalar_81_tready(m_axis_scalar_81_tready),
        .m_axis_scalar_82_aclk(m_axis_scalar_82_aclk),
        .m_axis_scalar_82_aresetn(m_axis_scalar_82_aresetn),
        .m_axis_scalar_82_tlast(m_axis_scalar_82_tlast),
        .m_axis_scalar_82_tvalid(m_axis_scalar_82_tvalid),
        .m_axis_scalar_82_tkeep(m_axis_scalar_82_tkeep),
        .m_axis_scalar_82_tstrb(m_axis_scalar_82_tstrb),
        .m_axis_scalar_82_tdata(m_axis_scalar_82_tdata),
        .m_axis_scalar_82_tready(m_axis_scalar_82_tready),
        .m_axis_scalar_83_aclk(m_axis_scalar_83_aclk),
        .m_axis_scalar_83_aresetn(m_axis_scalar_83_aresetn),
        .m_axis_scalar_83_tlast(m_axis_scalar_83_tlast),
        .m_axis_scalar_83_tvalid(m_axis_scalar_83_tvalid),
        .m_axis_scalar_83_tkeep(m_axis_scalar_83_tkeep),
        .m_axis_scalar_83_tstrb(m_axis_scalar_83_tstrb),
        .m_axis_scalar_83_tdata(m_axis_scalar_83_tdata),
        .m_axis_scalar_83_tready(m_axis_scalar_83_tready),
        .m_axis_scalar_84_aclk(m_axis_scalar_84_aclk),
        .m_axis_scalar_84_aresetn(m_axis_scalar_84_aresetn),
        .m_axis_scalar_84_tlast(m_axis_scalar_84_tlast),
        .m_axis_scalar_84_tvalid(m_axis_scalar_84_tvalid),
        .m_axis_scalar_84_tkeep(m_axis_scalar_84_tkeep),
        .m_axis_scalar_84_tstrb(m_axis_scalar_84_tstrb),
        .m_axis_scalar_84_tdata(m_axis_scalar_84_tdata),
        .m_axis_scalar_84_tready(m_axis_scalar_84_tready),
        .m_axis_scalar_85_aclk(m_axis_scalar_85_aclk),
        .m_axis_scalar_85_aresetn(m_axis_scalar_85_aresetn),
        .m_axis_scalar_85_tlast(m_axis_scalar_85_tlast),
        .m_axis_scalar_85_tvalid(m_axis_scalar_85_tvalid),
        .m_axis_scalar_85_tkeep(m_axis_scalar_85_tkeep),
        .m_axis_scalar_85_tstrb(m_axis_scalar_85_tstrb),
        .m_axis_scalar_85_tdata(m_axis_scalar_85_tdata),
        .m_axis_scalar_85_tready(m_axis_scalar_85_tready),
        .m_axis_scalar_86_aclk(m_axis_scalar_86_aclk),
        .m_axis_scalar_86_aresetn(m_axis_scalar_86_aresetn),
        .m_axis_scalar_86_tlast(m_axis_scalar_86_tlast),
        .m_axis_scalar_86_tvalid(m_axis_scalar_86_tvalid),
        .m_axis_scalar_86_tkeep(m_axis_scalar_86_tkeep),
        .m_axis_scalar_86_tstrb(m_axis_scalar_86_tstrb),
        .m_axis_scalar_86_tdata(m_axis_scalar_86_tdata),
        .m_axis_scalar_86_tready(m_axis_scalar_86_tready),
        .m_axis_scalar_87_aclk(m_axis_scalar_87_aclk),
        .m_axis_scalar_87_aresetn(m_axis_scalar_87_aresetn),
        .m_axis_scalar_87_tlast(m_axis_scalar_87_tlast),
        .m_axis_scalar_87_tvalid(m_axis_scalar_87_tvalid),
        .m_axis_scalar_87_tkeep(m_axis_scalar_87_tkeep),
        .m_axis_scalar_87_tstrb(m_axis_scalar_87_tstrb),
        .m_axis_scalar_87_tdata(m_axis_scalar_87_tdata),
        .m_axis_scalar_87_tready(m_axis_scalar_87_tready),
        .m_axis_scalar_88_aclk(m_axis_scalar_88_aclk),
        .m_axis_scalar_88_aresetn(m_axis_scalar_88_aresetn),
        .m_axis_scalar_88_tlast(m_axis_scalar_88_tlast),
        .m_axis_scalar_88_tvalid(m_axis_scalar_88_tvalid),
        .m_axis_scalar_88_tkeep(m_axis_scalar_88_tkeep),
        .m_axis_scalar_88_tstrb(m_axis_scalar_88_tstrb),
        .m_axis_scalar_88_tdata(m_axis_scalar_88_tdata),
        .m_axis_scalar_88_tready(m_axis_scalar_88_tready),
        .m_axis_scalar_89_aclk(m_axis_scalar_89_aclk),
        .m_axis_scalar_89_aresetn(m_axis_scalar_89_aresetn),
        .m_axis_scalar_89_tlast(m_axis_scalar_89_tlast),
        .m_axis_scalar_89_tvalid(m_axis_scalar_89_tvalid),
        .m_axis_scalar_89_tkeep(m_axis_scalar_89_tkeep),
        .m_axis_scalar_89_tstrb(m_axis_scalar_89_tstrb),
        .m_axis_scalar_89_tdata(m_axis_scalar_89_tdata),
        .m_axis_scalar_89_tready(m_axis_scalar_89_tready),
        .m_axis_scalar_90_aclk(m_axis_scalar_90_aclk),
        .m_axis_scalar_90_aresetn(m_axis_scalar_90_aresetn),
        .m_axis_scalar_90_tlast(m_axis_scalar_90_tlast),
        .m_axis_scalar_90_tvalid(m_axis_scalar_90_tvalid),
        .m_axis_scalar_90_tkeep(m_axis_scalar_90_tkeep),
        .m_axis_scalar_90_tstrb(m_axis_scalar_90_tstrb),
        .m_axis_scalar_90_tdata(m_axis_scalar_90_tdata),
        .m_axis_scalar_90_tready(m_axis_scalar_90_tready),
        .m_axis_scalar_91_aclk(m_axis_scalar_91_aclk),
        .m_axis_scalar_91_aresetn(m_axis_scalar_91_aresetn),
        .m_axis_scalar_91_tlast(m_axis_scalar_91_tlast),
        .m_axis_scalar_91_tvalid(m_axis_scalar_91_tvalid),
        .m_axis_scalar_91_tkeep(m_axis_scalar_91_tkeep),
        .m_axis_scalar_91_tstrb(m_axis_scalar_91_tstrb),
        .m_axis_scalar_91_tdata(m_axis_scalar_91_tdata),
        .m_axis_scalar_91_tready(m_axis_scalar_91_tready),
        .m_axis_scalar_92_aclk(m_axis_scalar_92_aclk),
        .m_axis_scalar_92_aresetn(m_axis_scalar_92_aresetn),
        .m_axis_scalar_92_tlast(m_axis_scalar_92_tlast),
        .m_axis_scalar_92_tvalid(m_axis_scalar_92_tvalid),
        .m_axis_scalar_92_tkeep(m_axis_scalar_92_tkeep),
        .m_axis_scalar_92_tstrb(m_axis_scalar_92_tstrb),
        .m_axis_scalar_92_tdata(m_axis_scalar_92_tdata),
        .m_axis_scalar_92_tready(m_axis_scalar_92_tready),
        .m_axis_scalar_93_aclk(m_axis_scalar_93_aclk),
        .m_axis_scalar_93_aresetn(m_axis_scalar_93_aresetn),
        .m_axis_scalar_93_tlast(m_axis_scalar_93_tlast),
        .m_axis_scalar_93_tvalid(m_axis_scalar_93_tvalid),
        .m_axis_scalar_93_tkeep(m_axis_scalar_93_tkeep),
        .m_axis_scalar_93_tstrb(m_axis_scalar_93_tstrb),
        .m_axis_scalar_93_tdata(m_axis_scalar_93_tdata),
        .m_axis_scalar_93_tready(m_axis_scalar_93_tready),
        .m_axis_scalar_94_aclk(m_axis_scalar_94_aclk),
        .m_axis_scalar_94_aresetn(m_axis_scalar_94_aresetn),
        .m_axis_scalar_94_tlast(m_axis_scalar_94_tlast),
        .m_axis_scalar_94_tvalid(m_axis_scalar_94_tvalid),
        .m_axis_scalar_94_tkeep(m_axis_scalar_94_tkeep),
        .m_axis_scalar_94_tstrb(m_axis_scalar_94_tstrb),
        .m_axis_scalar_94_tdata(m_axis_scalar_94_tdata),
        .m_axis_scalar_94_tready(m_axis_scalar_94_tready),
        .m_axis_scalar_95_aclk(m_axis_scalar_95_aclk),
        .m_axis_scalar_95_aresetn(m_axis_scalar_95_aresetn),
        .m_axis_scalar_95_tlast(m_axis_scalar_95_tlast),
        .m_axis_scalar_95_tvalid(m_axis_scalar_95_tvalid),
        .m_axis_scalar_95_tkeep(m_axis_scalar_95_tkeep),
        .m_axis_scalar_95_tstrb(m_axis_scalar_95_tstrb),
        .m_axis_scalar_95_tdata(m_axis_scalar_95_tdata),
        .m_axis_scalar_95_tready(m_axis_scalar_95_tready),
        .m_axis_scalar_96_aclk(m_axis_scalar_96_aclk),
        .m_axis_scalar_96_aresetn(m_axis_scalar_96_aresetn),
        .m_axis_scalar_96_tlast(m_axis_scalar_96_tlast),
        .m_axis_scalar_96_tvalid(m_axis_scalar_96_tvalid),
        .m_axis_scalar_96_tkeep(m_axis_scalar_96_tkeep),
        .m_axis_scalar_96_tstrb(m_axis_scalar_96_tstrb),
        .m_axis_scalar_96_tdata(m_axis_scalar_96_tdata),
        .m_axis_scalar_96_tready(m_axis_scalar_96_tready),
        .m_axis_scalar_97_aclk(m_axis_scalar_97_aclk),
        .m_axis_scalar_97_aresetn(m_axis_scalar_97_aresetn),
        .m_axis_scalar_97_tlast(m_axis_scalar_97_tlast),
        .m_axis_scalar_97_tvalid(m_axis_scalar_97_tvalid),
        .m_axis_scalar_97_tkeep(m_axis_scalar_97_tkeep),
        .m_axis_scalar_97_tstrb(m_axis_scalar_97_tstrb),
        .m_axis_scalar_97_tdata(m_axis_scalar_97_tdata),
        .m_axis_scalar_97_tready(m_axis_scalar_97_tready),
        .m_axis_scalar_98_aclk(m_axis_scalar_98_aclk),
        .m_axis_scalar_98_aresetn(m_axis_scalar_98_aresetn),
        .m_axis_scalar_98_tlast(m_axis_scalar_98_tlast),
        .m_axis_scalar_98_tvalid(m_axis_scalar_98_tvalid),
        .m_axis_scalar_98_tkeep(m_axis_scalar_98_tkeep),
        .m_axis_scalar_98_tstrb(m_axis_scalar_98_tstrb),
        .m_axis_scalar_98_tdata(m_axis_scalar_98_tdata),
        .m_axis_scalar_98_tready(m_axis_scalar_98_tready),
        .m_axis_scalar_99_aclk(m_axis_scalar_99_aclk),
        .m_axis_scalar_99_aresetn(m_axis_scalar_99_aresetn),
        .m_axis_scalar_99_tlast(m_axis_scalar_99_tlast),
        .m_axis_scalar_99_tvalid(m_axis_scalar_99_tvalid),
        .m_axis_scalar_99_tkeep(m_axis_scalar_99_tkeep),
        .m_axis_scalar_99_tstrb(m_axis_scalar_99_tstrb),
        .m_axis_scalar_99_tdata(m_axis_scalar_99_tdata),
        .m_axis_scalar_99_tready(m_axis_scalar_99_tready),
        .m_axis_scalar_100_aclk(m_axis_scalar_100_aclk),
        .m_axis_scalar_100_aresetn(m_axis_scalar_100_aresetn),
        .m_axis_scalar_100_tlast(m_axis_scalar_100_tlast),
        .m_axis_scalar_100_tvalid(m_axis_scalar_100_tvalid),
        .m_axis_scalar_100_tkeep(m_axis_scalar_100_tkeep),
        .m_axis_scalar_100_tstrb(m_axis_scalar_100_tstrb),
        .m_axis_scalar_100_tdata(m_axis_scalar_100_tdata),
        .m_axis_scalar_100_tready(m_axis_scalar_100_tready),
        .m_axis_scalar_101_aclk(m_axis_scalar_101_aclk),
        .m_axis_scalar_101_aresetn(m_axis_scalar_101_aresetn),
        .m_axis_scalar_101_tlast(m_axis_scalar_101_tlast),
        .m_axis_scalar_101_tvalid(m_axis_scalar_101_tvalid),
        .m_axis_scalar_101_tkeep(m_axis_scalar_101_tkeep),
        .m_axis_scalar_101_tstrb(m_axis_scalar_101_tstrb),
        .m_axis_scalar_101_tdata(m_axis_scalar_101_tdata),
        .m_axis_scalar_101_tready(m_axis_scalar_101_tready),
        .m_axis_scalar_102_aclk(m_axis_scalar_102_aclk),
        .m_axis_scalar_102_aresetn(m_axis_scalar_102_aresetn),
        .m_axis_scalar_102_tlast(m_axis_scalar_102_tlast),
        .m_axis_scalar_102_tvalid(m_axis_scalar_102_tvalid),
        .m_axis_scalar_102_tkeep(m_axis_scalar_102_tkeep),
        .m_axis_scalar_102_tstrb(m_axis_scalar_102_tstrb),
        .m_axis_scalar_102_tdata(m_axis_scalar_102_tdata),
        .m_axis_scalar_102_tready(m_axis_scalar_102_tready),
        .m_axis_scalar_103_aclk(m_axis_scalar_103_aclk),
        .m_axis_scalar_103_aresetn(m_axis_scalar_103_aresetn),
        .m_axis_scalar_103_tlast(m_axis_scalar_103_tlast),
        .m_axis_scalar_103_tvalid(m_axis_scalar_103_tvalid),
        .m_axis_scalar_103_tkeep(m_axis_scalar_103_tkeep),
        .m_axis_scalar_103_tstrb(m_axis_scalar_103_tstrb),
        .m_axis_scalar_103_tdata(m_axis_scalar_103_tdata),
        .m_axis_scalar_103_tready(m_axis_scalar_103_tready),
        .m_axis_scalar_104_aclk(m_axis_scalar_104_aclk),
        .m_axis_scalar_104_aresetn(m_axis_scalar_104_aresetn),
        .m_axis_scalar_104_tlast(m_axis_scalar_104_tlast),
        .m_axis_scalar_104_tvalid(m_axis_scalar_104_tvalid),
        .m_axis_scalar_104_tkeep(m_axis_scalar_104_tkeep),
        .m_axis_scalar_104_tstrb(m_axis_scalar_104_tstrb),
        .m_axis_scalar_104_tdata(m_axis_scalar_104_tdata),
        .m_axis_scalar_104_tready(m_axis_scalar_104_tready),
        .m_axis_scalar_105_aclk(m_axis_scalar_105_aclk),
        .m_axis_scalar_105_aresetn(m_axis_scalar_105_aresetn),
        .m_axis_scalar_105_tlast(m_axis_scalar_105_tlast),
        .m_axis_scalar_105_tvalid(m_axis_scalar_105_tvalid),
        .m_axis_scalar_105_tkeep(m_axis_scalar_105_tkeep),
        .m_axis_scalar_105_tstrb(m_axis_scalar_105_tstrb),
        .m_axis_scalar_105_tdata(m_axis_scalar_105_tdata),
        .m_axis_scalar_105_tready(m_axis_scalar_105_tready),
        .m_axis_scalar_106_aclk(m_axis_scalar_106_aclk),
        .m_axis_scalar_106_aresetn(m_axis_scalar_106_aresetn),
        .m_axis_scalar_106_tlast(m_axis_scalar_106_tlast),
        .m_axis_scalar_106_tvalid(m_axis_scalar_106_tvalid),
        .m_axis_scalar_106_tkeep(m_axis_scalar_106_tkeep),
        .m_axis_scalar_106_tstrb(m_axis_scalar_106_tstrb),
        .m_axis_scalar_106_tdata(m_axis_scalar_106_tdata),
        .m_axis_scalar_106_tready(m_axis_scalar_106_tready),
        .m_axis_scalar_107_aclk(m_axis_scalar_107_aclk),
        .m_axis_scalar_107_aresetn(m_axis_scalar_107_aresetn),
        .m_axis_scalar_107_tlast(m_axis_scalar_107_tlast),
        .m_axis_scalar_107_tvalid(m_axis_scalar_107_tvalid),
        .m_axis_scalar_107_tkeep(m_axis_scalar_107_tkeep),
        .m_axis_scalar_107_tstrb(m_axis_scalar_107_tstrb),
        .m_axis_scalar_107_tdata(m_axis_scalar_107_tdata),
        .m_axis_scalar_107_tready(m_axis_scalar_107_tready),
        .m_axis_scalar_108_aclk(m_axis_scalar_108_aclk),
        .m_axis_scalar_108_aresetn(m_axis_scalar_108_aresetn),
        .m_axis_scalar_108_tlast(m_axis_scalar_108_tlast),
        .m_axis_scalar_108_tvalid(m_axis_scalar_108_tvalid),
        .m_axis_scalar_108_tkeep(m_axis_scalar_108_tkeep),
        .m_axis_scalar_108_tstrb(m_axis_scalar_108_tstrb),
        .m_axis_scalar_108_tdata(m_axis_scalar_108_tdata),
        .m_axis_scalar_108_tready(m_axis_scalar_108_tready),
        .m_axis_scalar_109_aclk(m_axis_scalar_109_aclk),
        .m_axis_scalar_109_aresetn(m_axis_scalar_109_aresetn),
        .m_axis_scalar_109_tlast(m_axis_scalar_109_tlast),
        .m_axis_scalar_109_tvalid(m_axis_scalar_109_tvalid),
        .m_axis_scalar_109_tkeep(m_axis_scalar_109_tkeep),
        .m_axis_scalar_109_tstrb(m_axis_scalar_109_tstrb),
        .m_axis_scalar_109_tdata(m_axis_scalar_109_tdata),
        .m_axis_scalar_109_tready(m_axis_scalar_109_tready),
        .m_axis_scalar_110_aclk(m_axis_scalar_110_aclk),
        .m_axis_scalar_110_aresetn(m_axis_scalar_110_aresetn),
        .m_axis_scalar_110_tlast(m_axis_scalar_110_tlast),
        .m_axis_scalar_110_tvalid(m_axis_scalar_110_tvalid),
        .m_axis_scalar_110_tkeep(m_axis_scalar_110_tkeep),
        .m_axis_scalar_110_tstrb(m_axis_scalar_110_tstrb),
        .m_axis_scalar_110_tdata(m_axis_scalar_110_tdata),
        .m_axis_scalar_110_tready(m_axis_scalar_110_tready),
        .m_axis_scalar_111_aclk(m_axis_scalar_111_aclk),
        .m_axis_scalar_111_aresetn(m_axis_scalar_111_aresetn),
        .m_axis_scalar_111_tlast(m_axis_scalar_111_tlast),
        .m_axis_scalar_111_tvalid(m_axis_scalar_111_tvalid),
        .m_axis_scalar_111_tkeep(m_axis_scalar_111_tkeep),
        .m_axis_scalar_111_tstrb(m_axis_scalar_111_tstrb),
        .m_axis_scalar_111_tdata(m_axis_scalar_111_tdata),
        .m_axis_scalar_111_tready(m_axis_scalar_111_tready),
        .m_axis_scalar_112_aclk(m_axis_scalar_112_aclk),
        .m_axis_scalar_112_aresetn(m_axis_scalar_112_aresetn),
        .m_axis_scalar_112_tlast(m_axis_scalar_112_tlast),
        .m_axis_scalar_112_tvalid(m_axis_scalar_112_tvalid),
        .m_axis_scalar_112_tkeep(m_axis_scalar_112_tkeep),
        .m_axis_scalar_112_tstrb(m_axis_scalar_112_tstrb),
        .m_axis_scalar_112_tdata(m_axis_scalar_112_tdata),
        .m_axis_scalar_112_tready(m_axis_scalar_112_tready),
        .m_axis_scalar_113_aclk(m_axis_scalar_113_aclk),
        .m_axis_scalar_113_aresetn(m_axis_scalar_113_aresetn),
        .m_axis_scalar_113_tlast(m_axis_scalar_113_tlast),
        .m_axis_scalar_113_tvalid(m_axis_scalar_113_tvalid),
        .m_axis_scalar_113_tkeep(m_axis_scalar_113_tkeep),
        .m_axis_scalar_113_tstrb(m_axis_scalar_113_tstrb),
        .m_axis_scalar_113_tdata(m_axis_scalar_113_tdata),
        .m_axis_scalar_113_tready(m_axis_scalar_113_tready),
        .m_axis_scalar_114_aclk(m_axis_scalar_114_aclk),
        .m_axis_scalar_114_aresetn(m_axis_scalar_114_aresetn),
        .m_axis_scalar_114_tlast(m_axis_scalar_114_tlast),
        .m_axis_scalar_114_tvalid(m_axis_scalar_114_tvalid),
        .m_axis_scalar_114_tkeep(m_axis_scalar_114_tkeep),
        .m_axis_scalar_114_tstrb(m_axis_scalar_114_tstrb),
        .m_axis_scalar_114_tdata(m_axis_scalar_114_tdata),
        .m_axis_scalar_114_tready(m_axis_scalar_114_tready),
        .m_axis_scalar_115_aclk(m_axis_scalar_115_aclk),
        .m_axis_scalar_115_aresetn(m_axis_scalar_115_aresetn),
        .m_axis_scalar_115_tlast(m_axis_scalar_115_tlast),
        .m_axis_scalar_115_tvalid(m_axis_scalar_115_tvalid),
        .m_axis_scalar_115_tkeep(m_axis_scalar_115_tkeep),
        .m_axis_scalar_115_tstrb(m_axis_scalar_115_tstrb),
        .m_axis_scalar_115_tdata(m_axis_scalar_115_tdata),
        .m_axis_scalar_115_tready(m_axis_scalar_115_tready),
        .m_axis_scalar_116_aclk(m_axis_scalar_116_aclk),
        .m_axis_scalar_116_aresetn(m_axis_scalar_116_aresetn),
        .m_axis_scalar_116_tlast(m_axis_scalar_116_tlast),
        .m_axis_scalar_116_tvalid(m_axis_scalar_116_tvalid),
        .m_axis_scalar_116_tkeep(m_axis_scalar_116_tkeep),
        .m_axis_scalar_116_tstrb(m_axis_scalar_116_tstrb),
        .m_axis_scalar_116_tdata(m_axis_scalar_116_tdata),
        .m_axis_scalar_116_tready(m_axis_scalar_116_tready),
        .m_axis_scalar_117_aclk(m_axis_scalar_117_aclk),
        .m_axis_scalar_117_aresetn(m_axis_scalar_117_aresetn),
        .m_axis_scalar_117_tlast(m_axis_scalar_117_tlast),
        .m_axis_scalar_117_tvalid(m_axis_scalar_117_tvalid),
        .m_axis_scalar_117_tkeep(m_axis_scalar_117_tkeep),
        .m_axis_scalar_117_tstrb(m_axis_scalar_117_tstrb),
        .m_axis_scalar_117_tdata(m_axis_scalar_117_tdata),
        .m_axis_scalar_117_tready(m_axis_scalar_117_tready),
        .m_axis_scalar_118_aclk(m_axis_scalar_118_aclk),
        .m_axis_scalar_118_aresetn(m_axis_scalar_118_aresetn),
        .m_axis_scalar_118_tlast(m_axis_scalar_118_tlast),
        .m_axis_scalar_118_tvalid(m_axis_scalar_118_tvalid),
        .m_axis_scalar_118_tkeep(m_axis_scalar_118_tkeep),
        .m_axis_scalar_118_tstrb(m_axis_scalar_118_tstrb),
        .m_axis_scalar_118_tdata(m_axis_scalar_118_tdata),
        .m_axis_scalar_118_tready(m_axis_scalar_118_tready),
        .m_axis_scalar_119_aclk(m_axis_scalar_119_aclk),
        .m_axis_scalar_119_aresetn(m_axis_scalar_119_aresetn),
        .m_axis_scalar_119_tlast(m_axis_scalar_119_tlast),
        .m_axis_scalar_119_tvalid(m_axis_scalar_119_tvalid),
        .m_axis_scalar_119_tkeep(m_axis_scalar_119_tkeep),
        .m_axis_scalar_119_tstrb(m_axis_scalar_119_tstrb),
        .m_axis_scalar_119_tdata(m_axis_scalar_119_tdata),
        .m_axis_scalar_119_tready(m_axis_scalar_119_tready),
        .m_axis_scalar_120_aclk(m_axis_scalar_120_aclk),
        .m_axis_scalar_120_aresetn(m_axis_scalar_120_aresetn),
        .m_axis_scalar_120_tlast(m_axis_scalar_120_tlast),
        .m_axis_scalar_120_tvalid(m_axis_scalar_120_tvalid),
        .m_axis_scalar_120_tkeep(m_axis_scalar_120_tkeep),
        .m_axis_scalar_120_tstrb(m_axis_scalar_120_tstrb),
        .m_axis_scalar_120_tdata(m_axis_scalar_120_tdata),
        .m_axis_scalar_120_tready(m_axis_scalar_120_tready),
        .m_axis_scalar_121_aclk(m_axis_scalar_121_aclk),
        .m_axis_scalar_121_aresetn(m_axis_scalar_121_aresetn),
        .m_axis_scalar_121_tlast(m_axis_scalar_121_tlast),
        .m_axis_scalar_121_tvalid(m_axis_scalar_121_tvalid),
        .m_axis_scalar_121_tkeep(m_axis_scalar_121_tkeep),
        .m_axis_scalar_121_tstrb(m_axis_scalar_121_tstrb),
        .m_axis_scalar_121_tdata(m_axis_scalar_121_tdata),
        .m_axis_scalar_121_tready(m_axis_scalar_121_tready),
        .m_axis_scalar_122_aclk(m_axis_scalar_122_aclk),
        .m_axis_scalar_122_aresetn(m_axis_scalar_122_aresetn),
        .m_axis_scalar_122_tlast(m_axis_scalar_122_tlast),
        .m_axis_scalar_122_tvalid(m_axis_scalar_122_tvalid),
        .m_axis_scalar_122_tkeep(m_axis_scalar_122_tkeep),
        .m_axis_scalar_122_tstrb(m_axis_scalar_122_tstrb),
        .m_axis_scalar_122_tdata(m_axis_scalar_122_tdata),
        .m_axis_scalar_122_tready(m_axis_scalar_122_tready),
        .m_axis_scalar_123_aclk(m_axis_scalar_123_aclk),
        .m_axis_scalar_123_aresetn(m_axis_scalar_123_aresetn),
        .m_axis_scalar_123_tlast(m_axis_scalar_123_tlast),
        .m_axis_scalar_123_tvalid(m_axis_scalar_123_tvalid),
        .m_axis_scalar_123_tkeep(m_axis_scalar_123_tkeep),
        .m_axis_scalar_123_tstrb(m_axis_scalar_123_tstrb),
        .m_axis_scalar_123_tdata(m_axis_scalar_123_tdata),
        .m_axis_scalar_123_tready(m_axis_scalar_123_tready),
        .m_axis_scalar_124_aclk(m_axis_scalar_124_aclk),
        .m_axis_scalar_124_aresetn(m_axis_scalar_124_aresetn),
        .m_axis_scalar_124_tlast(m_axis_scalar_124_tlast),
        .m_axis_scalar_124_tvalid(m_axis_scalar_124_tvalid),
        .m_axis_scalar_124_tkeep(m_axis_scalar_124_tkeep),
        .m_axis_scalar_124_tstrb(m_axis_scalar_124_tstrb),
        .m_axis_scalar_124_tdata(m_axis_scalar_124_tdata),
        .m_axis_scalar_124_tready(m_axis_scalar_124_tready),
        .m_axis_scalar_125_aclk(m_axis_scalar_125_aclk),
        .m_axis_scalar_125_aresetn(m_axis_scalar_125_aresetn),
        .m_axis_scalar_125_tlast(m_axis_scalar_125_tlast),
        .m_axis_scalar_125_tvalid(m_axis_scalar_125_tvalid),
        .m_axis_scalar_125_tkeep(m_axis_scalar_125_tkeep),
        .m_axis_scalar_125_tstrb(m_axis_scalar_125_tstrb),
        .m_axis_scalar_125_tdata(m_axis_scalar_125_tdata),
        .m_axis_scalar_125_tready(m_axis_scalar_125_tready),
        .m_axis_scalar_126_aclk(m_axis_scalar_126_aclk),
        .m_axis_scalar_126_aresetn(m_axis_scalar_126_aresetn),
        .m_axis_scalar_126_tlast(m_axis_scalar_126_tlast),
        .m_axis_scalar_126_tvalid(m_axis_scalar_126_tvalid),
        .m_axis_scalar_126_tkeep(m_axis_scalar_126_tkeep),
        .m_axis_scalar_126_tstrb(m_axis_scalar_126_tstrb),
        .m_axis_scalar_126_tdata(m_axis_scalar_126_tdata),
        .m_axis_scalar_126_tready(m_axis_scalar_126_tready),
        .m_axis_scalar_127_aclk(m_axis_scalar_127_aclk),
        .m_axis_scalar_127_aresetn(m_axis_scalar_127_aresetn),
        .m_axis_scalar_127_tlast(m_axis_scalar_127_tlast),
        .m_axis_scalar_127_tvalid(m_axis_scalar_127_tvalid),
        .m_axis_scalar_127_tkeep(m_axis_scalar_127_tkeep),
        .m_axis_scalar_127_tstrb(m_axis_scalar_127_tstrb),
        .m_axis_scalar_127_tdata(m_axis_scalar_127_tdata),
        .m_axis_scalar_127_tready(m_axis_scalar_127_tready)
    );
    
    in_fifo_args #(
        .C_NUM_INPUT_FIFOs(C_NUM_INPUT_FIFOs),
        .S_AXIS_FIFO_0_WIDTH(S_AXIS_FIFO_0_WIDTH),
        .S_AXIS_FIFO_1_WIDTH(S_AXIS_FIFO_1_WIDTH),
        .S_AXIS_FIFO_2_WIDTH(S_AXIS_FIFO_2_WIDTH),
        .S_AXIS_FIFO_3_WIDTH(S_AXIS_FIFO_3_WIDTH),
        .S_AXIS_FIFO_4_WIDTH(S_AXIS_FIFO_4_WIDTH),
        .S_AXIS_FIFO_5_WIDTH(S_AXIS_FIFO_5_WIDTH),
        .S_AXIS_FIFO_6_WIDTH(S_AXIS_FIFO_6_WIDTH),
        .S_AXIS_FIFO_7_WIDTH(S_AXIS_FIFO_7_WIDTH),
        .S_AXIS_FIFO_8_WIDTH(S_AXIS_FIFO_8_WIDTH),
        .S_AXIS_FIFO_9_WIDTH(S_AXIS_FIFO_9_WIDTH),
        .S_AXIS_FIFO_10_WIDTH(S_AXIS_FIFO_10_WIDTH),
        .S_AXIS_FIFO_11_WIDTH(S_AXIS_FIFO_11_WIDTH),
        .S_AXIS_FIFO_12_WIDTH(S_AXIS_FIFO_12_WIDTH),
        .S_AXIS_FIFO_13_WIDTH(S_AXIS_FIFO_13_WIDTH),
        .S_AXIS_FIFO_14_WIDTH(S_AXIS_FIFO_14_WIDTH),
        .S_AXIS_FIFO_15_WIDTH(S_AXIS_FIFO_15_WIDTH),
        .S_AXIS_FIFO_16_WIDTH(S_AXIS_FIFO_16_WIDTH),
        .S_AXIS_FIFO_17_WIDTH(S_AXIS_FIFO_17_WIDTH),
        .S_AXIS_FIFO_18_WIDTH(S_AXIS_FIFO_18_WIDTH),
        .S_AXIS_FIFO_19_WIDTH(S_AXIS_FIFO_19_WIDTH),
        .S_AXIS_FIFO_20_WIDTH(S_AXIS_FIFO_20_WIDTH),
        .S_AXIS_FIFO_21_WIDTH(S_AXIS_FIFO_21_WIDTH),
        .S_AXIS_FIFO_22_WIDTH(S_AXIS_FIFO_22_WIDTH),
        .S_AXIS_FIFO_23_WIDTH(S_AXIS_FIFO_23_WIDTH),
        .S_AXIS_FIFO_24_WIDTH(S_AXIS_FIFO_24_WIDTH),
        .S_AXIS_FIFO_25_WIDTH(S_AXIS_FIFO_25_WIDTH),
        .S_AXIS_FIFO_26_WIDTH(S_AXIS_FIFO_26_WIDTH),
        .S_AXIS_FIFO_27_WIDTH(S_AXIS_FIFO_27_WIDTH),
        .S_AXIS_FIFO_28_WIDTH(S_AXIS_FIFO_28_WIDTH),
        .S_AXIS_FIFO_29_WIDTH(S_AXIS_FIFO_29_WIDTH),
        .S_AXIS_FIFO_30_WIDTH(S_AXIS_FIFO_30_WIDTH),
        .S_AXIS_FIFO_31_WIDTH(S_AXIS_FIFO_31_WIDTH),
        .S_AXIS_FIFO_32_WIDTH(S_AXIS_FIFO_32_WIDTH),
        .S_AXIS_FIFO_33_WIDTH(S_AXIS_FIFO_33_WIDTH),
        .S_AXIS_FIFO_34_WIDTH(S_AXIS_FIFO_34_WIDTH),
        .S_AXIS_FIFO_35_WIDTH(S_AXIS_FIFO_35_WIDTH),
        .S_AXIS_FIFO_36_WIDTH(S_AXIS_FIFO_36_WIDTH),
        .S_AXIS_FIFO_37_WIDTH(S_AXIS_FIFO_37_WIDTH),
        .S_AXIS_FIFO_38_WIDTH(S_AXIS_FIFO_38_WIDTH),
        .S_AXIS_FIFO_39_WIDTH(S_AXIS_FIFO_39_WIDTH),
        .S_AXIS_FIFO_40_WIDTH(S_AXIS_FIFO_40_WIDTH),
        .S_AXIS_FIFO_41_WIDTH(S_AXIS_FIFO_41_WIDTH),
        .S_AXIS_FIFO_42_WIDTH(S_AXIS_FIFO_42_WIDTH),
        .S_AXIS_FIFO_43_WIDTH(S_AXIS_FIFO_43_WIDTH),
        .S_AXIS_FIFO_44_WIDTH(S_AXIS_FIFO_44_WIDTH),
        .S_AXIS_FIFO_45_WIDTH(S_AXIS_FIFO_45_WIDTH),
        .S_AXIS_FIFO_46_WIDTH(S_AXIS_FIFO_46_WIDTH),
        .S_AXIS_FIFO_47_WIDTH(S_AXIS_FIFO_47_WIDTH),
        .S_AXIS_FIFO_48_WIDTH(S_AXIS_FIFO_48_WIDTH),
        .S_AXIS_FIFO_49_WIDTH(S_AXIS_FIFO_49_WIDTH),
        .S_AXIS_FIFO_50_WIDTH(S_AXIS_FIFO_50_WIDTH),
        .S_AXIS_FIFO_51_WIDTH(S_AXIS_FIFO_51_WIDTH),
        .S_AXIS_FIFO_52_WIDTH(S_AXIS_FIFO_52_WIDTH),
        .S_AXIS_FIFO_53_WIDTH(S_AXIS_FIFO_53_WIDTH),
        .S_AXIS_FIFO_54_WIDTH(S_AXIS_FIFO_54_WIDTH),
        .S_AXIS_FIFO_55_WIDTH(S_AXIS_FIFO_55_WIDTH),
        .S_AXIS_FIFO_56_WIDTH(S_AXIS_FIFO_56_WIDTH),
        .S_AXIS_FIFO_57_WIDTH(S_AXIS_FIFO_57_WIDTH),
        .S_AXIS_FIFO_58_WIDTH(S_AXIS_FIFO_58_WIDTH),
        .S_AXIS_FIFO_59_WIDTH(S_AXIS_FIFO_59_WIDTH),
        .S_AXIS_FIFO_60_WIDTH(S_AXIS_FIFO_60_WIDTH),
        .S_AXIS_FIFO_61_WIDTH(S_AXIS_FIFO_61_WIDTH),
        .S_AXIS_FIFO_62_WIDTH(S_AXIS_FIFO_62_WIDTH),
        .S_AXIS_FIFO_63_WIDTH(S_AXIS_FIFO_63_WIDTH),
        .S_AXIS_FIFO_64_WIDTH(S_AXIS_FIFO_64_WIDTH),
        .S_AXIS_FIFO_65_WIDTH(S_AXIS_FIFO_65_WIDTH),
        .S_AXIS_FIFO_66_WIDTH(S_AXIS_FIFO_66_WIDTH),
        .S_AXIS_FIFO_67_WIDTH(S_AXIS_FIFO_67_WIDTH),
        .S_AXIS_FIFO_68_WIDTH(S_AXIS_FIFO_68_WIDTH),
        .S_AXIS_FIFO_69_WIDTH(S_AXIS_FIFO_69_WIDTH),
        .S_AXIS_FIFO_70_WIDTH(S_AXIS_FIFO_70_WIDTH),
        .S_AXIS_FIFO_71_WIDTH(S_AXIS_FIFO_71_WIDTH),
        .S_AXIS_FIFO_72_WIDTH(S_AXIS_FIFO_72_WIDTH),
        .S_AXIS_FIFO_73_WIDTH(S_AXIS_FIFO_73_WIDTH),
        .S_AXIS_FIFO_74_WIDTH(S_AXIS_FIFO_74_WIDTH),
        .S_AXIS_FIFO_75_WIDTH(S_AXIS_FIFO_75_WIDTH),
        .S_AXIS_FIFO_76_WIDTH(S_AXIS_FIFO_76_WIDTH),
        .S_AXIS_FIFO_77_WIDTH(S_AXIS_FIFO_77_WIDTH),
        .S_AXIS_FIFO_78_WIDTH(S_AXIS_FIFO_78_WIDTH),
        .S_AXIS_FIFO_79_WIDTH(S_AXIS_FIFO_79_WIDTH),
        .S_AXIS_FIFO_80_WIDTH(S_AXIS_FIFO_80_WIDTH),
        .S_AXIS_FIFO_81_WIDTH(S_AXIS_FIFO_81_WIDTH),
        .S_AXIS_FIFO_82_WIDTH(S_AXIS_FIFO_82_WIDTH),
        .S_AXIS_FIFO_83_WIDTH(S_AXIS_FIFO_83_WIDTH),
        .S_AXIS_FIFO_84_WIDTH(S_AXIS_FIFO_84_WIDTH),
        .S_AXIS_FIFO_85_WIDTH(S_AXIS_FIFO_85_WIDTH),
        .S_AXIS_FIFO_86_WIDTH(S_AXIS_FIFO_86_WIDTH),
        .S_AXIS_FIFO_87_WIDTH(S_AXIS_FIFO_87_WIDTH),
        .S_AXIS_FIFO_88_WIDTH(S_AXIS_FIFO_88_WIDTH),
        .S_AXIS_FIFO_89_WIDTH(S_AXIS_FIFO_89_WIDTH),
        .S_AXIS_FIFO_90_WIDTH(S_AXIS_FIFO_90_WIDTH),
        .S_AXIS_FIFO_91_WIDTH(S_AXIS_FIFO_91_WIDTH),
        .S_AXIS_FIFO_92_WIDTH(S_AXIS_FIFO_92_WIDTH),
        .S_AXIS_FIFO_93_WIDTH(S_AXIS_FIFO_93_WIDTH),
        .S_AXIS_FIFO_94_WIDTH(S_AXIS_FIFO_94_WIDTH),
        .S_AXIS_FIFO_95_WIDTH(S_AXIS_FIFO_95_WIDTH),
        .S_AXIS_FIFO_96_WIDTH(S_AXIS_FIFO_96_WIDTH),
        .S_AXIS_FIFO_97_WIDTH(S_AXIS_FIFO_97_WIDTH),
        .S_AXIS_FIFO_98_WIDTH(S_AXIS_FIFO_98_WIDTH),
        .S_AXIS_FIFO_99_WIDTH(S_AXIS_FIFO_99_WIDTH),
        .S_AXIS_FIFO_100_WIDTH(S_AXIS_FIFO_100_WIDTH),
        .S_AXIS_FIFO_101_WIDTH(S_AXIS_FIFO_101_WIDTH),
        .S_AXIS_FIFO_102_WIDTH(S_AXIS_FIFO_102_WIDTH),
        .S_AXIS_FIFO_103_WIDTH(S_AXIS_FIFO_103_WIDTH),
        .S_AXIS_FIFO_104_WIDTH(S_AXIS_FIFO_104_WIDTH),
        .S_AXIS_FIFO_105_WIDTH(S_AXIS_FIFO_105_WIDTH),
        .S_AXIS_FIFO_106_WIDTH(S_AXIS_FIFO_106_WIDTH),
        .S_AXIS_FIFO_107_WIDTH(S_AXIS_FIFO_107_WIDTH),
        .S_AXIS_FIFO_108_WIDTH(S_AXIS_FIFO_108_WIDTH),
        .S_AXIS_FIFO_109_WIDTH(S_AXIS_FIFO_109_WIDTH),
        .S_AXIS_FIFO_110_WIDTH(S_AXIS_FIFO_110_WIDTH),
        .S_AXIS_FIFO_111_WIDTH(S_AXIS_FIFO_111_WIDTH),
        .S_AXIS_FIFO_112_WIDTH(S_AXIS_FIFO_112_WIDTH),
        .S_AXIS_FIFO_113_WIDTH(S_AXIS_FIFO_113_WIDTH),
        .S_AXIS_FIFO_114_WIDTH(S_AXIS_FIFO_114_WIDTH),
        .S_AXIS_FIFO_115_WIDTH(S_AXIS_FIFO_115_WIDTH),
        .S_AXIS_FIFO_116_WIDTH(S_AXIS_FIFO_116_WIDTH),
        .S_AXIS_FIFO_117_WIDTH(S_AXIS_FIFO_117_WIDTH),
        .S_AXIS_FIFO_118_WIDTH(S_AXIS_FIFO_118_WIDTH),
        .S_AXIS_FIFO_119_WIDTH(S_AXIS_FIFO_119_WIDTH),
        .S_AXIS_FIFO_120_WIDTH(S_AXIS_FIFO_120_WIDTH),
        .S_AXIS_FIFO_121_WIDTH(S_AXIS_FIFO_121_WIDTH),
        .S_AXIS_FIFO_122_WIDTH(S_AXIS_FIFO_122_WIDTH),
        .S_AXIS_FIFO_123_WIDTH(S_AXIS_FIFO_123_WIDTH),
        .S_AXIS_FIFO_124_WIDTH(S_AXIS_FIFO_124_WIDTH),
        .S_AXIS_FIFO_125_WIDTH(S_AXIS_FIFO_125_WIDTH),
        .S_AXIS_FIFO_126_WIDTH(S_AXIS_FIFO_126_WIDTH),
        .S_AXIS_FIFO_127_WIDTH(S_AXIS_FIFO_127_WIDTH),
        .S_AXIS_FIFO_0_DEPTH(S_AXIS_FIFO_0_DEPTH),
        .S_AXIS_FIFO_1_DEPTH(S_AXIS_FIFO_1_DEPTH),
        .S_AXIS_FIFO_2_DEPTH(S_AXIS_FIFO_2_DEPTH),
        .S_AXIS_FIFO_3_DEPTH(S_AXIS_FIFO_3_DEPTH),
        .S_AXIS_FIFO_4_DEPTH(S_AXIS_FIFO_4_DEPTH),
        .S_AXIS_FIFO_5_DEPTH(S_AXIS_FIFO_5_DEPTH),
        .S_AXIS_FIFO_6_DEPTH(S_AXIS_FIFO_6_DEPTH),
        .S_AXIS_FIFO_7_DEPTH(S_AXIS_FIFO_7_DEPTH),
        .S_AXIS_FIFO_8_DEPTH(S_AXIS_FIFO_8_DEPTH),
        .S_AXIS_FIFO_9_DEPTH(S_AXIS_FIFO_9_DEPTH),
        .S_AXIS_FIFO_10_DEPTH(S_AXIS_FIFO_10_DEPTH),
        .S_AXIS_FIFO_11_DEPTH(S_AXIS_FIFO_11_DEPTH),
        .S_AXIS_FIFO_12_DEPTH(S_AXIS_FIFO_12_DEPTH),
        .S_AXIS_FIFO_13_DEPTH(S_AXIS_FIFO_13_DEPTH),
        .S_AXIS_FIFO_14_DEPTH(S_AXIS_FIFO_14_DEPTH),
        .S_AXIS_FIFO_15_DEPTH(S_AXIS_FIFO_15_DEPTH),
        .S_AXIS_FIFO_16_DEPTH(S_AXIS_FIFO_16_DEPTH),
        .S_AXIS_FIFO_17_DEPTH(S_AXIS_FIFO_17_DEPTH),
        .S_AXIS_FIFO_18_DEPTH(S_AXIS_FIFO_18_DEPTH),
        .S_AXIS_FIFO_19_DEPTH(S_AXIS_FIFO_19_DEPTH),
        .S_AXIS_FIFO_20_DEPTH(S_AXIS_FIFO_20_DEPTH),
        .S_AXIS_FIFO_21_DEPTH(S_AXIS_FIFO_21_DEPTH),
        .S_AXIS_FIFO_22_DEPTH(S_AXIS_FIFO_22_DEPTH),
        .S_AXIS_FIFO_23_DEPTH(S_AXIS_FIFO_23_DEPTH),
        .S_AXIS_FIFO_24_DEPTH(S_AXIS_FIFO_24_DEPTH),
        .S_AXIS_FIFO_25_DEPTH(S_AXIS_FIFO_25_DEPTH),
        .S_AXIS_FIFO_26_DEPTH(S_AXIS_FIFO_26_DEPTH),
        .S_AXIS_FIFO_27_DEPTH(S_AXIS_FIFO_27_DEPTH),
        .S_AXIS_FIFO_28_DEPTH(S_AXIS_FIFO_28_DEPTH),
        .S_AXIS_FIFO_29_DEPTH(S_AXIS_FIFO_29_DEPTH),
        .S_AXIS_FIFO_30_DEPTH(S_AXIS_FIFO_30_DEPTH),
        .S_AXIS_FIFO_31_DEPTH(S_AXIS_FIFO_31_DEPTH),
        .S_AXIS_FIFO_32_DEPTH(S_AXIS_FIFO_32_DEPTH),
        .S_AXIS_FIFO_33_DEPTH(S_AXIS_FIFO_33_DEPTH),
        .S_AXIS_FIFO_34_DEPTH(S_AXIS_FIFO_34_DEPTH),
        .S_AXIS_FIFO_35_DEPTH(S_AXIS_FIFO_35_DEPTH),
        .S_AXIS_FIFO_36_DEPTH(S_AXIS_FIFO_36_DEPTH),
        .S_AXIS_FIFO_37_DEPTH(S_AXIS_FIFO_37_DEPTH),
        .S_AXIS_FIFO_38_DEPTH(S_AXIS_FIFO_38_DEPTH),
        .S_AXIS_FIFO_39_DEPTH(S_AXIS_FIFO_39_DEPTH),
        .S_AXIS_FIFO_40_DEPTH(S_AXIS_FIFO_40_DEPTH),
        .S_AXIS_FIFO_41_DEPTH(S_AXIS_FIFO_41_DEPTH),
        .S_AXIS_FIFO_42_DEPTH(S_AXIS_FIFO_42_DEPTH),
        .S_AXIS_FIFO_43_DEPTH(S_AXIS_FIFO_43_DEPTH),
        .S_AXIS_FIFO_44_DEPTH(S_AXIS_FIFO_44_DEPTH),
        .S_AXIS_FIFO_45_DEPTH(S_AXIS_FIFO_45_DEPTH),
        .S_AXIS_FIFO_46_DEPTH(S_AXIS_FIFO_46_DEPTH),
        .S_AXIS_FIFO_47_DEPTH(S_AXIS_FIFO_47_DEPTH),
        .S_AXIS_FIFO_48_DEPTH(S_AXIS_FIFO_48_DEPTH),
        .S_AXIS_FIFO_49_DEPTH(S_AXIS_FIFO_49_DEPTH),
        .S_AXIS_FIFO_50_DEPTH(S_AXIS_FIFO_50_DEPTH),
        .S_AXIS_FIFO_51_DEPTH(S_AXIS_FIFO_51_DEPTH),
        .S_AXIS_FIFO_52_DEPTH(S_AXIS_FIFO_52_DEPTH),
        .S_AXIS_FIFO_53_DEPTH(S_AXIS_FIFO_53_DEPTH),
        .S_AXIS_FIFO_54_DEPTH(S_AXIS_FIFO_54_DEPTH),
        .S_AXIS_FIFO_55_DEPTH(S_AXIS_FIFO_55_DEPTH),
        .S_AXIS_FIFO_56_DEPTH(S_AXIS_FIFO_56_DEPTH),
        .S_AXIS_FIFO_57_DEPTH(S_AXIS_FIFO_57_DEPTH),
        .S_AXIS_FIFO_58_DEPTH(S_AXIS_FIFO_58_DEPTH),
        .S_AXIS_FIFO_59_DEPTH(S_AXIS_FIFO_59_DEPTH),
        .S_AXIS_FIFO_60_DEPTH(S_AXIS_FIFO_60_DEPTH),
        .S_AXIS_FIFO_61_DEPTH(S_AXIS_FIFO_61_DEPTH),
        .S_AXIS_FIFO_62_DEPTH(S_AXIS_FIFO_62_DEPTH),
        .S_AXIS_FIFO_63_DEPTH(S_AXIS_FIFO_63_DEPTH),
        .S_AXIS_FIFO_64_DEPTH(S_AXIS_FIFO_64_DEPTH),
        .S_AXIS_FIFO_65_DEPTH(S_AXIS_FIFO_65_DEPTH),
        .S_AXIS_FIFO_66_DEPTH(S_AXIS_FIFO_66_DEPTH),
        .S_AXIS_FIFO_67_DEPTH(S_AXIS_FIFO_67_DEPTH),
        .S_AXIS_FIFO_68_DEPTH(S_AXIS_FIFO_68_DEPTH),
        .S_AXIS_FIFO_69_DEPTH(S_AXIS_FIFO_69_DEPTH),
        .S_AXIS_FIFO_70_DEPTH(S_AXIS_FIFO_70_DEPTH),
        .S_AXIS_FIFO_71_DEPTH(S_AXIS_FIFO_71_DEPTH),
        .S_AXIS_FIFO_72_DEPTH(S_AXIS_FIFO_72_DEPTH),
        .S_AXIS_FIFO_73_DEPTH(S_AXIS_FIFO_73_DEPTH),
        .S_AXIS_FIFO_74_DEPTH(S_AXIS_FIFO_74_DEPTH),
        .S_AXIS_FIFO_75_DEPTH(S_AXIS_FIFO_75_DEPTH),
        .S_AXIS_FIFO_76_DEPTH(S_AXIS_FIFO_76_DEPTH),
        .S_AXIS_FIFO_77_DEPTH(S_AXIS_FIFO_77_DEPTH),
        .S_AXIS_FIFO_78_DEPTH(S_AXIS_FIFO_78_DEPTH),
        .S_AXIS_FIFO_79_DEPTH(S_AXIS_FIFO_79_DEPTH),
        .S_AXIS_FIFO_80_DEPTH(S_AXIS_FIFO_80_DEPTH),
        .S_AXIS_FIFO_81_DEPTH(S_AXIS_FIFO_81_DEPTH),
        .S_AXIS_FIFO_82_DEPTH(S_AXIS_FIFO_82_DEPTH),
        .S_AXIS_FIFO_83_DEPTH(S_AXIS_FIFO_83_DEPTH),
        .S_AXIS_FIFO_84_DEPTH(S_AXIS_FIFO_84_DEPTH),
        .S_AXIS_FIFO_85_DEPTH(S_AXIS_FIFO_85_DEPTH),
        .S_AXIS_FIFO_86_DEPTH(S_AXIS_FIFO_86_DEPTH),
        .S_AXIS_FIFO_87_DEPTH(S_AXIS_FIFO_87_DEPTH),
        .S_AXIS_FIFO_88_DEPTH(S_AXIS_FIFO_88_DEPTH),
        .S_AXIS_FIFO_89_DEPTH(S_AXIS_FIFO_89_DEPTH),
        .S_AXIS_FIFO_90_DEPTH(S_AXIS_FIFO_90_DEPTH),
        .S_AXIS_FIFO_91_DEPTH(S_AXIS_FIFO_91_DEPTH),
        .S_AXIS_FIFO_92_DEPTH(S_AXIS_FIFO_92_DEPTH),
        .S_AXIS_FIFO_93_DEPTH(S_AXIS_FIFO_93_DEPTH),
        .S_AXIS_FIFO_94_DEPTH(S_AXIS_FIFO_94_DEPTH),
        .S_AXIS_FIFO_95_DEPTH(S_AXIS_FIFO_95_DEPTH),
        .S_AXIS_FIFO_96_DEPTH(S_AXIS_FIFO_96_DEPTH),
        .S_AXIS_FIFO_97_DEPTH(S_AXIS_FIFO_97_DEPTH),
        .S_AXIS_FIFO_98_DEPTH(S_AXIS_FIFO_98_DEPTH),
        .S_AXIS_FIFO_99_DEPTH(S_AXIS_FIFO_99_DEPTH),
        .S_AXIS_FIFO_100_DEPTH(S_AXIS_FIFO_100_DEPTH),
        .S_AXIS_FIFO_101_DEPTH(S_AXIS_FIFO_101_DEPTH),
        .S_AXIS_FIFO_102_DEPTH(S_AXIS_FIFO_102_DEPTH),
        .S_AXIS_FIFO_103_DEPTH(S_AXIS_FIFO_103_DEPTH),
        .S_AXIS_FIFO_104_DEPTH(S_AXIS_FIFO_104_DEPTH),
        .S_AXIS_FIFO_105_DEPTH(S_AXIS_FIFO_105_DEPTH),
        .S_AXIS_FIFO_106_DEPTH(S_AXIS_FIFO_106_DEPTH),
        .S_AXIS_FIFO_107_DEPTH(S_AXIS_FIFO_107_DEPTH),
        .S_AXIS_FIFO_108_DEPTH(S_AXIS_FIFO_108_DEPTH),
        .S_AXIS_FIFO_109_DEPTH(S_AXIS_FIFO_109_DEPTH),
        .S_AXIS_FIFO_110_DEPTH(S_AXIS_FIFO_110_DEPTH),
        .S_AXIS_FIFO_111_DEPTH(S_AXIS_FIFO_111_DEPTH),
        .S_AXIS_FIFO_112_DEPTH(S_AXIS_FIFO_112_DEPTH),
        .S_AXIS_FIFO_113_DEPTH(S_AXIS_FIFO_113_DEPTH),
        .S_AXIS_FIFO_114_DEPTH(S_AXIS_FIFO_114_DEPTH),
        .S_AXIS_FIFO_115_DEPTH(S_AXIS_FIFO_115_DEPTH),
        .S_AXIS_FIFO_116_DEPTH(S_AXIS_FIFO_116_DEPTH),
        .S_AXIS_FIFO_117_DEPTH(S_AXIS_FIFO_117_DEPTH),
        .S_AXIS_FIFO_118_DEPTH(S_AXIS_FIFO_118_DEPTH),
        .S_AXIS_FIFO_119_DEPTH(S_AXIS_FIFO_119_DEPTH),
        .S_AXIS_FIFO_120_DEPTH(S_AXIS_FIFO_120_DEPTH),
        .S_AXIS_FIFO_121_DEPTH(S_AXIS_FIFO_121_DEPTH),
        .S_AXIS_FIFO_122_DEPTH(S_AXIS_FIFO_122_DEPTH),
        .S_AXIS_FIFO_123_DEPTH(S_AXIS_FIFO_123_DEPTH),
        .S_AXIS_FIFO_124_DEPTH(S_AXIS_FIFO_124_DEPTH),
        .S_AXIS_FIFO_125_DEPTH(S_AXIS_FIFO_125_DEPTH),
        .S_AXIS_FIFO_126_DEPTH(S_AXIS_FIFO_126_DEPTH),
        .S_AXIS_FIFO_127_DEPTH(S_AXIS_FIFO_127_DEPTH),
        .S_AXIS_FIFO_0_IS_ASYNC(S_AXIS_FIFO_0_IS_ASYNC),
        .S_AXIS_FIFO_1_IS_ASYNC(S_AXIS_FIFO_1_IS_ASYNC),
        .S_AXIS_FIFO_2_IS_ASYNC(S_AXIS_FIFO_2_IS_ASYNC),
        .S_AXIS_FIFO_3_IS_ASYNC(S_AXIS_FIFO_3_IS_ASYNC),
        .S_AXIS_FIFO_4_IS_ASYNC(S_AXIS_FIFO_4_IS_ASYNC),
        .S_AXIS_FIFO_5_IS_ASYNC(S_AXIS_FIFO_5_IS_ASYNC),
        .S_AXIS_FIFO_6_IS_ASYNC(S_AXIS_FIFO_6_IS_ASYNC),
        .S_AXIS_FIFO_7_IS_ASYNC(S_AXIS_FIFO_7_IS_ASYNC),
        .S_AXIS_FIFO_8_IS_ASYNC(S_AXIS_FIFO_8_IS_ASYNC),
        .S_AXIS_FIFO_9_IS_ASYNC(S_AXIS_FIFO_9_IS_ASYNC),
        .S_AXIS_FIFO_10_IS_ASYNC(S_AXIS_FIFO_10_IS_ASYNC),
        .S_AXIS_FIFO_11_IS_ASYNC(S_AXIS_FIFO_11_IS_ASYNC),
        .S_AXIS_FIFO_12_IS_ASYNC(S_AXIS_FIFO_12_IS_ASYNC),
        .S_AXIS_FIFO_13_IS_ASYNC(S_AXIS_FIFO_13_IS_ASYNC),
        .S_AXIS_FIFO_14_IS_ASYNC(S_AXIS_FIFO_14_IS_ASYNC),
        .S_AXIS_FIFO_15_IS_ASYNC(S_AXIS_FIFO_15_IS_ASYNC),
        .S_AXIS_FIFO_16_IS_ASYNC(S_AXIS_FIFO_16_IS_ASYNC),
        .S_AXIS_FIFO_17_IS_ASYNC(S_AXIS_FIFO_17_IS_ASYNC),
        .S_AXIS_FIFO_18_IS_ASYNC(S_AXIS_FIFO_18_IS_ASYNC),
        .S_AXIS_FIFO_19_IS_ASYNC(S_AXIS_FIFO_19_IS_ASYNC),
        .S_AXIS_FIFO_20_IS_ASYNC(S_AXIS_FIFO_20_IS_ASYNC),
        .S_AXIS_FIFO_21_IS_ASYNC(S_AXIS_FIFO_21_IS_ASYNC),
        .S_AXIS_FIFO_22_IS_ASYNC(S_AXIS_FIFO_22_IS_ASYNC),
        .S_AXIS_FIFO_23_IS_ASYNC(S_AXIS_FIFO_23_IS_ASYNC),
        .S_AXIS_FIFO_24_IS_ASYNC(S_AXIS_FIFO_24_IS_ASYNC),
        .S_AXIS_FIFO_25_IS_ASYNC(S_AXIS_FIFO_25_IS_ASYNC),
        .S_AXIS_FIFO_26_IS_ASYNC(S_AXIS_FIFO_26_IS_ASYNC),
        .S_AXIS_FIFO_27_IS_ASYNC(S_AXIS_FIFO_27_IS_ASYNC),
        .S_AXIS_FIFO_28_IS_ASYNC(S_AXIS_FIFO_28_IS_ASYNC),
        .S_AXIS_FIFO_29_IS_ASYNC(S_AXIS_FIFO_29_IS_ASYNC),
        .S_AXIS_FIFO_30_IS_ASYNC(S_AXIS_FIFO_30_IS_ASYNC),
        .S_AXIS_FIFO_31_IS_ASYNC(S_AXIS_FIFO_31_IS_ASYNC),
        .S_AXIS_FIFO_32_IS_ASYNC(S_AXIS_FIFO_32_IS_ASYNC),
        .S_AXIS_FIFO_33_IS_ASYNC(S_AXIS_FIFO_33_IS_ASYNC),
        .S_AXIS_FIFO_34_IS_ASYNC(S_AXIS_FIFO_34_IS_ASYNC),
        .S_AXIS_FIFO_35_IS_ASYNC(S_AXIS_FIFO_35_IS_ASYNC),
        .S_AXIS_FIFO_36_IS_ASYNC(S_AXIS_FIFO_36_IS_ASYNC),
        .S_AXIS_FIFO_37_IS_ASYNC(S_AXIS_FIFO_37_IS_ASYNC),
        .S_AXIS_FIFO_38_IS_ASYNC(S_AXIS_FIFO_38_IS_ASYNC),
        .S_AXIS_FIFO_39_IS_ASYNC(S_AXIS_FIFO_39_IS_ASYNC),
        .S_AXIS_FIFO_40_IS_ASYNC(S_AXIS_FIFO_40_IS_ASYNC),
        .S_AXIS_FIFO_41_IS_ASYNC(S_AXIS_FIFO_41_IS_ASYNC),
        .S_AXIS_FIFO_42_IS_ASYNC(S_AXIS_FIFO_42_IS_ASYNC),
        .S_AXIS_FIFO_43_IS_ASYNC(S_AXIS_FIFO_43_IS_ASYNC),
        .S_AXIS_FIFO_44_IS_ASYNC(S_AXIS_FIFO_44_IS_ASYNC),
        .S_AXIS_FIFO_45_IS_ASYNC(S_AXIS_FIFO_45_IS_ASYNC),
        .S_AXIS_FIFO_46_IS_ASYNC(S_AXIS_FIFO_46_IS_ASYNC),
        .S_AXIS_FIFO_47_IS_ASYNC(S_AXIS_FIFO_47_IS_ASYNC),
        .S_AXIS_FIFO_48_IS_ASYNC(S_AXIS_FIFO_48_IS_ASYNC),
        .S_AXIS_FIFO_49_IS_ASYNC(S_AXIS_FIFO_49_IS_ASYNC),
        .S_AXIS_FIFO_50_IS_ASYNC(S_AXIS_FIFO_50_IS_ASYNC),
        .S_AXIS_FIFO_51_IS_ASYNC(S_AXIS_FIFO_51_IS_ASYNC),
        .S_AXIS_FIFO_52_IS_ASYNC(S_AXIS_FIFO_52_IS_ASYNC),
        .S_AXIS_FIFO_53_IS_ASYNC(S_AXIS_FIFO_53_IS_ASYNC),
        .S_AXIS_FIFO_54_IS_ASYNC(S_AXIS_FIFO_54_IS_ASYNC),
        .S_AXIS_FIFO_55_IS_ASYNC(S_AXIS_FIFO_55_IS_ASYNC),
        .S_AXIS_FIFO_56_IS_ASYNC(S_AXIS_FIFO_56_IS_ASYNC),
        .S_AXIS_FIFO_57_IS_ASYNC(S_AXIS_FIFO_57_IS_ASYNC),
        .S_AXIS_FIFO_58_IS_ASYNC(S_AXIS_FIFO_58_IS_ASYNC),
        .S_AXIS_FIFO_59_IS_ASYNC(S_AXIS_FIFO_59_IS_ASYNC),
        .S_AXIS_FIFO_60_IS_ASYNC(S_AXIS_FIFO_60_IS_ASYNC),
        .S_AXIS_FIFO_61_IS_ASYNC(S_AXIS_FIFO_61_IS_ASYNC),
        .S_AXIS_FIFO_62_IS_ASYNC(S_AXIS_FIFO_62_IS_ASYNC),
        .S_AXIS_FIFO_63_IS_ASYNC(S_AXIS_FIFO_63_IS_ASYNC),
        .S_AXIS_FIFO_64_IS_ASYNC(S_AXIS_FIFO_64_IS_ASYNC),
        .S_AXIS_FIFO_65_IS_ASYNC(S_AXIS_FIFO_65_IS_ASYNC),
        .S_AXIS_FIFO_66_IS_ASYNC(S_AXIS_FIFO_66_IS_ASYNC),
        .S_AXIS_FIFO_67_IS_ASYNC(S_AXIS_FIFO_67_IS_ASYNC),
        .S_AXIS_FIFO_68_IS_ASYNC(S_AXIS_FIFO_68_IS_ASYNC),
        .S_AXIS_FIFO_69_IS_ASYNC(S_AXIS_FIFO_69_IS_ASYNC),
        .S_AXIS_FIFO_70_IS_ASYNC(S_AXIS_FIFO_70_IS_ASYNC),
        .S_AXIS_FIFO_71_IS_ASYNC(S_AXIS_FIFO_71_IS_ASYNC),
        .S_AXIS_FIFO_72_IS_ASYNC(S_AXIS_FIFO_72_IS_ASYNC),
        .S_AXIS_FIFO_73_IS_ASYNC(S_AXIS_FIFO_73_IS_ASYNC),
        .S_AXIS_FIFO_74_IS_ASYNC(S_AXIS_FIFO_74_IS_ASYNC),
        .S_AXIS_FIFO_75_IS_ASYNC(S_AXIS_FIFO_75_IS_ASYNC),
        .S_AXIS_FIFO_76_IS_ASYNC(S_AXIS_FIFO_76_IS_ASYNC),
        .S_AXIS_FIFO_77_IS_ASYNC(S_AXIS_FIFO_77_IS_ASYNC),
        .S_AXIS_FIFO_78_IS_ASYNC(S_AXIS_FIFO_78_IS_ASYNC),
        .S_AXIS_FIFO_79_IS_ASYNC(S_AXIS_FIFO_79_IS_ASYNC),
        .S_AXIS_FIFO_80_IS_ASYNC(S_AXIS_FIFO_80_IS_ASYNC),
        .S_AXIS_FIFO_81_IS_ASYNC(S_AXIS_FIFO_81_IS_ASYNC),
        .S_AXIS_FIFO_82_IS_ASYNC(S_AXIS_FIFO_82_IS_ASYNC),
        .S_AXIS_FIFO_83_IS_ASYNC(S_AXIS_FIFO_83_IS_ASYNC),
        .S_AXIS_FIFO_84_IS_ASYNC(S_AXIS_FIFO_84_IS_ASYNC),
        .S_AXIS_FIFO_85_IS_ASYNC(S_AXIS_FIFO_85_IS_ASYNC),
        .S_AXIS_FIFO_86_IS_ASYNC(S_AXIS_FIFO_86_IS_ASYNC),
        .S_AXIS_FIFO_87_IS_ASYNC(S_AXIS_FIFO_87_IS_ASYNC),
        .S_AXIS_FIFO_88_IS_ASYNC(S_AXIS_FIFO_88_IS_ASYNC),
        .S_AXIS_FIFO_89_IS_ASYNC(S_AXIS_FIFO_89_IS_ASYNC),
        .S_AXIS_FIFO_90_IS_ASYNC(S_AXIS_FIFO_90_IS_ASYNC),
        .S_AXIS_FIFO_91_IS_ASYNC(S_AXIS_FIFO_91_IS_ASYNC),
        .S_AXIS_FIFO_92_IS_ASYNC(S_AXIS_FIFO_92_IS_ASYNC),
        .S_AXIS_FIFO_93_IS_ASYNC(S_AXIS_FIFO_93_IS_ASYNC),
        .S_AXIS_FIFO_94_IS_ASYNC(S_AXIS_FIFO_94_IS_ASYNC),
        .S_AXIS_FIFO_95_IS_ASYNC(S_AXIS_FIFO_95_IS_ASYNC),
        .S_AXIS_FIFO_96_IS_ASYNC(S_AXIS_FIFO_96_IS_ASYNC),
        .S_AXIS_FIFO_97_IS_ASYNC(S_AXIS_FIFO_97_IS_ASYNC),
        .S_AXIS_FIFO_98_IS_ASYNC(S_AXIS_FIFO_98_IS_ASYNC),
        .S_AXIS_FIFO_99_IS_ASYNC(S_AXIS_FIFO_99_IS_ASYNC),
        .S_AXIS_FIFO_100_IS_ASYNC(S_AXIS_FIFO_100_IS_ASYNC),
        .S_AXIS_FIFO_101_IS_ASYNC(S_AXIS_FIFO_101_IS_ASYNC),
        .S_AXIS_FIFO_102_IS_ASYNC(S_AXIS_FIFO_102_IS_ASYNC),
        .S_AXIS_FIFO_103_IS_ASYNC(S_AXIS_FIFO_103_IS_ASYNC),
        .S_AXIS_FIFO_104_IS_ASYNC(S_AXIS_FIFO_104_IS_ASYNC),
        .S_AXIS_FIFO_105_IS_ASYNC(S_AXIS_FIFO_105_IS_ASYNC),
        .S_AXIS_FIFO_106_IS_ASYNC(S_AXIS_FIFO_106_IS_ASYNC),
        .S_AXIS_FIFO_107_IS_ASYNC(S_AXIS_FIFO_107_IS_ASYNC),
        .S_AXIS_FIFO_108_IS_ASYNC(S_AXIS_FIFO_108_IS_ASYNC),
        .S_AXIS_FIFO_109_IS_ASYNC(S_AXIS_FIFO_109_IS_ASYNC),
        .S_AXIS_FIFO_110_IS_ASYNC(S_AXIS_FIFO_110_IS_ASYNC),
        .S_AXIS_FIFO_111_IS_ASYNC(S_AXIS_FIFO_111_IS_ASYNC),
        .S_AXIS_FIFO_112_IS_ASYNC(S_AXIS_FIFO_112_IS_ASYNC),
        .S_AXIS_FIFO_113_IS_ASYNC(S_AXIS_FIFO_113_IS_ASYNC),
        .S_AXIS_FIFO_114_IS_ASYNC(S_AXIS_FIFO_114_IS_ASYNC),
        .S_AXIS_FIFO_115_IS_ASYNC(S_AXIS_FIFO_115_IS_ASYNC),
        .S_AXIS_FIFO_116_IS_ASYNC(S_AXIS_FIFO_116_IS_ASYNC),
        .S_AXIS_FIFO_117_IS_ASYNC(S_AXIS_FIFO_117_IS_ASYNC),
        .S_AXIS_FIFO_118_IS_ASYNC(S_AXIS_FIFO_118_IS_ASYNC),
        .S_AXIS_FIFO_119_IS_ASYNC(S_AXIS_FIFO_119_IS_ASYNC),
        .S_AXIS_FIFO_120_IS_ASYNC(S_AXIS_FIFO_120_IS_ASYNC),
        .S_AXIS_FIFO_121_IS_ASYNC(S_AXIS_FIFO_121_IS_ASYNC),
        .S_AXIS_FIFO_122_IS_ASYNC(S_AXIS_FIFO_122_IS_ASYNC),
        .S_AXIS_FIFO_123_IS_ASYNC(S_AXIS_FIFO_123_IS_ASYNC),
        .S_AXIS_FIFO_124_IS_ASYNC(S_AXIS_FIFO_124_IS_ASYNC),
        .S_AXIS_FIFO_125_IS_ASYNC(S_AXIS_FIFO_125_IS_ASYNC),
        .S_AXIS_FIFO_126_IS_ASYNC(S_AXIS_FIFO_126_IS_ASYNC),
        .S_AXIS_FIFO_127_IS_ASYNC(S_AXIS_FIFO_127_IS_ASYNC),
        .S_AXIS_FIFO_0_BYTE_WIDTH(S_AXIS_FIFO_0_BYTE_WIDTH),
        .S_AXIS_FIFO_1_BYTE_WIDTH(S_AXIS_FIFO_1_BYTE_WIDTH),
        .S_AXIS_FIFO_2_BYTE_WIDTH(S_AXIS_FIFO_2_BYTE_WIDTH),
        .S_AXIS_FIFO_3_BYTE_WIDTH(S_AXIS_FIFO_3_BYTE_WIDTH),
        .S_AXIS_FIFO_4_BYTE_WIDTH(S_AXIS_FIFO_4_BYTE_WIDTH),
        .S_AXIS_FIFO_5_BYTE_WIDTH(S_AXIS_FIFO_5_BYTE_WIDTH),
        .S_AXIS_FIFO_6_BYTE_WIDTH(S_AXIS_FIFO_6_BYTE_WIDTH),
        .S_AXIS_FIFO_7_BYTE_WIDTH(S_AXIS_FIFO_7_BYTE_WIDTH),
        .S_AXIS_FIFO_8_BYTE_WIDTH(S_AXIS_FIFO_8_BYTE_WIDTH),
        .S_AXIS_FIFO_9_BYTE_WIDTH(S_AXIS_FIFO_9_BYTE_WIDTH),
        .S_AXIS_FIFO_10_BYTE_WIDTH(S_AXIS_FIFO_10_BYTE_WIDTH),
        .S_AXIS_FIFO_11_BYTE_WIDTH(S_AXIS_FIFO_11_BYTE_WIDTH),
        .S_AXIS_FIFO_12_BYTE_WIDTH(S_AXIS_FIFO_12_BYTE_WIDTH),
        .S_AXIS_FIFO_13_BYTE_WIDTH(S_AXIS_FIFO_13_BYTE_WIDTH),
        .S_AXIS_FIFO_14_BYTE_WIDTH(S_AXIS_FIFO_14_BYTE_WIDTH),
        .S_AXIS_FIFO_15_BYTE_WIDTH(S_AXIS_FIFO_15_BYTE_WIDTH),
        .S_AXIS_FIFO_16_BYTE_WIDTH(S_AXIS_FIFO_16_BYTE_WIDTH),
        .S_AXIS_FIFO_17_BYTE_WIDTH(S_AXIS_FIFO_17_BYTE_WIDTH),
        .S_AXIS_FIFO_18_BYTE_WIDTH(S_AXIS_FIFO_18_BYTE_WIDTH),
        .S_AXIS_FIFO_19_BYTE_WIDTH(S_AXIS_FIFO_19_BYTE_WIDTH),
        .S_AXIS_FIFO_20_BYTE_WIDTH(S_AXIS_FIFO_20_BYTE_WIDTH),
        .S_AXIS_FIFO_21_BYTE_WIDTH(S_AXIS_FIFO_21_BYTE_WIDTH),
        .S_AXIS_FIFO_22_BYTE_WIDTH(S_AXIS_FIFO_22_BYTE_WIDTH),
        .S_AXIS_FIFO_23_BYTE_WIDTH(S_AXIS_FIFO_23_BYTE_WIDTH),
        .S_AXIS_FIFO_24_BYTE_WIDTH(S_AXIS_FIFO_24_BYTE_WIDTH),
        .S_AXIS_FIFO_25_BYTE_WIDTH(S_AXIS_FIFO_25_BYTE_WIDTH),
        .S_AXIS_FIFO_26_BYTE_WIDTH(S_AXIS_FIFO_26_BYTE_WIDTH),
        .S_AXIS_FIFO_27_BYTE_WIDTH(S_AXIS_FIFO_27_BYTE_WIDTH),
        .S_AXIS_FIFO_28_BYTE_WIDTH(S_AXIS_FIFO_28_BYTE_WIDTH),
        .S_AXIS_FIFO_29_BYTE_WIDTH(S_AXIS_FIFO_29_BYTE_WIDTH),
        .S_AXIS_FIFO_30_BYTE_WIDTH(S_AXIS_FIFO_30_BYTE_WIDTH),
        .S_AXIS_FIFO_31_BYTE_WIDTH(S_AXIS_FIFO_31_BYTE_WIDTH),
        .S_AXIS_FIFO_32_BYTE_WIDTH(S_AXIS_FIFO_32_BYTE_WIDTH),
        .S_AXIS_FIFO_33_BYTE_WIDTH(S_AXIS_FIFO_33_BYTE_WIDTH),
        .S_AXIS_FIFO_34_BYTE_WIDTH(S_AXIS_FIFO_34_BYTE_WIDTH),
        .S_AXIS_FIFO_35_BYTE_WIDTH(S_AXIS_FIFO_35_BYTE_WIDTH),
        .S_AXIS_FIFO_36_BYTE_WIDTH(S_AXIS_FIFO_36_BYTE_WIDTH),
        .S_AXIS_FIFO_37_BYTE_WIDTH(S_AXIS_FIFO_37_BYTE_WIDTH),
        .S_AXIS_FIFO_38_BYTE_WIDTH(S_AXIS_FIFO_38_BYTE_WIDTH),
        .S_AXIS_FIFO_39_BYTE_WIDTH(S_AXIS_FIFO_39_BYTE_WIDTH),
        .S_AXIS_FIFO_40_BYTE_WIDTH(S_AXIS_FIFO_40_BYTE_WIDTH),
        .S_AXIS_FIFO_41_BYTE_WIDTH(S_AXIS_FIFO_41_BYTE_WIDTH),
        .S_AXIS_FIFO_42_BYTE_WIDTH(S_AXIS_FIFO_42_BYTE_WIDTH),
        .S_AXIS_FIFO_43_BYTE_WIDTH(S_AXIS_FIFO_43_BYTE_WIDTH),
        .S_AXIS_FIFO_44_BYTE_WIDTH(S_AXIS_FIFO_44_BYTE_WIDTH),
        .S_AXIS_FIFO_45_BYTE_WIDTH(S_AXIS_FIFO_45_BYTE_WIDTH),
        .S_AXIS_FIFO_46_BYTE_WIDTH(S_AXIS_FIFO_46_BYTE_WIDTH),
        .S_AXIS_FIFO_47_BYTE_WIDTH(S_AXIS_FIFO_47_BYTE_WIDTH),
        .S_AXIS_FIFO_48_BYTE_WIDTH(S_AXIS_FIFO_48_BYTE_WIDTH),
        .S_AXIS_FIFO_49_BYTE_WIDTH(S_AXIS_FIFO_49_BYTE_WIDTH),
        .S_AXIS_FIFO_50_BYTE_WIDTH(S_AXIS_FIFO_50_BYTE_WIDTH),
        .S_AXIS_FIFO_51_BYTE_WIDTH(S_AXIS_FIFO_51_BYTE_WIDTH),
        .S_AXIS_FIFO_52_BYTE_WIDTH(S_AXIS_FIFO_52_BYTE_WIDTH),
        .S_AXIS_FIFO_53_BYTE_WIDTH(S_AXIS_FIFO_53_BYTE_WIDTH),
        .S_AXIS_FIFO_54_BYTE_WIDTH(S_AXIS_FIFO_54_BYTE_WIDTH),
        .S_AXIS_FIFO_55_BYTE_WIDTH(S_AXIS_FIFO_55_BYTE_WIDTH),
        .S_AXIS_FIFO_56_BYTE_WIDTH(S_AXIS_FIFO_56_BYTE_WIDTH),
        .S_AXIS_FIFO_57_BYTE_WIDTH(S_AXIS_FIFO_57_BYTE_WIDTH),
        .S_AXIS_FIFO_58_BYTE_WIDTH(S_AXIS_FIFO_58_BYTE_WIDTH),
        .S_AXIS_FIFO_59_BYTE_WIDTH(S_AXIS_FIFO_59_BYTE_WIDTH),
        .S_AXIS_FIFO_60_BYTE_WIDTH(S_AXIS_FIFO_60_BYTE_WIDTH),
        .S_AXIS_FIFO_61_BYTE_WIDTH(S_AXIS_FIFO_61_BYTE_WIDTH),
        .S_AXIS_FIFO_62_BYTE_WIDTH(S_AXIS_FIFO_62_BYTE_WIDTH),
        .S_AXIS_FIFO_63_BYTE_WIDTH(S_AXIS_FIFO_63_BYTE_WIDTH),
        .S_AXIS_FIFO_64_BYTE_WIDTH(S_AXIS_FIFO_64_BYTE_WIDTH),
        .S_AXIS_FIFO_65_BYTE_WIDTH(S_AXIS_FIFO_65_BYTE_WIDTH),
        .S_AXIS_FIFO_66_BYTE_WIDTH(S_AXIS_FIFO_66_BYTE_WIDTH),
        .S_AXIS_FIFO_67_BYTE_WIDTH(S_AXIS_FIFO_67_BYTE_WIDTH),
        .S_AXIS_FIFO_68_BYTE_WIDTH(S_AXIS_FIFO_68_BYTE_WIDTH),
        .S_AXIS_FIFO_69_BYTE_WIDTH(S_AXIS_FIFO_69_BYTE_WIDTH),
        .S_AXIS_FIFO_70_BYTE_WIDTH(S_AXIS_FIFO_70_BYTE_WIDTH),
        .S_AXIS_FIFO_71_BYTE_WIDTH(S_AXIS_FIFO_71_BYTE_WIDTH),
        .S_AXIS_FIFO_72_BYTE_WIDTH(S_AXIS_FIFO_72_BYTE_WIDTH),
        .S_AXIS_FIFO_73_BYTE_WIDTH(S_AXIS_FIFO_73_BYTE_WIDTH),
        .S_AXIS_FIFO_74_BYTE_WIDTH(S_AXIS_FIFO_74_BYTE_WIDTH),
        .S_AXIS_FIFO_75_BYTE_WIDTH(S_AXIS_FIFO_75_BYTE_WIDTH),
        .S_AXIS_FIFO_76_BYTE_WIDTH(S_AXIS_FIFO_76_BYTE_WIDTH),
        .S_AXIS_FIFO_77_BYTE_WIDTH(S_AXIS_FIFO_77_BYTE_WIDTH),
        .S_AXIS_FIFO_78_BYTE_WIDTH(S_AXIS_FIFO_78_BYTE_WIDTH),
        .S_AXIS_FIFO_79_BYTE_WIDTH(S_AXIS_FIFO_79_BYTE_WIDTH),
        .S_AXIS_FIFO_80_BYTE_WIDTH(S_AXIS_FIFO_80_BYTE_WIDTH),
        .S_AXIS_FIFO_81_BYTE_WIDTH(S_AXIS_FIFO_81_BYTE_WIDTH),
        .S_AXIS_FIFO_82_BYTE_WIDTH(S_AXIS_FIFO_82_BYTE_WIDTH),
        .S_AXIS_FIFO_83_BYTE_WIDTH(S_AXIS_FIFO_83_BYTE_WIDTH),
        .S_AXIS_FIFO_84_BYTE_WIDTH(S_AXIS_FIFO_84_BYTE_WIDTH),
        .S_AXIS_FIFO_85_BYTE_WIDTH(S_AXIS_FIFO_85_BYTE_WIDTH),
        .S_AXIS_FIFO_86_BYTE_WIDTH(S_AXIS_FIFO_86_BYTE_WIDTH),
        .S_AXIS_FIFO_87_BYTE_WIDTH(S_AXIS_FIFO_87_BYTE_WIDTH),
        .S_AXIS_FIFO_88_BYTE_WIDTH(S_AXIS_FIFO_88_BYTE_WIDTH),
        .S_AXIS_FIFO_89_BYTE_WIDTH(S_AXIS_FIFO_89_BYTE_WIDTH),
        .S_AXIS_FIFO_90_BYTE_WIDTH(S_AXIS_FIFO_90_BYTE_WIDTH),
        .S_AXIS_FIFO_91_BYTE_WIDTH(S_AXIS_FIFO_91_BYTE_WIDTH),
        .S_AXIS_FIFO_92_BYTE_WIDTH(S_AXIS_FIFO_92_BYTE_WIDTH),
        .S_AXIS_FIFO_93_BYTE_WIDTH(S_AXIS_FIFO_93_BYTE_WIDTH),
        .S_AXIS_FIFO_94_BYTE_WIDTH(S_AXIS_FIFO_94_BYTE_WIDTH),
        .S_AXIS_FIFO_95_BYTE_WIDTH(S_AXIS_FIFO_95_BYTE_WIDTH),
        .S_AXIS_FIFO_96_BYTE_WIDTH(S_AXIS_FIFO_96_BYTE_WIDTH),
        .S_AXIS_FIFO_97_BYTE_WIDTH(S_AXIS_FIFO_97_BYTE_WIDTH),
        .S_AXIS_FIFO_98_BYTE_WIDTH(S_AXIS_FIFO_98_BYTE_WIDTH),
        .S_AXIS_FIFO_99_BYTE_WIDTH(S_AXIS_FIFO_99_BYTE_WIDTH),
        .S_AXIS_FIFO_100_BYTE_WIDTH(S_AXIS_FIFO_100_BYTE_WIDTH),
        .S_AXIS_FIFO_101_BYTE_WIDTH(S_AXIS_FIFO_101_BYTE_WIDTH),
        .S_AXIS_FIFO_102_BYTE_WIDTH(S_AXIS_FIFO_102_BYTE_WIDTH),
        .S_AXIS_FIFO_103_BYTE_WIDTH(S_AXIS_FIFO_103_BYTE_WIDTH),
        .S_AXIS_FIFO_104_BYTE_WIDTH(S_AXIS_FIFO_104_BYTE_WIDTH),
        .S_AXIS_FIFO_105_BYTE_WIDTH(S_AXIS_FIFO_105_BYTE_WIDTH),
        .S_AXIS_FIFO_106_BYTE_WIDTH(S_AXIS_FIFO_106_BYTE_WIDTH),
        .S_AXIS_FIFO_107_BYTE_WIDTH(S_AXIS_FIFO_107_BYTE_WIDTH),
        .S_AXIS_FIFO_108_BYTE_WIDTH(S_AXIS_FIFO_108_BYTE_WIDTH),
        .S_AXIS_FIFO_109_BYTE_WIDTH(S_AXIS_FIFO_109_BYTE_WIDTH),
        .S_AXIS_FIFO_110_BYTE_WIDTH(S_AXIS_FIFO_110_BYTE_WIDTH),
        .S_AXIS_FIFO_111_BYTE_WIDTH(S_AXIS_FIFO_111_BYTE_WIDTH),
        .S_AXIS_FIFO_112_BYTE_WIDTH(S_AXIS_FIFO_112_BYTE_WIDTH),
        .S_AXIS_FIFO_113_BYTE_WIDTH(S_AXIS_FIFO_113_BYTE_WIDTH),
        .S_AXIS_FIFO_114_BYTE_WIDTH(S_AXIS_FIFO_114_BYTE_WIDTH),
        .S_AXIS_FIFO_115_BYTE_WIDTH(S_AXIS_FIFO_115_BYTE_WIDTH),
        .S_AXIS_FIFO_116_BYTE_WIDTH(S_AXIS_FIFO_116_BYTE_WIDTH),
        .S_AXIS_FIFO_117_BYTE_WIDTH(S_AXIS_FIFO_117_BYTE_WIDTH),
        .S_AXIS_FIFO_118_BYTE_WIDTH(S_AXIS_FIFO_118_BYTE_WIDTH),
        .S_AXIS_FIFO_119_BYTE_WIDTH(S_AXIS_FIFO_119_BYTE_WIDTH),
        .S_AXIS_FIFO_120_BYTE_WIDTH(S_AXIS_FIFO_120_BYTE_WIDTH),
        .S_AXIS_FIFO_121_BYTE_WIDTH(S_AXIS_FIFO_121_BYTE_WIDTH),
        .S_AXIS_FIFO_122_BYTE_WIDTH(S_AXIS_FIFO_122_BYTE_WIDTH),
        .S_AXIS_FIFO_123_BYTE_WIDTH(S_AXIS_FIFO_123_BYTE_WIDTH),
        .S_AXIS_FIFO_124_BYTE_WIDTH(S_AXIS_FIFO_124_BYTE_WIDTH),
        .S_AXIS_FIFO_125_BYTE_WIDTH(S_AXIS_FIFO_125_BYTE_WIDTH),
        .S_AXIS_FIFO_126_BYTE_WIDTH(S_AXIS_FIFO_126_BYTE_WIDTH),
        .S_AXIS_FIFO_127_BYTE_WIDTH(S_AXIS_FIFO_127_BYTE_WIDTH),
        .S_AXIS_FIFO_0_DMWIDTH(S_AXIS_FIFO_0_DMWIDTH),
        .S_AXIS_FIFO_1_DMWIDTH(S_AXIS_FIFO_1_DMWIDTH),
        .S_AXIS_FIFO_2_DMWIDTH(S_AXIS_FIFO_2_DMWIDTH),
        .S_AXIS_FIFO_3_DMWIDTH(S_AXIS_FIFO_3_DMWIDTH),
        .S_AXIS_FIFO_4_DMWIDTH(S_AXIS_FIFO_4_DMWIDTH),
        .S_AXIS_FIFO_5_DMWIDTH(S_AXIS_FIFO_5_DMWIDTH),
        .S_AXIS_FIFO_6_DMWIDTH(S_AXIS_FIFO_6_DMWIDTH),
        .S_AXIS_FIFO_7_DMWIDTH(S_AXIS_FIFO_7_DMWIDTH),
        .S_AXIS_FIFO_8_DMWIDTH(S_AXIS_FIFO_8_DMWIDTH),
        .S_AXIS_FIFO_9_DMWIDTH(S_AXIS_FIFO_9_DMWIDTH),
        .S_AXIS_FIFO_10_DMWIDTH(S_AXIS_FIFO_10_DMWIDTH),
        .S_AXIS_FIFO_11_DMWIDTH(S_AXIS_FIFO_11_DMWIDTH),
        .S_AXIS_FIFO_12_DMWIDTH(S_AXIS_FIFO_12_DMWIDTH),
        .S_AXIS_FIFO_13_DMWIDTH(S_AXIS_FIFO_13_DMWIDTH),
        .S_AXIS_FIFO_14_DMWIDTH(S_AXIS_FIFO_14_DMWIDTH),
        .S_AXIS_FIFO_15_DMWIDTH(S_AXIS_FIFO_15_DMWIDTH),
        .S_AXIS_FIFO_16_DMWIDTH(S_AXIS_FIFO_16_DMWIDTH),
        .S_AXIS_FIFO_17_DMWIDTH(S_AXIS_FIFO_17_DMWIDTH),
        .S_AXIS_FIFO_18_DMWIDTH(S_AXIS_FIFO_18_DMWIDTH),
        .S_AXIS_FIFO_19_DMWIDTH(S_AXIS_FIFO_19_DMWIDTH),
        .S_AXIS_FIFO_20_DMWIDTH(S_AXIS_FIFO_20_DMWIDTH),
        .S_AXIS_FIFO_21_DMWIDTH(S_AXIS_FIFO_21_DMWIDTH),
        .S_AXIS_FIFO_22_DMWIDTH(S_AXIS_FIFO_22_DMWIDTH),
        .S_AXIS_FIFO_23_DMWIDTH(S_AXIS_FIFO_23_DMWIDTH),
        .S_AXIS_FIFO_24_DMWIDTH(S_AXIS_FIFO_24_DMWIDTH),
        .S_AXIS_FIFO_25_DMWIDTH(S_AXIS_FIFO_25_DMWIDTH),
        .S_AXIS_FIFO_26_DMWIDTH(S_AXIS_FIFO_26_DMWIDTH),
        .S_AXIS_FIFO_27_DMWIDTH(S_AXIS_FIFO_27_DMWIDTH),
        .S_AXIS_FIFO_28_DMWIDTH(S_AXIS_FIFO_28_DMWIDTH),
        .S_AXIS_FIFO_29_DMWIDTH(S_AXIS_FIFO_29_DMWIDTH),
        .S_AXIS_FIFO_30_DMWIDTH(S_AXIS_FIFO_30_DMWIDTH),
        .S_AXIS_FIFO_31_DMWIDTH(S_AXIS_FIFO_31_DMWIDTH),
        .S_AXIS_FIFO_32_DMWIDTH(S_AXIS_FIFO_32_DMWIDTH),
        .S_AXIS_FIFO_33_DMWIDTH(S_AXIS_FIFO_33_DMWIDTH),
        .S_AXIS_FIFO_34_DMWIDTH(S_AXIS_FIFO_34_DMWIDTH),
        .S_AXIS_FIFO_35_DMWIDTH(S_AXIS_FIFO_35_DMWIDTH),
        .S_AXIS_FIFO_36_DMWIDTH(S_AXIS_FIFO_36_DMWIDTH),
        .S_AXIS_FIFO_37_DMWIDTH(S_AXIS_FIFO_37_DMWIDTH),
        .S_AXIS_FIFO_38_DMWIDTH(S_AXIS_FIFO_38_DMWIDTH),
        .S_AXIS_FIFO_39_DMWIDTH(S_AXIS_FIFO_39_DMWIDTH),
        .S_AXIS_FIFO_40_DMWIDTH(S_AXIS_FIFO_40_DMWIDTH),
        .S_AXIS_FIFO_41_DMWIDTH(S_AXIS_FIFO_41_DMWIDTH),
        .S_AXIS_FIFO_42_DMWIDTH(S_AXIS_FIFO_42_DMWIDTH),
        .S_AXIS_FIFO_43_DMWIDTH(S_AXIS_FIFO_43_DMWIDTH),
        .S_AXIS_FIFO_44_DMWIDTH(S_AXIS_FIFO_44_DMWIDTH),
        .S_AXIS_FIFO_45_DMWIDTH(S_AXIS_FIFO_45_DMWIDTH),
        .S_AXIS_FIFO_46_DMWIDTH(S_AXIS_FIFO_46_DMWIDTH),
        .S_AXIS_FIFO_47_DMWIDTH(S_AXIS_FIFO_47_DMWIDTH),
        .S_AXIS_FIFO_48_DMWIDTH(S_AXIS_FIFO_48_DMWIDTH),
        .S_AXIS_FIFO_49_DMWIDTH(S_AXIS_FIFO_49_DMWIDTH),
        .S_AXIS_FIFO_50_DMWIDTH(S_AXIS_FIFO_50_DMWIDTH),
        .S_AXIS_FIFO_51_DMWIDTH(S_AXIS_FIFO_51_DMWIDTH),
        .S_AXIS_FIFO_52_DMWIDTH(S_AXIS_FIFO_52_DMWIDTH),
        .S_AXIS_FIFO_53_DMWIDTH(S_AXIS_FIFO_53_DMWIDTH),
        .S_AXIS_FIFO_54_DMWIDTH(S_AXIS_FIFO_54_DMWIDTH),
        .S_AXIS_FIFO_55_DMWIDTH(S_AXIS_FIFO_55_DMWIDTH),
        .S_AXIS_FIFO_56_DMWIDTH(S_AXIS_FIFO_56_DMWIDTH),
        .S_AXIS_FIFO_57_DMWIDTH(S_AXIS_FIFO_57_DMWIDTH),
        .S_AXIS_FIFO_58_DMWIDTH(S_AXIS_FIFO_58_DMWIDTH),
        .S_AXIS_FIFO_59_DMWIDTH(S_AXIS_FIFO_59_DMWIDTH),
        .S_AXIS_FIFO_60_DMWIDTH(S_AXIS_FIFO_60_DMWIDTH),
        .S_AXIS_FIFO_61_DMWIDTH(S_AXIS_FIFO_61_DMWIDTH),
        .S_AXIS_FIFO_62_DMWIDTH(S_AXIS_FIFO_62_DMWIDTH),
        .S_AXIS_FIFO_63_DMWIDTH(S_AXIS_FIFO_63_DMWIDTH),
        .S_AXIS_FIFO_64_DMWIDTH(S_AXIS_FIFO_64_DMWIDTH),
        .S_AXIS_FIFO_65_DMWIDTH(S_AXIS_FIFO_65_DMWIDTH),
        .S_AXIS_FIFO_66_DMWIDTH(S_AXIS_FIFO_66_DMWIDTH),
        .S_AXIS_FIFO_67_DMWIDTH(S_AXIS_FIFO_67_DMWIDTH),
        .S_AXIS_FIFO_68_DMWIDTH(S_AXIS_FIFO_68_DMWIDTH),
        .S_AXIS_FIFO_69_DMWIDTH(S_AXIS_FIFO_69_DMWIDTH),
        .S_AXIS_FIFO_70_DMWIDTH(S_AXIS_FIFO_70_DMWIDTH),
        .S_AXIS_FIFO_71_DMWIDTH(S_AXIS_FIFO_71_DMWIDTH),
        .S_AXIS_FIFO_72_DMWIDTH(S_AXIS_FIFO_72_DMWIDTH),
        .S_AXIS_FIFO_73_DMWIDTH(S_AXIS_FIFO_73_DMWIDTH),
        .S_AXIS_FIFO_74_DMWIDTH(S_AXIS_FIFO_74_DMWIDTH),
        .S_AXIS_FIFO_75_DMWIDTH(S_AXIS_FIFO_75_DMWIDTH),
        .S_AXIS_FIFO_76_DMWIDTH(S_AXIS_FIFO_76_DMWIDTH),
        .S_AXIS_FIFO_77_DMWIDTH(S_AXIS_FIFO_77_DMWIDTH),
        .S_AXIS_FIFO_78_DMWIDTH(S_AXIS_FIFO_78_DMWIDTH),
        .S_AXIS_FIFO_79_DMWIDTH(S_AXIS_FIFO_79_DMWIDTH),
        .S_AXIS_FIFO_80_DMWIDTH(S_AXIS_FIFO_80_DMWIDTH),
        .S_AXIS_FIFO_81_DMWIDTH(S_AXIS_FIFO_81_DMWIDTH),
        .S_AXIS_FIFO_82_DMWIDTH(S_AXIS_FIFO_82_DMWIDTH),
        .S_AXIS_FIFO_83_DMWIDTH(S_AXIS_FIFO_83_DMWIDTH),
        .S_AXIS_FIFO_84_DMWIDTH(S_AXIS_FIFO_84_DMWIDTH),
        .S_AXIS_FIFO_85_DMWIDTH(S_AXIS_FIFO_85_DMWIDTH),
        .S_AXIS_FIFO_86_DMWIDTH(S_AXIS_FIFO_86_DMWIDTH),
        .S_AXIS_FIFO_87_DMWIDTH(S_AXIS_FIFO_87_DMWIDTH),
        .S_AXIS_FIFO_88_DMWIDTH(S_AXIS_FIFO_88_DMWIDTH),
        .S_AXIS_FIFO_89_DMWIDTH(S_AXIS_FIFO_89_DMWIDTH),
        .S_AXIS_FIFO_90_DMWIDTH(S_AXIS_FIFO_90_DMWIDTH),
        .S_AXIS_FIFO_91_DMWIDTH(S_AXIS_FIFO_91_DMWIDTH),
        .S_AXIS_FIFO_92_DMWIDTH(S_AXIS_FIFO_92_DMWIDTH),
        .S_AXIS_FIFO_93_DMWIDTH(S_AXIS_FIFO_93_DMWIDTH),
        .S_AXIS_FIFO_94_DMWIDTH(S_AXIS_FIFO_94_DMWIDTH),
        .S_AXIS_FIFO_95_DMWIDTH(S_AXIS_FIFO_95_DMWIDTH),
        .S_AXIS_FIFO_96_DMWIDTH(S_AXIS_FIFO_96_DMWIDTH),
        .S_AXIS_FIFO_97_DMWIDTH(S_AXIS_FIFO_97_DMWIDTH),
        .S_AXIS_FIFO_98_DMWIDTH(S_AXIS_FIFO_98_DMWIDTH),
        .S_AXIS_FIFO_99_DMWIDTH(S_AXIS_FIFO_99_DMWIDTH),
        .S_AXIS_FIFO_100_DMWIDTH(S_AXIS_FIFO_100_DMWIDTH),
        .S_AXIS_FIFO_101_DMWIDTH(S_AXIS_FIFO_101_DMWIDTH),
        .S_AXIS_FIFO_102_DMWIDTH(S_AXIS_FIFO_102_DMWIDTH),
        .S_AXIS_FIFO_103_DMWIDTH(S_AXIS_FIFO_103_DMWIDTH),
        .S_AXIS_FIFO_104_DMWIDTH(S_AXIS_FIFO_104_DMWIDTH),
        .S_AXIS_FIFO_105_DMWIDTH(S_AXIS_FIFO_105_DMWIDTH),
        .S_AXIS_FIFO_106_DMWIDTH(S_AXIS_FIFO_106_DMWIDTH),
        .S_AXIS_FIFO_107_DMWIDTH(S_AXIS_FIFO_107_DMWIDTH),
        .S_AXIS_FIFO_108_DMWIDTH(S_AXIS_FIFO_108_DMWIDTH),
        .S_AXIS_FIFO_109_DMWIDTH(S_AXIS_FIFO_109_DMWIDTH),
        .S_AXIS_FIFO_110_DMWIDTH(S_AXIS_FIFO_110_DMWIDTH),
        .S_AXIS_FIFO_111_DMWIDTH(S_AXIS_FIFO_111_DMWIDTH),
        .S_AXIS_FIFO_112_DMWIDTH(S_AXIS_FIFO_112_DMWIDTH),
        .S_AXIS_FIFO_113_DMWIDTH(S_AXIS_FIFO_113_DMWIDTH),
        .S_AXIS_FIFO_114_DMWIDTH(S_AXIS_FIFO_114_DMWIDTH),
        .S_AXIS_FIFO_115_DMWIDTH(S_AXIS_FIFO_115_DMWIDTH),
        .S_AXIS_FIFO_116_DMWIDTH(S_AXIS_FIFO_116_DMWIDTH),
        .S_AXIS_FIFO_117_DMWIDTH(S_AXIS_FIFO_117_DMWIDTH),
        .S_AXIS_FIFO_118_DMWIDTH(S_AXIS_FIFO_118_DMWIDTH),
        .S_AXIS_FIFO_119_DMWIDTH(S_AXIS_FIFO_119_DMWIDTH),
        .S_AXIS_FIFO_120_DMWIDTH(S_AXIS_FIFO_120_DMWIDTH),
        .S_AXIS_FIFO_121_DMWIDTH(S_AXIS_FIFO_121_DMWIDTH),
        .S_AXIS_FIFO_122_DMWIDTH(S_AXIS_FIFO_122_DMWIDTH),
        .S_AXIS_FIFO_123_DMWIDTH(S_AXIS_FIFO_123_DMWIDTH),
        .S_AXIS_FIFO_124_DMWIDTH(S_AXIS_FIFO_124_DMWIDTH),
        .S_AXIS_FIFO_125_DMWIDTH(S_AXIS_FIFO_125_DMWIDTH),
        .S_AXIS_FIFO_126_DMWIDTH(S_AXIS_FIFO_126_DMWIDTH),
        .S_AXIS_FIFO_127_DMWIDTH(S_AXIS_FIFO_127_DMWIDTH)
    ) in_fifo_args_i (
        .acc_clk(acc_aclk),
        .acc_aresetn(acc_aresetn),
        .in_fifo_allow(infifo_ctrl_allow),
        .s_axis_fifo_0_aclk(s_axis_fifo_0_aclk),
        .s_axis_fifo_0_aresetn(s_axis_fifo_0_aresetn),
        .s_axis_fifo_0_tlast(s_axis_fifo_0_tlast),
        .s_axis_fifo_0_tvalid(s_axis_fifo_0_tvalid),
        .s_axis_fifo_0_tkeep(s_axis_fifo_0_tkeep),
        .s_axis_fifo_0_tstrb(s_axis_fifo_0_tstrb),
        .s_axis_fifo_0_tdata(s_axis_fifo_0_tdata),
        .s_axis_fifo_0_tready(s_axis_fifo_0_tready),
        .ap_fifo_iarg_0_empty_n(ap_fifo_iarg_0_empty_n),
        .ap_fifo_iarg_0_dout(ap_fifo_iarg_0_dout),
        .ap_fifo_iarg_0_read(ap_fifo_iarg_0_read),
        .s_axis_fifo_1_aclk(s_axis_fifo_1_aclk),
        .s_axis_fifo_1_aresetn(s_axis_fifo_1_aresetn),
        .s_axis_fifo_1_tlast(s_axis_fifo_1_tlast),
        .s_axis_fifo_1_tvalid(s_axis_fifo_1_tvalid),
        .s_axis_fifo_1_tkeep(s_axis_fifo_1_tkeep),
        .s_axis_fifo_1_tstrb(s_axis_fifo_1_tstrb),
        .s_axis_fifo_1_tdata(s_axis_fifo_1_tdata),
        .s_axis_fifo_1_tready(s_axis_fifo_1_tready),
        .ap_fifo_iarg_1_empty_n(ap_fifo_iarg_1_empty_n),
        .ap_fifo_iarg_1_dout(ap_fifo_iarg_1_dout),
        .ap_fifo_iarg_1_read(ap_fifo_iarg_1_read),
        .s_axis_fifo_2_aclk(s_axis_fifo_2_aclk),
        .s_axis_fifo_2_aresetn(s_axis_fifo_2_aresetn),
        .s_axis_fifo_2_tlast(s_axis_fifo_2_tlast),
        .s_axis_fifo_2_tvalid(s_axis_fifo_2_tvalid),
        .s_axis_fifo_2_tkeep(s_axis_fifo_2_tkeep),
        .s_axis_fifo_2_tstrb(s_axis_fifo_2_tstrb),
        .s_axis_fifo_2_tdata(s_axis_fifo_2_tdata),
        .s_axis_fifo_2_tready(s_axis_fifo_2_tready),
        .ap_fifo_iarg_2_empty_n(ap_fifo_iarg_2_empty_n),
        .ap_fifo_iarg_2_dout(ap_fifo_iarg_2_dout),
        .ap_fifo_iarg_2_read(ap_fifo_iarg_2_read),
        .s_axis_fifo_3_aclk(s_axis_fifo_3_aclk),
        .s_axis_fifo_3_aresetn(s_axis_fifo_3_aresetn),
        .s_axis_fifo_3_tlast(s_axis_fifo_3_tlast),
        .s_axis_fifo_3_tvalid(s_axis_fifo_3_tvalid),
        .s_axis_fifo_3_tkeep(s_axis_fifo_3_tkeep),
        .s_axis_fifo_3_tstrb(s_axis_fifo_3_tstrb),
        .s_axis_fifo_3_tdata(s_axis_fifo_3_tdata),
        .s_axis_fifo_3_tready(s_axis_fifo_3_tready),
        .ap_fifo_iarg_3_empty_n(ap_fifo_iarg_3_empty_n),
        .ap_fifo_iarg_3_dout(ap_fifo_iarg_3_dout),
        .ap_fifo_iarg_3_read(ap_fifo_iarg_3_read),
        .s_axis_fifo_4_aclk(s_axis_fifo_4_aclk),
        .s_axis_fifo_4_aresetn(s_axis_fifo_4_aresetn),
        .s_axis_fifo_4_tlast(s_axis_fifo_4_tlast),
        .s_axis_fifo_4_tvalid(s_axis_fifo_4_tvalid),
        .s_axis_fifo_4_tkeep(s_axis_fifo_4_tkeep),
        .s_axis_fifo_4_tstrb(s_axis_fifo_4_tstrb),
        .s_axis_fifo_4_tdata(s_axis_fifo_4_tdata),
        .s_axis_fifo_4_tready(s_axis_fifo_4_tready),
        .ap_fifo_iarg_4_empty_n(ap_fifo_iarg_4_empty_n),
        .ap_fifo_iarg_4_dout(ap_fifo_iarg_4_dout),
        .ap_fifo_iarg_4_read(ap_fifo_iarg_4_read),
        .s_axis_fifo_5_aclk(s_axis_fifo_5_aclk),
        .s_axis_fifo_5_aresetn(s_axis_fifo_5_aresetn),
        .s_axis_fifo_5_tlast(s_axis_fifo_5_tlast),
        .s_axis_fifo_5_tvalid(s_axis_fifo_5_tvalid),
        .s_axis_fifo_5_tkeep(s_axis_fifo_5_tkeep),
        .s_axis_fifo_5_tstrb(s_axis_fifo_5_tstrb),
        .s_axis_fifo_5_tdata(s_axis_fifo_5_tdata),
        .s_axis_fifo_5_tready(s_axis_fifo_5_tready),
        .ap_fifo_iarg_5_empty_n(ap_fifo_iarg_5_empty_n),
        .ap_fifo_iarg_5_dout(ap_fifo_iarg_5_dout),
        .ap_fifo_iarg_5_read(ap_fifo_iarg_5_read),
        .s_axis_fifo_6_aclk(s_axis_fifo_6_aclk),
        .s_axis_fifo_6_aresetn(s_axis_fifo_6_aresetn),
        .s_axis_fifo_6_tlast(s_axis_fifo_6_tlast),
        .s_axis_fifo_6_tvalid(s_axis_fifo_6_tvalid),
        .s_axis_fifo_6_tkeep(s_axis_fifo_6_tkeep),
        .s_axis_fifo_6_tstrb(s_axis_fifo_6_tstrb),
        .s_axis_fifo_6_tdata(s_axis_fifo_6_tdata),
        .s_axis_fifo_6_tready(s_axis_fifo_6_tready),
        .ap_fifo_iarg_6_empty_n(ap_fifo_iarg_6_empty_n),
        .ap_fifo_iarg_6_dout(ap_fifo_iarg_6_dout),
        .ap_fifo_iarg_6_read(ap_fifo_iarg_6_read),
        .s_axis_fifo_7_aclk(s_axis_fifo_7_aclk),
        .s_axis_fifo_7_aresetn(s_axis_fifo_7_aresetn),
        .s_axis_fifo_7_tlast(s_axis_fifo_7_tlast),
        .s_axis_fifo_7_tvalid(s_axis_fifo_7_tvalid),
        .s_axis_fifo_7_tkeep(s_axis_fifo_7_tkeep),
        .s_axis_fifo_7_tstrb(s_axis_fifo_7_tstrb),
        .s_axis_fifo_7_tdata(s_axis_fifo_7_tdata),
        .s_axis_fifo_7_tready(s_axis_fifo_7_tready),
        .ap_fifo_iarg_7_empty_n(ap_fifo_iarg_7_empty_n),
        .ap_fifo_iarg_7_dout(ap_fifo_iarg_7_dout),
        .ap_fifo_iarg_7_read(ap_fifo_iarg_7_read),
        .s_axis_fifo_8_aclk(s_axis_fifo_8_aclk),
        .s_axis_fifo_8_aresetn(s_axis_fifo_8_aresetn),
        .s_axis_fifo_8_tlast(s_axis_fifo_8_tlast),
        .s_axis_fifo_8_tvalid(s_axis_fifo_8_tvalid),
        .s_axis_fifo_8_tkeep(s_axis_fifo_8_tkeep),
        .s_axis_fifo_8_tstrb(s_axis_fifo_8_tstrb),
        .s_axis_fifo_8_tdata(s_axis_fifo_8_tdata),
        .s_axis_fifo_8_tready(s_axis_fifo_8_tready),
        .ap_fifo_iarg_8_empty_n(ap_fifo_iarg_8_empty_n),
        .ap_fifo_iarg_8_dout(ap_fifo_iarg_8_dout),
        .ap_fifo_iarg_8_read(ap_fifo_iarg_8_read),
        .s_axis_fifo_9_aclk(s_axis_fifo_9_aclk),
        .s_axis_fifo_9_aresetn(s_axis_fifo_9_aresetn),
        .s_axis_fifo_9_tlast(s_axis_fifo_9_tlast),
        .s_axis_fifo_9_tvalid(s_axis_fifo_9_tvalid),
        .s_axis_fifo_9_tkeep(s_axis_fifo_9_tkeep),
        .s_axis_fifo_9_tstrb(s_axis_fifo_9_tstrb),
        .s_axis_fifo_9_tdata(s_axis_fifo_9_tdata),
        .s_axis_fifo_9_tready(s_axis_fifo_9_tready),
        .ap_fifo_iarg_9_empty_n(ap_fifo_iarg_9_empty_n),
        .ap_fifo_iarg_9_dout(ap_fifo_iarg_9_dout),
        .ap_fifo_iarg_9_read(ap_fifo_iarg_9_read),
        .s_axis_fifo_10_aclk(s_axis_fifo_10_aclk),
        .s_axis_fifo_10_aresetn(s_axis_fifo_10_aresetn),
        .s_axis_fifo_10_tlast(s_axis_fifo_10_tlast),
        .s_axis_fifo_10_tvalid(s_axis_fifo_10_tvalid),
        .s_axis_fifo_10_tkeep(s_axis_fifo_10_tkeep),
        .s_axis_fifo_10_tstrb(s_axis_fifo_10_tstrb),
        .s_axis_fifo_10_tdata(s_axis_fifo_10_tdata),
        .s_axis_fifo_10_tready(s_axis_fifo_10_tready),
        .ap_fifo_iarg_10_empty_n(ap_fifo_iarg_10_empty_n),
        .ap_fifo_iarg_10_dout(ap_fifo_iarg_10_dout),
        .ap_fifo_iarg_10_read(ap_fifo_iarg_10_read),
        .s_axis_fifo_11_aclk(s_axis_fifo_11_aclk),
        .s_axis_fifo_11_aresetn(s_axis_fifo_11_aresetn),
        .s_axis_fifo_11_tlast(s_axis_fifo_11_tlast),
        .s_axis_fifo_11_tvalid(s_axis_fifo_11_tvalid),
        .s_axis_fifo_11_tkeep(s_axis_fifo_11_tkeep),
        .s_axis_fifo_11_tstrb(s_axis_fifo_11_tstrb),
        .s_axis_fifo_11_tdata(s_axis_fifo_11_tdata),
        .s_axis_fifo_11_tready(s_axis_fifo_11_tready),
        .ap_fifo_iarg_11_empty_n(ap_fifo_iarg_11_empty_n),
        .ap_fifo_iarg_11_dout(ap_fifo_iarg_11_dout),
        .ap_fifo_iarg_11_read(ap_fifo_iarg_11_read),
        .s_axis_fifo_12_aclk(s_axis_fifo_12_aclk),
        .s_axis_fifo_12_aresetn(s_axis_fifo_12_aresetn),
        .s_axis_fifo_12_tlast(s_axis_fifo_12_tlast),
        .s_axis_fifo_12_tvalid(s_axis_fifo_12_tvalid),
        .s_axis_fifo_12_tkeep(s_axis_fifo_12_tkeep),
        .s_axis_fifo_12_tstrb(s_axis_fifo_12_tstrb),
        .s_axis_fifo_12_tdata(s_axis_fifo_12_tdata),
        .s_axis_fifo_12_tready(s_axis_fifo_12_tready),
        .ap_fifo_iarg_12_empty_n(ap_fifo_iarg_12_empty_n),
        .ap_fifo_iarg_12_dout(ap_fifo_iarg_12_dout),
        .ap_fifo_iarg_12_read(ap_fifo_iarg_12_read),
        .s_axis_fifo_13_aclk(s_axis_fifo_13_aclk),
        .s_axis_fifo_13_aresetn(s_axis_fifo_13_aresetn),
        .s_axis_fifo_13_tlast(s_axis_fifo_13_tlast),
        .s_axis_fifo_13_tvalid(s_axis_fifo_13_tvalid),
        .s_axis_fifo_13_tkeep(s_axis_fifo_13_tkeep),
        .s_axis_fifo_13_tstrb(s_axis_fifo_13_tstrb),
        .s_axis_fifo_13_tdata(s_axis_fifo_13_tdata),
        .s_axis_fifo_13_tready(s_axis_fifo_13_tready),
        .ap_fifo_iarg_13_empty_n(ap_fifo_iarg_13_empty_n),
        .ap_fifo_iarg_13_dout(ap_fifo_iarg_13_dout),
        .ap_fifo_iarg_13_read(ap_fifo_iarg_13_read),
        .s_axis_fifo_14_aclk(s_axis_fifo_14_aclk),
        .s_axis_fifo_14_aresetn(s_axis_fifo_14_aresetn),
        .s_axis_fifo_14_tlast(s_axis_fifo_14_tlast),
        .s_axis_fifo_14_tvalid(s_axis_fifo_14_tvalid),
        .s_axis_fifo_14_tkeep(s_axis_fifo_14_tkeep),
        .s_axis_fifo_14_tstrb(s_axis_fifo_14_tstrb),
        .s_axis_fifo_14_tdata(s_axis_fifo_14_tdata),
        .s_axis_fifo_14_tready(s_axis_fifo_14_tready),
        .ap_fifo_iarg_14_empty_n(ap_fifo_iarg_14_empty_n),
        .ap_fifo_iarg_14_dout(ap_fifo_iarg_14_dout),
        .ap_fifo_iarg_14_read(ap_fifo_iarg_14_read),
        .s_axis_fifo_15_aclk(s_axis_fifo_15_aclk),
        .s_axis_fifo_15_aresetn(s_axis_fifo_15_aresetn),
        .s_axis_fifo_15_tlast(s_axis_fifo_15_tlast),
        .s_axis_fifo_15_tvalid(s_axis_fifo_15_tvalid),
        .s_axis_fifo_15_tkeep(s_axis_fifo_15_tkeep),
        .s_axis_fifo_15_tstrb(s_axis_fifo_15_tstrb),
        .s_axis_fifo_15_tdata(s_axis_fifo_15_tdata),
        .s_axis_fifo_15_tready(s_axis_fifo_15_tready),
        .ap_fifo_iarg_15_empty_n(ap_fifo_iarg_15_empty_n),
        .ap_fifo_iarg_15_dout(ap_fifo_iarg_15_dout),
        .ap_fifo_iarg_15_read(ap_fifo_iarg_15_read),
        .s_axis_fifo_16_aclk(s_axis_fifo_16_aclk),
        .s_axis_fifo_16_aresetn(s_axis_fifo_16_aresetn),
        .s_axis_fifo_16_tlast(s_axis_fifo_16_tlast),
        .s_axis_fifo_16_tvalid(s_axis_fifo_16_tvalid),
        .s_axis_fifo_16_tkeep(s_axis_fifo_16_tkeep),
        .s_axis_fifo_16_tstrb(s_axis_fifo_16_tstrb),
        .s_axis_fifo_16_tdata(s_axis_fifo_16_tdata),
        .s_axis_fifo_16_tready(s_axis_fifo_16_tready),
        .ap_fifo_iarg_16_empty_n(ap_fifo_iarg_16_empty_n),
        .ap_fifo_iarg_16_dout(ap_fifo_iarg_16_dout),
        .ap_fifo_iarg_16_read(ap_fifo_iarg_16_read),
        .s_axis_fifo_17_aclk(s_axis_fifo_17_aclk),
        .s_axis_fifo_17_aresetn(s_axis_fifo_17_aresetn),
        .s_axis_fifo_17_tlast(s_axis_fifo_17_tlast),
        .s_axis_fifo_17_tvalid(s_axis_fifo_17_tvalid),
        .s_axis_fifo_17_tkeep(s_axis_fifo_17_tkeep),
        .s_axis_fifo_17_tstrb(s_axis_fifo_17_tstrb),
        .s_axis_fifo_17_tdata(s_axis_fifo_17_tdata),
        .s_axis_fifo_17_tready(s_axis_fifo_17_tready),
        .ap_fifo_iarg_17_empty_n(ap_fifo_iarg_17_empty_n),
        .ap_fifo_iarg_17_dout(ap_fifo_iarg_17_dout),
        .ap_fifo_iarg_17_read(ap_fifo_iarg_17_read),
        .s_axis_fifo_18_aclk(s_axis_fifo_18_aclk),
        .s_axis_fifo_18_aresetn(s_axis_fifo_18_aresetn),
        .s_axis_fifo_18_tlast(s_axis_fifo_18_tlast),
        .s_axis_fifo_18_tvalid(s_axis_fifo_18_tvalid),
        .s_axis_fifo_18_tkeep(s_axis_fifo_18_tkeep),
        .s_axis_fifo_18_tstrb(s_axis_fifo_18_tstrb),
        .s_axis_fifo_18_tdata(s_axis_fifo_18_tdata),
        .s_axis_fifo_18_tready(s_axis_fifo_18_tready),
        .ap_fifo_iarg_18_empty_n(ap_fifo_iarg_18_empty_n),
        .ap_fifo_iarg_18_dout(ap_fifo_iarg_18_dout),
        .ap_fifo_iarg_18_read(ap_fifo_iarg_18_read),
        .s_axis_fifo_19_aclk(s_axis_fifo_19_aclk),
        .s_axis_fifo_19_aresetn(s_axis_fifo_19_aresetn),
        .s_axis_fifo_19_tlast(s_axis_fifo_19_tlast),
        .s_axis_fifo_19_tvalid(s_axis_fifo_19_tvalid),
        .s_axis_fifo_19_tkeep(s_axis_fifo_19_tkeep),
        .s_axis_fifo_19_tstrb(s_axis_fifo_19_tstrb),
        .s_axis_fifo_19_tdata(s_axis_fifo_19_tdata),
        .s_axis_fifo_19_tready(s_axis_fifo_19_tready),
        .ap_fifo_iarg_19_empty_n(ap_fifo_iarg_19_empty_n),
        .ap_fifo_iarg_19_dout(ap_fifo_iarg_19_dout),
        .ap_fifo_iarg_19_read(ap_fifo_iarg_19_read),
        .s_axis_fifo_20_aclk(s_axis_fifo_20_aclk),
        .s_axis_fifo_20_aresetn(s_axis_fifo_20_aresetn),
        .s_axis_fifo_20_tlast(s_axis_fifo_20_tlast),
        .s_axis_fifo_20_tvalid(s_axis_fifo_20_tvalid),
        .s_axis_fifo_20_tkeep(s_axis_fifo_20_tkeep),
        .s_axis_fifo_20_tstrb(s_axis_fifo_20_tstrb),
        .s_axis_fifo_20_tdata(s_axis_fifo_20_tdata),
        .s_axis_fifo_20_tready(s_axis_fifo_20_tready),
        .ap_fifo_iarg_20_empty_n(ap_fifo_iarg_20_empty_n),
        .ap_fifo_iarg_20_dout(ap_fifo_iarg_20_dout),
        .ap_fifo_iarg_20_read(ap_fifo_iarg_20_read),
        .s_axis_fifo_21_aclk(s_axis_fifo_21_aclk),
        .s_axis_fifo_21_aresetn(s_axis_fifo_21_aresetn),
        .s_axis_fifo_21_tlast(s_axis_fifo_21_tlast),
        .s_axis_fifo_21_tvalid(s_axis_fifo_21_tvalid),
        .s_axis_fifo_21_tkeep(s_axis_fifo_21_tkeep),
        .s_axis_fifo_21_tstrb(s_axis_fifo_21_tstrb),
        .s_axis_fifo_21_tdata(s_axis_fifo_21_tdata),
        .s_axis_fifo_21_tready(s_axis_fifo_21_tready),
        .ap_fifo_iarg_21_empty_n(ap_fifo_iarg_21_empty_n),
        .ap_fifo_iarg_21_dout(ap_fifo_iarg_21_dout),
        .ap_fifo_iarg_21_read(ap_fifo_iarg_21_read),
        .s_axis_fifo_22_aclk(s_axis_fifo_22_aclk),
        .s_axis_fifo_22_aresetn(s_axis_fifo_22_aresetn),
        .s_axis_fifo_22_tlast(s_axis_fifo_22_tlast),
        .s_axis_fifo_22_tvalid(s_axis_fifo_22_tvalid),
        .s_axis_fifo_22_tkeep(s_axis_fifo_22_tkeep),
        .s_axis_fifo_22_tstrb(s_axis_fifo_22_tstrb),
        .s_axis_fifo_22_tdata(s_axis_fifo_22_tdata),
        .s_axis_fifo_22_tready(s_axis_fifo_22_tready),
        .ap_fifo_iarg_22_empty_n(ap_fifo_iarg_22_empty_n),
        .ap_fifo_iarg_22_dout(ap_fifo_iarg_22_dout),
        .ap_fifo_iarg_22_read(ap_fifo_iarg_22_read),
        .s_axis_fifo_23_aclk(s_axis_fifo_23_aclk),
        .s_axis_fifo_23_aresetn(s_axis_fifo_23_aresetn),
        .s_axis_fifo_23_tlast(s_axis_fifo_23_tlast),
        .s_axis_fifo_23_tvalid(s_axis_fifo_23_tvalid),
        .s_axis_fifo_23_tkeep(s_axis_fifo_23_tkeep),
        .s_axis_fifo_23_tstrb(s_axis_fifo_23_tstrb),
        .s_axis_fifo_23_tdata(s_axis_fifo_23_tdata),
        .s_axis_fifo_23_tready(s_axis_fifo_23_tready),
        .ap_fifo_iarg_23_empty_n(ap_fifo_iarg_23_empty_n),
        .ap_fifo_iarg_23_dout(ap_fifo_iarg_23_dout),
        .ap_fifo_iarg_23_read(ap_fifo_iarg_23_read),
        .s_axis_fifo_24_aclk(s_axis_fifo_24_aclk),
        .s_axis_fifo_24_aresetn(s_axis_fifo_24_aresetn),
        .s_axis_fifo_24_tlast(s_axis_fifo_24_tlast),
        .s_axis_fifo_24_tvalid(s_axis_fifo_24_tvalid),
        .s_axis_fifo_24_tkeep(s_axis_fifo_24_tkeep),
        .s_axis_fifo_24_tstrb(s_axis_fifo_24_tstrb),
        .s_axis_fifo_24_tdata(s_axis_fifo_24_tdata),
        .s_axis_fifo_24_tready(s_axis_fifo_24_tready),
        .ap_fifo_iarg_24_empty_n(ap_fifo_iarg_24_empty_n),
        .ap_fifo_iarg_24_dout(ap_fifo_iarg_24_dout),
        .ap_fifo_iarg_24_read(ap_fifo_iarg_24_read),
        .s_axis_fifo_25_aclk(s_axis_fifo_25_aclk),
        .s_axis_fifo_25_aresetn(s_axis_fifo_25_aresetn),
        .s_axis_fifo_25_tlast(s_axis_fifo_25_tlast),
        .s_axis_fifo_25_tvalid(s_axis_fifo_25_tvalid),
        .s_axis_fifo_25_tkeep(s_axis_fifo_25_tkeep),
        .s_axis_fifo_25_tstrb(s_axis_fifo_25_tstrb),
        .s_axis_fifo_25_tdata(s_axis_fifo_25_tdata),
        .s_axis_fifo_25_tready(s_axis_fifo_25_tready),
        .ap_fifo_iarg_25_empty_n(ap_fifo_iarg_25_empty_n),
        .ap_fifo_iarg_25_dout(ap_fifo_iarg_25_dout),
        .ap_fifo_iarg_25_read(ap_fifo_iarg_25_read),
        .s_axis_fifo_26_aclk(s_axis_fifo_26_aclk),
        .s_axis_fifo_26_aresetn(s_axis_fifo_26_aresetn),
        .s_axis_fifo_26_tlast(s_axis_fifo_26_tlast),
        .s_axis_fifo_26_tvalid(s_axis_fifo_26_tvalid),
        .s_axis_fifo_26_tkeep(s_axis_fifo_26_tkeep),
        .s_axis_fifo_26_tstrb(s_axis_fifo_26_tstrb),
        .s_axis_fifo_26_tdata(s_axis_fifo_26_tdata),
        .s_axis_fifo_26_tready(s_axis_fifo_26_tready),
        .ap_fifo_iarg_26_empty_n(ap_fifo_iarg_26_empty_n),
        .ap_fifo_iarg_26_dout(ap_fifo_iarg_26_dout),
        .ap_fifo_iarg_26_read(ap_fifo_iarg_26_read),
        .s_axis_fifo_27_aclk(s_axis_fifo_27_aclk),
        .s_axis_fifo_27_aresetn(s_axis_fifo_27_aresetn),
        .s_axis_fifo_27_tlast(s_axis_fifo_27_tlast),
        .s_axis_fifo_27_tvalid(s_axis_fifo_27_tvalid),
        .s_axis_fifo_27_tkeep(s_axis_fifo_27_tkeep),
        .s_axis_fifo_27_tstrb(s_axis_fifo_27_tstrb),
        .s_axis_fifo_27_tdata(s_axis_fifo_27_tdata),
        .s_axis_fifo_27_tready(s_axis_fifo_27_tready),
        .ap_fifo_iarg_27_empty_n(ap_fifo_iarg_27_empty_n),
        .ap_fifo_iarg_27_dout(ap_fifo_iarg_27_dout),
        .ap_fifo_iarg_27_read(ap_fifo_iarg_27_read),
        .s_axis_fifo_28_aclk(s_axis_fifo_28_aclk),
        .s_axis_fifo_28_aresetn(s_axis_fifo_28_aresetn),
        .s_axis_fifo_28_tlast(s_axis_fifo_28_tlast),
        .s_axis_fifo_28_tvalid(s_axis_fifo_28_tvalid),
        .s_axis_fifo_28_tkeep(s_axis_fifo_28_tkeep),
        .s_axis_fifo_28_tstrb(s_axis_fifo_28_tstrb),
        .s_axis_fifo_28_tdata(s_axis_fifo_28_tdata),
        .s_axis_fifo_28_tready(s_axis_fifo_28_tready),
        .ap_fifo_iarg_28_empty_n(ap_fifo_iarg_28_empty_n),
        .ap_fifo_iarg_28_dout(ap_fifo_iarg_28_dout),
        .ap_fifo_iarg_28_read(ap_fifo_iarg_28_read),
        .s_axis_fifo_29_aclk(s_axis_fifo_29_aclk),
        .s_axis_fifo_29_aresetn(s_axis_fifo_29_aresetn),
        .s_axis_fifo_29_tlast(s_axis_fifo_29_tlast),
        .s_axis_fifo_29_tvalid(s_axis_fifo_29_tvalid),
        .s_axis_fifo_29_tkeep(s_axis_fifo_29_tkeep),
        .s_axis_fifo_29_tstrb(s_axis_fifo_29_tstrb),
        .s_axis_fifo_29_tdata(s_axis_fifo_29_tdata),
        .s_axis_fifo_29_tready(s_axis_fifo_29_tready),
        .ap_fifo_iarg_29_empty_n(ap_fifo_iarg_29_empty_n),
        .ap_fifo_iarg_29_dout(ap_fifo_iarg_29_dout),
        .ap_fifo_iarg_29_read(ap_fifo_iarg_29_read),
        .s_axis_fifo_30_aclk(s_axis_fifo_30_aclk),
        .s_axis_fifo_30_aresetn(s_axis_fifo_30_aresetn),
        .s_axis_fifo_30_tlast(s_axis_fifo_30_tlast),
        .s_axis_fifo_30_tvalid(s_axis_fifo_30_tvalid),
        .s_axis_fifo_30_tkeep(s_axis_fifo_30_tkeep),
        .s_axis_fifo_30_tstrb(s_axis_fifo_30_tstrb),
        .s_axis_fifo_30_tdata(s_axis_fifo_30_tdata),
        .s_axis_fifo_30_tready(s_axis_fifo_30_tready),
        .ap_fifo_iarg_30_empty_n(ap_fifo_iarg_30_empty_n),
        .ap_fifo_iarg_30_dout(ap_fifo_iarg_30_dout),
        .ap_fifo_iarg_30_read(ap_fifo_iarg_30_read),
        .s_axis_fifo_31_aclk(s_axis_fifo_31_aclk),
        .s_axis_fifo_31_aresetn(s_axis_fifo_31_aresetn),
        .s_axis_fifo_31_tlast(s_axis_fifo_31_tlast),
        .s_axis_fifo_31_tvalid(s_axis_fifo_31_tvalid),
        .s_axis_fifo_31_tkeep(s_axis_fifo_31_tkeep),
        .s_axis_fifo_31_tstrb(s_axis_fifo_31_tstrb),
        .s_axis_fifo_31_tdata(s_axis_fifo_31_tdata),
        .s_axis_fifo_31_tready(s_axis_fifo_31_tready),
        .ap_fifo_iarg_31_empty_n(ap_fifo_iarg_31_empty_n),
        .ap_fifo_iarg_31_dout(ap_fifo_iarg_31_dout),
        .ap_fifo_iarg_31_read(ap_fifo_iarg_31_read),
        .s_axis_fifo_32_aclk(s_axis_fifo_32_aclk),
        .s_axis_fifo_32_aresetn(s_axis_fifo_32_aresetn),
        .s_axis_fifo_32_tlast(s_axis_fifo_32_tlast),
        .s_axis_fifo_32_tvalid(s_axis_fifo_32_tvalid),
        .s_axis_fifo_32_tkeep(s_axis_fifo_32_tkeep),
        .s_axis_fifo_32_tstrb(s_axis_fifo_32_tstrb),
        .s_axis_fifo_32_tdata(s_axis_fifo_32_tdata),
        .s_axis_fifo_32_tready(s_axis_fifo_32_tready),
        .ap_fifo_iarg_32_empty_n(ap_fifo_iarg_32_empty_n),
        .ap_fifo_iarg_32_dout(ap_fifo_iarg_32_dout),
        .ap_fifo_iarg_32_read(ap_fifo_iarg_32_read),
        .s_axis_fifo_33_aclk(s_axis_fifo_33_aclk),
        .s_axis_fifo_33_aresetn(s_axis_fifo_33_aresetn),
        .s_axis_fifo_33_tlast(s_axis_fifo_33_tlast),
        .s_axis_fifo_33_tvalid(s_axis_fifo_33_tvalid),
        .s_axis_fifo_33_tkeep(s_axis_fifo_33_tkeep),
        .s_axis_fifo_33_tstrb(s_axis_fifo_33_tstrb),
        .s_axis_fifo_33_tdata(s_axis_fifo_33_tdata),
        .s_axis_fifo_33_tready(s_axis_fifo_33_tready),
        .ap_fifo_iarg_33_empty_n(ap_fifo_iarg_33_empty_n),
        .ap_fifo_iarg_33_dout(ap_fifo_iarg_33_dout),
        .ap_fifo_iarg_33_read(ap_fifo_iarg_33_read),
        .s_axis_fifo_34_aclk(s_axis_fifo_34_aclk),
        .s_axis_fifo_34_aresetn(s_axis_fifo_34_aresetn),
        .s_axis_fifo_34_tlast(s_axis_fifo_34_tlast),
        .s_axis_fifo_34_tvalid(s_axis_fifo_34_tvalid),
        .s_axis_fifo_34_tkeep(s_axis_fifo_34_tkeep),
        .s_axis_fifo_34_tstrb(s_axis_fifo_34_tstrb),
        .s_axis_fifo_34_tdata(s_axis_fifo_34_tdata),
        .s_axis_fifo_34_tready(s_axis_fifo_34_tready),
        .ap_fifo_iarg_34_empty_n(ap_fifo_iarg_34_empty_n),
        .ap_fifo_iarg_34_dout(ap_fifo_iarg_34_dout),
        .ap_fifo_iarg_34_read(ap_fifo_iarg_34_read),
        .s_axis_fifo_35_aclk(s_axis_fifo_35_aclk),
        .s_axis_fifo_35_aresetn(s_axis_fifo_35_aresetn),
        .s_axis_fifo_35_tlast(s_axis_fifo_35_tlast),
        .s_axis_fifo_35_tvalid(s_axis_fifo_35_tvalid),
        .s_axis_fifo_35_tkeep(s_axis_fifo_35_tkeep),
        .s_axis_fifo_35_tstrb(s_axis_fifo_35_tstrb),
        .s_axis_fifo_35_tdata(s_axis_fifo_35_tdata),
        .s_axis_fifo_35_tready(s_axis_fifo_35_tready),
        .ap_fifo_iarg_35_empty_n(ap_fifo_iarg_35_empty_n),
        .ap_fifo_iarg_35_dout(ap_fifo_iarg_35_dout),
        .ap_fifo_iarg_35_read(ap_fifo_iarg_35_read),
        .s_axis_fifo_36_aclk(s_axis_fifo_36_aclk),
        .s_axis_fifo_36_aresetn(s_axis_fifo_36_aresetn),
        .s_axis_fifo_36_tlast(s_axis_fifo_36_tlast),
        .s_axis_fifo_36_tvalid(s_axis_fifo_36_tvalid),
        .s_axis_fifo_36_tkeep(s_axis_fifo_36_tkeep),
        .s_axis_fifo_36_tstrb(s_axis_fifo_36_tstrb),
        .s_axis_fifo_36_tdata(s_axis_fifo_36_tdata),
        .s_axis_fifo_36_tready(s_axis_fifo_36_tready),
        .ap_fifo_iarg_36_empty_n(ap_fifo_iarg_36_empty_n),
        .ap_fifo_iarg_36_dout(ap_fifo_iarg_36_dout),
        .ap_fifo_iarg_36_read(ap_fifo_iarg_36_read),
        .s_axis_fifo_37_aclk(s_axis_fifo_37_aclk),
        .s_axis_fifo_37_aresetn(s_axis_fifo_37_aresetn),
        .s_axis_fifo_37_tlast(s_axis_fifo_37_tlast),
        .s_axis_fifo_37_tvalid(s_axis_fifo_37_tvalid),
        .s_axis_fifo_37_tkeep(s_axis_fifo_37_tkeep),
        .s_axis_fifo_37_tstrb(s_axis_fifo_37_tstrb),
        .s_axis_fifo_37_tdata(s_axis_fifo_37_tdata),
        .s_axis_fifo_37_tready(s_axis_fifo_37_tready),
        .ap_fifo_iarg_37_empty_n(ap_fifo_iarg_37_empty_n),
        .ap_fifo_iarg_37_dout(ap_fifo_iarg_37_dout),
        .ap_fifo_iarg_37_read(ap_fifo_iarg_37_read),
        .s_axis_fifo_38_aclk(s_axis_fifo_38_aclk),
        .s_axis_fifo_38_aresetn(s_axis_fifo_38_aresetn),
        .s_axis_fifo_38_tlast(s_axis_fifo_38_tlast),
        .s_axis_fifo_38_tvalid(s_axis_fifo_38_tvalid),
        .s_axis_fifo_38_tkeep(s_axis_fifo_38_tkeep),
        .s_axis_fifo_38_tstrb(s_axis_fifo_38_tstrb),
        .s_axis_fifo_38_tdata(s_axis_fifo_38_tdata),
        .s_axis_fifo_38_tready(s_axis_fifo_38_tready),
        .ap_fifo_iarg_38_empty_n(ap_fifo_iarg_38_empty_n),
        .ap_fifo_iarg_38_dout(ap_fifo_iarg_38_dout),
        .ap_fifo_iarg_38_read(ap_fifo_iarg_38_read),
        .s_axis_fifo_39_aclk(s_axis_fifo_39_aclk),
        .s_axis_fifo_39_aresetn(s_axis_fifo_39_aresetn),
        .s_axis_fifo_39_tlast(s_axis_fifo_39_tlast),
        .s_axis_fifo_39_tvalid(s_axis_fifo_39_tvalid),
        .s_axis_fifo_39_tkeep(s_axis_fifo_39_tkeep),
        .s_axis_fifo_39_tstrb(s_axis_fifo_39_tstrb),
        .s_axis_fifo_39_tdata(s_axis_fifo_39_tdata),
        .s_axis_fifo_39_tready(s_axis_fifo_39_tready),
        .ap_fifo_iarg_39_empty_n(ap_fifo_iarg_39_empty_n),
        .ap_fifo_iarg_39_dout(ap_fifo_iarg_39_dout),
        .ap_fifo_iarg_39_read(ap_fifo_iarg_39_read),
        .s_axis_fifo_40_aclk(s_axis_fifo_40_aclk),
        .s_axis_fifo_40_aresetn(s_axis_fifo_40_aresetn),
        .s_axis_fifo_40_tlast(s_axis_fifo_40_tlast),
        .s_axis_fifo_40_tvalid(s_axis_fifo_40_tvalid),
        .s_axis_fifo_40_tkeep(s_axis_fifo_40_tkeep),
        .s_axis_fifo_40_tstrb(s_axis_fifo_40_tstrb),
        .s_axis_fifo_40_tdata(s_axis_fifo_40_tdata),
        .s_axis_fifo_40_tready(s_axis_fifo_40_tready),
        .ap_fifo_iarg_40_empty_n(ap_fifo_iarg_40_empty_n),
        .ap_fifo_iarg_40_dout(ap_fifo_iarg_40_dout),
        .ap_fifo_iarg_40_read(ap_fifo_iarg_40_read),
        .s_axis_fifo_41_aclk(s_axis_fifo_41_aclk),
        .s_axis_fifo_41_aresetn(s_axis_fifo_41_aresetn),
        .s_axis_fifo_41_tlast(s_axis_fifo_41_tlast),
        .s_axis_fifo_41_tvalid(s_axis_fifo_41_tvalid),
        .s_axis_fifo_41_tkeep(s_axis_fifo_41_tkeep),
        .s_axis_fifo_41_tstrb(s_axis_fifo_41_tstrb),
        .s_axis_fifo_41_tdata(s_axis_fifo_41_tdata),
        .s_axis_fifo_41_tready(s_axis_fifo_41_tready),
        .ap_fifo_iarg_41_empty_n(ap_fifo_iarg_41_empty_n),
        .ap_fifo_iarg_41_dout(ap_fifo_iarg_41_dout),
        .ap_fifo_iarg_41_read(ap_fifo_iarg_41_read),
        .s_axis_fifo_42_aclk(s_axis_fifo_42_aclk),
        .s_axis_fifo_42_aresetn(s_axis_fifo_42_aresetn),
        .s_axis_fifo_42_tlast(s_axis_fifo_42_tlast),
        .s_axis_fifo_42_tvalid(s_axis_fifo_42_tvalid),
        .s_axis_fifo_42_tkeep(s_axis_fifo_42_tkeep),
        .s_axis_fifo_42_tstrb(s_axis_fifo_42_tstrb),
        .s_axis_fifo_42_tdata(s_axis_fifo_42_tdata),
        .s_axis_fifo_42_tready(s_axis_fifo_42_tready),
        .ap_fifo_iarg_42_empty_n(ap_fifo_iarg_42_empty_n),
        .ap_fifo_iarg_42_dout(ap_fifo_iarg_42_dout),
        .ap_fifo_iarg_42_read(ap_fifo_iarg_42_read),
        .s_axis_fifo_43_aclk(s_axis_fifo_43_aclk),
        .s_axis_fifo_43_aresetn(s_axis_fifo_43_aresetn),
        .s_axis_fifo_43_tlast(s_axis_fifo_43_tlast),
        .s_axis_fifo_43_tvalid(s_axis_fifo_43_tvalid),
        .s_axis_fifo_43_tkeep(s_axis_fifo_43_tkeep),
        .s_axis_fifo_43_tstrb(s_axis_fifo_43_tstrb),
        .s_axis_fifo_43_tdata(s_axis_fifo_43_tdata),
        .s_axis_fifo_43_tready(s_axis_fifo_43_tready),
        .ap_fifo_iarg_43_empty_n(ap_fifo_iarg_43_empty_n),
        .ap_fifo_iarg_43_dout(ap_fifo_iarg_43_dout),
        .ap_fifo_iarg_43_read(ap_fifo_iarg_43_read),
        .s_axis_fifo_44_aclk(s_axis_fifo_44_aclk),
        .s_axis_fifo_44_aresetn(s_axis_fifo_44_aresetn),
        .s_axis_fifo_44_tlast(s_axis_fifo_44_tlast),
        .s_axis_fifo_44_tvalid(s_axis_fifo_44_tvalid),
        .s_axis_fifo_44_tkeep(s_axis_fifo_44_tkeep),
        .s_axis_fifo_44_tstrb(s_axis_fifo_44_tstrb),
        .s_axis_fifo_44_tdata(s_axis_fifo_44_tdata),
        .s_axis_fifo_44_tready(s_axis_fifo_44_tready),
        .ap_fifo_iarg_44_empty_n(ap_fifo_iarg_44_empty_n),
        .ap_fifo_iarg_44_dout(ap_fifo_iarg_44_dout),
        .ap_fifo_iarg_44_read(ap_fifo_iarg_44_read),
        .s_axis_fifo_45_aclk(s_axis_fifo_45_aclk),
        .s_axis_fifo_45_aresetn(s_axis_fifo_45_aresetn),
        .s_axis_fifo_45_tlast(s_axis_fifo_45_tlast),
        .s_axis_fifo_45_tvalid(s_axis_fifo_45_tvalid),
        .s_axis_fifo_45_tkeep(s_axis_fifo_45_tkeep),
        .s_axis_fifo_45_tstrb(s_axis_fifo_45_tstrb),
        .s_axis_fifo_45_tdata(s_axis_fifo_45_tdata),
        .s_axis_fifo_45_tready(s_axis_fifo_45_tready),
        .ap_fifo_iarg_45_empty_n(ap_fifo_iarg_45_empty_n),
        .ap_fifo_iarg_45_dout(ap_fifo_iarg_45_dout),
        .ap_fifo_iarg_45_read(ap_fifo_iarg_45_read),
        .s_axis_fifo_46_aclk(s_axis_fifo_46_aclk),
        .s_axis_fifo_46_aresetn(s_axis_fifo_46_aresetn),
        .s_axis_fifo_46_tlast(s_axis_fifo_46_tlast),
        .s_axis_fifo_46_tvalid(s_axis_fifo_46_tvalid),
        .s_axis_fifo_46_tkeep(s_axis_fifo_46_tkeep),
        .s_axis_fifo_46_tstrb(s_axis_fifo_46_tstrb),
        .s_axis_fifo_46_tdata(s_axis_fifo_46_tdata),
        .s_axis_fifo_46_tready(s_axis_fifo_46_tready),
        .ap_fifo_iarg_46_empty_n(ap_fifo_iarg_46_empty_n),
        .ap_fifo_iarg_46_dout(ap_fifo_iarg_46_dout),
        .ap_fifo_iarg_46_read(ap_fifo_iarg_46_read),
        .s_axis_fifo_47_aclk(s_axis_fifo_47_aclk),
        .s_axis_fifo_47_aresetn(s_axis_fifo_47_aresetn),
        .s_axis_fifo_47_tlast(s_axis_fifo_47_tlast),
        .s_axis_fifo_47_tvalid(s_axis_fifo_47_tvalid),
        .s_axis_fifo_47_tkeep(s_axis_fifo_47_tkeep),
        .s_axis_fifo_47_tstrb(s_axis_fifo_47_tstrb),
        .s_axis_fifo_47_tdata(s_axis_fifo_47_tdata),
        .s_axis_fifo_47_tready(s_axis_fifo_47_tready),
        .ap_fifo_iarg_47_empty_n(ap_fifo_iarg_47_empty_n),
        .ap_fifo_iarg_47_dout(ap_fifo_iarg_47_dout),
        .ap_fifo_iarg_47_read(ap_fifo_iarg_47_read),
        .s_axis_fifo_48_aclk(s_axis_fifo_48_aclk),
        .s_axis_fifo_48_aresetn(s_axis_fifo_48_aresetn),
        .s_axis_fifo_48_tlast(s_axis_fifo_48_tlast),
        .s_axis_fifo_48_tvalid(s_axis_fifo_48_tvalid),
        .s_axis_fifo_48_tkeep(s_axis_fifo_48_tkeep),
        .s_axis_fifo_48_tstrb(s_axis_fifo_48_tstrb),
        .s_axis_fifo_48_tdata(s_axis_fifo_48_tdata),
        .s_axis_fifo_48_tready(s_axis_fifo_48_tready),
        .ap_fifo_iarg_48_empty_n(ap_fifo_iarg_48_empty_n),
        .ap_fifo_iarg_48_dout(ap_fifo_iarg_48_dout),
        .ap_fifo_iarg_48_read(ap_fifo_iarg_48_read),
        .s_axis_fifo_49_aclk(s_axis_fifo_49_aclk),
        .s_axis_fifo_49_aresetn(s_axis_fifo_49_aresetn),
        .s_axis_fifo_49_tlast(s_axis_fifo_49_tlast),
        .s_axis_fifo_49_tvalid(s_axis_fifo_49_tvalid),
        .s_axis_fifo_49_tkeep(s_axis_fifo_49_tkeep),
        .s_axis_fifo_49_tstrb(s_axis_fifo_49_tstrb),
        .s_axis_fifo_49_tdata(s_axis_fifo_49_tdata),
        .s_axis_fifo_49_tready(s_axis_fifo_49_tready),
        .ap_fifo_iarg_49_empty_n(ap_fifo_iarg_49_empty_n),
        .ap_fifo_iarg_49_dout(ap_fifo_iarg_49_dout),
        .ap_fifo_iarg_49_read(ap_fifo_iarg_49_read),
        .s_axis_fifo_50_aclk(s_axis_fifo_50_aclk),
        .s_axis_fifo_50_aresetn(s_axis_fifo_50_aresetn),
        .s_axis_fifo_50_tlast(s_axis_fifo_50_tlast),
        .s_axis_fifo_50_tvalid(s_axis_fifo_50_tvalid),
        .s_axis_fifo_50_tkeep(s_axis_fifo_50_tkeep),
        .s_axis_fifo_50_tstrb(s_axis_fifo_50_tstrb),
        .s_axis_fifo_50_tdata(s_axis_fifo_50_tdata),
        .s_axis_fifo_50_tready(s_axis_fifo_50_tready),
        .ap_fifo_iarg_50_empty_n(ap_fifo_iarg_50_empty_n),
        .ap_fifo_iarg_50_dout(ap_fifo_iarg_50_dout),
        .ap_fifo_iarg_50_read(ap_fifo_iarg_50_read),
        .s_axis_fifo_51_aclk(s_axis_fifo_51_aclk),
        .s_axis_fifo_51_aresetn(s_axis_fifo_51_aresetn),
        .s_axis_fifo_51_tlast(s_axis_fifo_51_tlast),
        .s_axis_fifo_51_tvalid(s_axis_fifo_51_tvalid),
        .s_axis_fifo_51_tkeep(s_axis_fifo_51_tkeep),
        .s_axis_fifo_51_tstrb(s_axis_fifo_51_tstrb),
        .s_axis_fifo_51_tdata(s_axis_fifo_51_tdata),
        .s_axis_fifo_51_tready(s_axis_fifo_51_tready),
        .ap_fifo_iarg_51_empty_n(ap_fifo_iarg_51_empty_n),
        .ap_fifo_iarg_51_dout(ap_fifo_iarg_51_dout),
        .ap_fifo_iarg_51_read(ap_fifo_iarg_51_read),
        .s_axis_fifo_52_aclk(s_axis_fifo_52_aclk),
        .s_axis_fifo_52_aresetn(s_axis_fifo_52_aresetn),
        .s_axis_fifo_52_tlast(s_axis_fifo_52_tlast),
        .s_axis_fifo_52_tvalid(s_axis_fifo_52_tvalid),
        .s_axis_fifo_52_tkeep(s_axis_fifo_52_tkeep),
        .s_axis_fifo_52_tstrb(s_axis_fifo_52_tstrb),
        .s_axis_fifo_52_tdata(s_axis_fifo_52_tdata),
        .s_axis_fifo_52_tready(s_axis_fifo_52_tready),
        .ap_fifo_iarg_52_empty_n(ap_fifo_iarg_52_empty_n),
        .ap_fifo_iarg_52_dout(ap_fifo_iarg_52_dout),
        .ap_fifo_iarg_52_read(ap_fifo_iarg_52_read),
        .s_axis_fifo_53_aclk(s_axis_fifo_53_aclk),
        .s_axis_fifo_53_aresetn(s_axis_fifo_53_aresetn),
        .s_axis_fifo_53_tlast(s_axis_fifo_53_tlast),
        .s_axis_fifo_53_tvalid(s_axis_fifo_53_tvalid),
        .s_axis_fifo_53_tkeep(s_axis_fifo_53_tkeep),
        .s_axis_fifo_53_tstrb(s_axis_fifo_53_tstrb),
        .s_axis_fifo_53_tdata(s_axis_fifo_53_tdata),
        .s_axis_fifo_53_tready(s_axis_fifo_53_tready),
        .ap_fifo_iarg_53_empty_n(ap_fifo_iarg_53_empty_n),
        .ap_fifo_iarg_53_dout(ap_fifo_iarg_53_dout),
        .ap_fifo_iarg_53_read(ap_fifo_iarg_53_read),
        .s_axis_fifo_54_aclk(s_axis_fifo_54_aclk),
        .s_axis_fifo_54_aresetn(s_axis_fifo_54_aresetn),
        .s_axis_fifo_54_tlast(s_axis_fifo_54_tlast),
        .s_axis_fifo_54_tvalid(s_axis_fifo_54_tvalid),
        .s_axis_fifo_54_tkeep(s_axis_fifo_54_tkeep),
        .s_axis_fifo_54_tstrb(s_axis_fifo_54_tstrb),
        .s_axis_fifo_54_tdata(s_axis_fifo_54_tdata),
        .s_axis_fifo_54_tready(s_axis_fifo_54_tready),
        .ap_fifo_iarg_54_empty_n(ap_fifo_iarg_54_empty_n),
        .ap_fifo_iarg_54_dout(ap_fifo_iarg_54_dout),
        .ap_fifo_iarg_54_read(ap_fifo_iarg_54_read),
        .s_axis_fifo_55_aclk(s_axis_fifo_55_aclk),
        .s_axis_fifo_55_aresetn(s_axis_fifo_55_aresetn),
        .s_axis_fifo_55_tlast(s_axis_fifo_55_tlast),
        .s_axis_fifo_55_tvalid(s_axis_fifo_55_tvalid),
        .s_axis_fifo_55_tkeep(s_axis_fifo_55_tkeep),
        .s_axis_fifo_55_tstrb(s_axis_fifo_55_tstrb),
        .s_axis_fifo_55_tdata(s_axis_fifo_55_tdata),
        .s_axis_fifo_55_tready(s_axis_fifo_55_tready),
        .ap_fifo_iarg_55_empty_n(ap_fifo_iarg_55_empty_n),
        .ap_fifo_iarg_55_dout(ap_fifo_iarg_55_dout),
        .ap_fifo_iarg_55_read(ap_fifo_iarg_55_read),
        .s_axis_fifo_56_aclk(s_axis_fifo_56_aclk),
        .s_axis_fifo_56_aresetn(s_axis_fifo_56_aresetn),
        .s_axis_fifo_56_tlast(s_axis_fifo_56_tlast),
        .s_axis_fifo_56_tvalid(s_axis_fifo_56_tvalid),
        .s_axis_fifo_56_tkeep(s_axis_fifo_56_tkeep),
        .s_axis_fifo_56_tstrb(s_axis_fifo_56_tstrb),
        .s_axis_fifo_56_tdata(s_axis_fifo_56_tdata),
        .s_axis_fifo_56_tready(s_axis_fifo_56_tready),
        .ap_fifo_iarg_56_empty_n(ap_fifo_iarg_56_empty_n),
        .ap_fifo_iarg_56_dout(ap_fifo_iarg_56_dout),
        .ap_fifo_iarg_56_read(ap_fifo_iarg_56_read),
        .s_axis_fifo_57_aclk(s_axis_fifo_57_aclk),
        .s_axis_fifo_57_aresetn(s_axis_fifo_57_aresetn),
        .s_axis_fifo_57_tlast(s_axis_fifo_57_tlast),
        .s_axis_fifo_57_tvalid(s_axis_fifo_57_tvalid),
        .s_axis_fifo_57_tkeep(s_axis_fifo_57_tkeep),
        .s_axis_fifo_57_tstrb(s_axis_fifo_57_tstrb),
        .s_axis_fifo_57_tdata(s_axis_fifo_57_tdata),
        .s_axis_fifo_57_tready(s_axis_fifo_57_tready),
        .ap_fifo_iarg_57_empty_n(ap_fifo_iarg_57_empty_n),
        .ap_fifo_iarg_57_dout(ap_fifo_iarg_57_dout),
        .ap_fifo_iarg_57_read(ap_fifo_iarg_57_read),
        .s_axis_fifo_58_aclk(s_axis_fifo_58_aclk),
        .s_axis_fifo_58_aresetn(s_axis_fifo_58_aresetn),
        .s_axis_fifo_58_tlast(s_axis_fifo_58_tlast),
        .s_axis_fifo_58_tvalid(s_axis_fifo_58_tvalid),
        .s_axis_fifo_58_tkeep(s_axis_fifo_58_tkeep),
        .s_axis_fifo_58_tstrb(s_axis_fifo_58_tstrb),
        .s_axis_fifo_58_tdata(s_axis_fifo_58_tdata),
        .s_axis_fifo_58_tready(s_axis_fifo_58_tready),
        .ap_fifo_iarg_58_empty_n(ap_fifo_iarg_58_empty_n),
        .ap_fifo_iarg_58_dout(ap_fifo_iarg_58_dout),
        .ap_fifo_iarg_58_read(ap_fifo_iarg_58_read),
        .s_axis_fifo_59_aclk(s_axis_fifo_59_aclk),
        .s_axis_fifo_59_aresetn(s_axis_fifo_59_aresetn),
        .s_axis_fifo_59_tlast(s_axis_fifo_59_tlast),
        .s_axis_fifo_59_tvalid(s_axis_fifo_59_tvalid),
        .s_axis_fifo_59_tkeep(s_axis_fifo_59_tkeep),
        .s_axis_fifo_59_tstrb(s_axis_fifo_59_tstrb),
        .s_axis_fifo_59_tdata(s_axis_fifo_59_tdata),
        .s_axis_fifo_59_tready(s_axis_fifo_59_tready),
        .ap_fifo_iarg_59_empty_n(ap_fifo_iarg_59_empty_n),
        .ap_fifo_iarg_59_dout(ap_fifo_iarg_59_dout),
        .ap_fifo_iarg_59_read(ap_fifo_iarg_59_read),
        .s_axis_fifo_60_aclk(s_axis_fifo_60_aclk),
        .s_axis_fifo_60_aresetn(s_axis_fifo_60_aresetn),
        .s_axis_fifo_60_tlast(s_axis_fifo_60_tlast),
        .s_axis_fifo_60_tvalid(s_axis_fifo_60_tvalid),
        .s_axis_fifo_60_tkeep(s_axis_fifo_60_tkeep),
        .s_axis_fifo_60_tstrb(s_axis_fifo_60_tstrb),
        .s_axis_fifo_60_tdata(s_axis_fifo_60_tdata),
        .s_axis_fifo_60_tready(s_axis_fifo_60_tready),
        .ap_fifo_iarg_60_empty_n(ap_fifo_iarg_60_empty_n),
        .ap_fifo_iarg_60_dout(ap_fifo_iarg_60_dout),
        .ap_fifo_iarg_60_read(ap_fifo_iarg_60_read),
        .s_axis_fifo_61_aclk(s_axis_fifo_61_aclk),
        .s_axis_fifo_61_aresetn(s_axis_fifo_61_aresetn),
        .s_axis_fifo_61_tlast(s_axis_fifo_61_tlast),
        .s_axis_fifo_61_tvalid(s_axis_fifo_61_tvalid),
        .s_axis_fifo_61_tkeep(s_axis_fifo_61_tkeep),
        .s_axis_fifo_61_tstrb(s_axis_fifo_61_tstrb),
        .s_axis_fifo_61_tdata(s_axis_fifo_61_tdata),
        .s_axis_fifo_61_tready(s_axis_fifo_61_tready),
        .ap_fifo_iarg_61_empty_n(ap_fifo_iarg_61_empty_n),
        .ap_fifo_iarg_61_dout(ap_fifo_iarg_61_dout),
        .ap_fifo_iarg_61_read(ap_fifo_iarg_61_read),
        .s_axis_fifo_62_aclk(s_axis_fifo_62_aclk),
        .s_axis_fifo_62_aresetn(s_axis_fifo_62_aresetn),
        .s_axis_fifo_62_tlast(s_axis_fifo_62_tlast),
        .s_axis_fifo_62_tvalid(s_axis_fifo_62_tvalid),
        .s_axis_fifo_62_tkeep(s_axis_fifo_62_tkeep),
        .s_axis_fifo_62_tstrb(s_axis_fifo_62_tstrb),
        .s_axis_fifo_62_tdata(s_axis_fifo_62_tdata),
        .s_axis_fifo_62_tready(s_axis_fifo_62_tready),
        .ap_fifo_iarg_62_empty_n(ap_fifo_iarg_62_empty_n),
        .ap_fifo_iarg_62_dout(ap_fifo_iarg_62_dout),
        .ap_fifo_iarg_62_read(ap_fifo_iarg_62_read),
        .s_axis_fifo_63_aclk(s_axis_fifo_63_aclk),
        .s_axis_fifo_63_aresetn(s_axis_fifo_63_aresetn),
        .s_axis_fifo_63_tlast(s_axis_fifo_63_tlast),
        .s_axis_fifo_63_tvalid(s_axis_fifo_63_tvalid),
        .s_axis_fifo_63_tkeep(s_axis_fifo_63_tkeep),
        .s_axis_fifo_63_tstrb(s_axis_fifo_63_tstrb),
        .s_axis_fifo_63_tdata(s_axis_fifo_63_tdata),
        .s_axis_fifo_63_tready(s_axis_fifo_63_tready),
        .ap_fifo_iarg_63_empty_n(ap_fifo_iarg_63_empty_n),
        .ap_fifo_iarg_63_dout(ap_fifo_iarg_63_dout),
        .ap_fifo_iarg_63_read(ap_fifo_iarg_63_read),
        .s_axis_fifo_64_aclk(s_axis_fifo_64_aclk),
        .s_axis_fifo_64_aresetn(s_axis_fifo_64_aresetn),
        .s_axis_fifo_64_tlast(s_axis_fifo_64_tlast),
        .s_axis_fifo_64_tvalid(s_axis_fifo_64_tvalid),
        .s_axis_fifo_64_tkeep(s_axis_fifo_64_tkeep),
        .s_axis_fifo_64_tstrb(s_axis_fifo_64_tstrb),
        .s_axis_fifo_64_tdata(s_axis_fifo_64_tdata),
        .s_axis_fifo_64_tready(s_axis_fifo_64_tready),
        .ap_fifo_iarg_64_empty_n(ap_fifo_iarg_64_empty_n),
        .ap_fifo_iarg_64_dout(ap_fifo_iarg_64_dout),
        .ap_fifo_iarg_64_read(ap_fifo_iarg_64_read),
        .s_axis_fifo_65_aclk(s_axis_fifo_65_aclk),
        .s_axis_fifo_65_aresetn(s_axis_fifo_65_aresetn),
        .s_axis_fifo_65_tlast(s_axis_fifo_65_tlast),
        .s_axis_fifo_65_tvalid(s_axis_fifo_65_tvalid),
        .s_axis_fifo_65_tkeep(s_axis_fifo_65_tkeep),
        .s_axis_fifo_65_tstrb(s_axis_fifo_65_tstrb),
        .s_axis_fifo_65_tdata(s_axis_fifo_65_tdata),
        .s_axis_fifo_65_tready(s_axis_fifo_65_tready),
        .ap_fifo_iarg_65_empty_n(ap_fifo_iarg_65_empty_n),
        .ap_fifo_iarg_65_dout(ap_fifo_iarg_65_dout),
        .ap_fifo_iarg_65_read(ap_fifo_iarg_65_read),
        .s_axis_fifo_66_aclk(s_axis_fifo_66_aclk),
        .s_axis_fifo_66_aresetn(s_axis_fifo_66_aresetn),
        .s_axis_fifo_66_tlast(s_axis_fifo_66_tlast),
        .s_axis_fifo_66_tvalid(s_axis_fifo_66_tvalid),
        .s_axis_fifo_66_tkeep(s_axis_fifo_66_tkeep),
        .s_axis_fifo_66_tstrb(s_axis_fifo_66_tstrb),
        .s_axis_fifo_66_tdata(s_axis_fifo_66_tdata),
        .s_axis_fifo_66_tready(s_axis_fifo_66_tready),
        .ap_fifo_iarg_66_empty_n(ap_fifo_iarg_66_empty_n),
        .ap_fifo_iarg_66_dout(ap_fifo_iarg_66_dout),
        .ap_fifo_iarg_66_read(ap_fifo_iarg_66_read),
        .s_axis_fifo_67_aclk(s_axis_fifo_67_aclk),
        .s_axis_fifo_67_aresetn(s_axis_fifo_67_aresetn),
        .s_axis_fifo_67_tlast(s_axis_fifo_67_tlast),
        .s_axis_fifo_67_tvalid(s_axis_fifo_67_tvalid),
        .s_axis_fifo_67_tkeep(s_axis_fifo_67_tkeep),
        .s_axis_fifo_67_tstrb(s_axis_fifo_67_tstrb),
        .s_axis_fifo_67_tdata(s_axis_fifo_67_tdata),
        .s_axis_fifo_67_tready(s_axis_fifo_67_tready),
        .ap_fifo_iarg_67_empty_n(ap_fifo_iarg_67_empty_n),
        .ap_fifo_iarg_67_dout(ap_fifo_iarg_67_dout),
        .ap_fifo_iarg_67_read(ap_fifo_iarg_67_read),
        .s_axis_fifo_68_aclk(s_axis_fifo_68_aclk),
        .s_axis_fifo_68_aresetn(s_axis_fifo_68_aresetn),
        .s_axis_fifo_68_tlast(s_axis_fifo_68_tlast),
        .s_axis_fifo_68_tvalid(s_axis_fifo_68_tvalid),
        .s_axis_fifo_68_tkeep(s_axis_fifo_68_tkeep),
        .s_axis_fifo_68_tstrb(s_axis_fifo_68_tstrb),
        .s_axis_fifo_68_tdata(s_axis_fifo_68_tdata),
        .s_axis_fifo_68_tready(s_axis_fifo_68_tready),
        .ap_fifo_iarg_68_empty_n(ap_fifo_iarg_68_empty_n),
        .ap_fifo_iarg_68_dout(ap_fifo_iarg_68_dout),
        .ap_fifo_iarg_68_read(ap_fifo_iarg_68_read),
        .s_axis_fifo_69_aclk(s_axis_fifo_69_aclk),
        .s_axis_fifo_69_aresetn(s_axis_fifo_69_aresetn),
        .s_axis_fifo_69_tlast(s_axis_fifo_69_tlast),
        .s_axis_fifo_69_tvalid(s_axis_fifo_69_tvalid),
        .s_axis_fifo_69_tkeep(s_axis_fifo_69_tkeep),
        .s_axis_fifo_69_tstrb(s_axis_fifo_69_tstrb),
        .s_axis_fifo_69_tdata(s_axis_fifo_69_tdata),
        .s_axis_fifo_69_tready(s_axis_fifo_69_tready),
        .ap_fifo_iarg_69_empty_n(ap_fifo_iarg_69_empty_n),
        .ap_fifo_iarg_69_dout(ap_fifo_iarg_69_dout),
        .ap_fifo_iarg_69_read(ap_fifo_iarg_69_read),
        .s_axis_fifo_70_aclk(s_axis_fifo_70_aclk),
        .s_axis_fifo_70_aresetn(s_axis_fifo_70_aresetn),
        .s_axis_fifo_70_tlast(s_axis_fifo_70_tlast),
        .s_axis_fifo_70_tvalid(s_axis_fifo_70_tvalid),
        .s_axis_fifo_70_tkeep(s_axis_fifo_70_tkeep),
        .s_axis_fifo_70_tstrb(s_axis_fifo_70_tstrb),
        .s_axis_fifo_70_tdata(s_axis_fifo_70_tdata),
        .s_axis_fifo_70_tready(s_axis_fifo_70_tready),
        .ap_fifo_iarg_70_empty_n(ap_fifo_iarg_70_empty_n),
        .ap_fifo_iarg_70_dout(ap_fifo_iarg_70_dout),
        .ap_fifo_iarg_70_read(ap_fifo_iarg_70_read),
        .s_axis_fifo_71_aclk(s_axis_fifo_71_aclk),
        .s_axis_fifo_71_aresetn(s_axis_fifo_71_aresetn),
        .s_axis_fifo_71_tlast(s_axis_fifo_71_tlast),
        .s_axis_fifo_71_tvalid(s_axis_fifo_71_tvalid),
        .s_axis_fifo_71_tkeep(s_axis_fifo_71_tkeep),
        .s_axis_fifo_71_tstrb(s_axis_fifo_71_tstrb),
        .s_axis_fifo_71_tdata(s_axis_fifo_71_tdata),
        .s_axis_fifo_71_tready(s_axis_fifo_71_tready),
        .ap_fifo_iarg_71_empty_n(ap_fifo_iarg_71_empty_n),
        .ap_fifo_iarg_71_dout(ap_fifo_iarg_71_dout),
        .ap_fifo_iarg_71_read(ap_fifo_iarg_71_read),
        .s_axis_fifo_72_aclk(s_axis_fifo_72_aclk),
        .s_axis_fifo_72_aresetn(s_axis_fifo_72_aresetn),
        .s_axis_fifo_72_tlast(s_axis_fifo_72_tlast),
        .s_axis_fifo_72_tvalid(s_axis_fifo_72_tvalid),
        .s_axis_fifo_72_tkeep(s_axis_fifo_72_tkeep),
        .s_axis_fifo_72_tstrb(s_axis_fifo_72_tstrb),
        .s_axis_fifo_72_tdata(s_axis_fifo_72_tdata),
        .s_axis_fifo_72_tready(s_axis_fifo_72_tready),
        .ap_fifo_iarg_72_empty_n(ap_fifo_iarg_72_empty_n),
        .ap_fifo_iarg_72_dout(ap_fifo_iarg_72_dout),
        .ap_fifo_iarg_72_read(ap_fifo_iarg_72_read),
        .s_axis_fifo_73_aclk(s_axis_fifo_73_aclk),
        .s_axis_fifo_73_aresetn(s_axis_fifo_73_aresetn),
        .s_axis_fifo_73_tlast(s_axis_fifo_73_tlast),
        .s_axis_fifo_73_tvalid(s_axis_fifo_73_tvalid),
        .s_axis_fifo_73_tkeep(s_axis_fifo_73_tkeep),
        .s_axis_fifo_73_tstrb(s_axis_fifo_73_tstrb),
        .s_axis_fifo_73_tdata(s_axis_fifo_73_tdata),
        .s_axis_fifo_73_tready(s_axis_fifo_73_tready),
        .ap_fifo_iarg_73_empty_n(ap_fifo_iarg_73_empty_n),
        .ap_fifo_iarg_73_dout(ap_fifo_iarg_73_dout),
        .ap_fifo_iarg_73_read(ap_fifo_iarg_73_read),
        .s_axis_fifo_74_aclk(s_axis_fifo_74_aclk),
        .s_axis_fifo_74_aresetn(s_axis_fifo_74_aresetn),
        .s_axis_fifo_74_tlast(s_axis_fifo_74_tlast),
        .s_axis_fifo_74_tvalid(s_axis_fifo_74_tvalid),
        .s_axis_fifo_74_tkeep(s_axis_fifo_74_tkeep),
        .s_axis_fifo_74_tstrb(s_axis_fifo_74_tstrb),
        .s_axis_fifo_74_tdata(s_axis_fifo_74_tdata),
        .s_axis_fifo_74_tready(s_axis_fifo_74_tready),
        .ap_fifo_iarg_74_empty_n(ap_fifo_iarg_74_empty_n),
        .ap_fifo_iarg_74_dout(ap_fifo_iarg_74_dout),
        .ap_fifo_iarg_74_read(ap_fifo_iarg_74_read),
        .s_axis_fifo_75_aclk(s_axis_fifo_75_aclk),
        .s_axis_fifo_75_aresetn(s_axis_fifo_75_aresetn),
        .s_axis_fifo_75_tlast(s_axis_fifo_75_tlast),
        .s_axis_fifo_75_tvalid(s_axis_fifo_75_tvalid),
        .s_axis_fifo_75_tkeep(s_axis_fifo_75_tkeep),
        .s_axis_fifo_75_tstrb(s_axis_fifo_75_tstrb),
        .s_axis_fifo_75_tdata(s_axis_fifo_75_tdata),
        .s_axis_fifo_75_tready(s_axis_fifo_75_tready),
        .ap_fifo_iarg_75_empty_n(ap_fifo_iarg_75_empty_n),
        .ap_fifo_iarg_75_dout(ap_fifo_iarg_75_dout),
        .ap_fifo_iarg_75_read(ap_fifo_iarg_75_read),
        .s_axis_fifo_76_aclk(s_axis_fifo_76_aclk),
        .s_axis_fifo_76_aresetn(s_axis_fifo_76_aresetn),
        .s_axis_fifo_76_tlast(s_axis_fifo_76_tlast),
        .s_axis_fifo_76_tvalid(s_axis_fifo_76_tvalid),
        .s_axis_fifo_76_tkeep(s_axis_fifo_76_tkeep),
        .s_axis_fifo_76_tstrb(s_axis_fifo_76_tstrb),
        .s_axis_fifo_76_tdata(s_axis_fifo_76_tdata),
        .s_axis_fifo_76_tready(s_axis_fifo_76_tready),
        .ap_fifo_iarg_76_empty_n(ap_fifo_iarg_76_empty_n),
        .ap_fifo_iarg_76_dout(ap_fifo_iarg_76_dout),
        .ap_fifo_iarg_76_read(ap_fifo_iarg_76_read),
        .s_axis_fifo_77_aclk(s_axis_fifo_77_aclk),
        .s_axis_fifo_77_aresetn(s_axis_fifo_77_aresetn),
        .s_axis_fifo_77_tlast(s_axis_fifo_77_tlast),
        .s_axis_fifo_77_tvalid(s_axis_fifo_77_tvalid),
        .s_axis_fifo_77_tkeep(s_axis_fifo_77_tkeep),
        .s_axis_fifo_77_tstrb(s_axis_fifo_77_tstrb),
        .s_axis_fifo_77_tdata(s_axis_fifo_77_tdata),
        .s_axis_fifo_77_tready(s_axis_fifo_77_tready),
        .ap_fifo_iarg_77_empty_n(ap_fifo_iarg_77_empty_n),
        .ap_fifo_iarg_77_dout(ap_fifo_iarg_77_dout),
        .ap_fifo_iarg_77_read(ap_fifo_iarg_77_read),
        .s_axis_fifo_78_aclk(s_axis_fifo_78_aclk),
        .s_axis_fifo_78_aresetn(s_axis_fifo_78_aresetn),
        .s_axis_fifo_78_tlast(s_axis_fifo_78_tlast),
        .s_axis_fifo_78_tvalid(s_axis_fifo_78_tvalid),
        .s_axis_fifo_78_tkeep(s_axis_fifo_78_tkeep),
        .s_axis_fifo_78_tstrb(s_axis_fifo_78_tstrb),
        .s_axis_fifo_78_tdata(s_axis_fifo_78_tdata),
        .s_axis_fifo_78_tready(s_axis_fifo_78_tready),
        .ap_fifo_iarg_78_empty_n(ap_fifo_iarg_78_empty_n),
        .ap_fifo_iarg_78_dout(ap_fifo_iarg_78_dout),
        .ap_fifo_iarg_78_read(ap_fifo_iarg_78_read),
        .s_axis_fifo_79_aclk(s_axis_fifo_79_aclk),
        .s_axis_fifo_79_aresetn(s_axis_fifo_79_aresetn),
        .s_axis_fifo_79_tlast(s_axis_fifo_79_tlast),
        .s_axis_fifo_79_tvalid(s_axis_fifo_79_tvalid),
        .s_axis_fifo_79_tkeep(s_axis_fifo_79_tkeep),
        .s_axis_fifo_79_tstrb(s_axis_fifo_79_tstrb),
        .s_axis_fifo_79_tdata(s_axis_fifo_79_tdata),
        .s_axis_fifo_79_tready(s_axis_fifo_79_tready),
        .ap_fifo_iarg_79_empty_n(ap_fifo_iarg_79_empty_n),
        .ap_fifo_iarg_79_dout(ap_fifo_iarg_79_dout),
        .ap_fifo_iarg_79_read(ap_fifo_iarg_79_read),
        .s_axis_fifo_80_aclk(s_axis_fifo_80_aclk),
        .s_axis_fifo_80_aresetn(s_axis_fifo_80_aresetn),
        .s_axis_fifo_80_tlast(s_axis_fifo_80_tlast),
        .s_axis_fifo_80_tvalid(s_axis_fifo_80_tvalid),
        .s_axis_fifo_80_tkeep(s_axis_fifo_80_tkeep),
        .s_axis_fifo_80_tstrb(s_axis_fifo_80_tstrb),
        .s_axis_fifo_80_tdata(s_axis_fifo_80_tdata),
        .s_axis_fifo_80_tready(s_axis_fifo_80_tready),
        .ap_fifo_iarg_80_empty_n(ap_fifo_iarg_80_empty_n),
        .ap_fifo_iarg_80_dout(ap_fifo_iarg_80_dout),
        .ap_fifo_iarg_80_read(ap_fifo_iarg_80_read),
        .s_axis_fifo_81_aclk(s_axis_fifo_81_aclk),
        .s_axis_fifo_81_aresetn(s_axis_fifo_81_aresetn),
        .s_axis_fifo_81_tlast(s_axis_fifo_81_tlast),
        .s_axis_fifo_81_tvalid(s_axis_fifo_81_tvalid),
        .s_axis_fifo_81_tkeep(s_axis_fifo_81_tkeep),
        .s_axis_fifo_81_tstrb(s_axis_fifo_81_tstrb),
        .s_axis_fifo_81_tdata(s_axis_fifo_81_tdata),
        .s_axis_fifo_81_tready(s_axis_fifo_81_tready),
        .ap_fifo_iarg_81_empty_n(ap_fifo_iarg_81_empty_n),
        .ap_fifo_iarg_81_dout(ap_fifo_iarg_81_dout),
        .ap_fifo_iarg_81_read(ap_fifo_iarg_81_read),
        .s_axis_fifo_82_aclk(s_axis_fifo_82_aclk),
        .s_axis_fifo_82_aresetn(s_axis_fifo_82_aresetn),
        .s_axis_fifo_82_tlast(s_axis_fifo_82_tlast),
        .s_axis_fifo_82_tvalid(s_axis_fifo_82_tvalid),
        .s_axis_fifo_82_tkeep(s_axis_fifo_82_tkeep),
        .s_axis_fifo_82_tstrb(s_axis_fifo_82_tstrb),
        .s_axis_fifo_82_tdata(s_axis_fifo_82_tdata),
        .s_axis_fifo_82_tready(s_axis_fifo_82_tready),
        .ap_fifo_iarg_82_empty_n(ap_fifo_iarg_82_empty_n),
        .ap_fifo_iarg_82_dout(ap_fifo_iarg_82_dout),
        .ap_fifo_iarg_82_read(ap_fifo_iarg_82_read),
        .s_axis_fifo_83_aclk(s_axis_fifo_83_aclk),
        .s_axis_fifo_83_aresetn(s_axis_fifo_83_aresetn),
        .s_axis_fifo_83_tlast(s_axis_fifo_83_tlast),
        .s_axis_fifo_83_tvalid(s_axis_fifo_83_tvalid),
        .s_axis_fifo_83_tkeep(s_axis_fifo_83_tkeep),
        .s_axis_fifo_83_tstrb(s_axis_fifo_83_tstrb),
        .s_axis_fifo_83_tdata(s_axis_fifo_83_tdata),
        .s_axis_fifo_83_tready(s_axis_fifo_83_tready),
        .ap_fifo_iarg_83_empty_n(ap_fifo_iarg_83_empty_n),
        .ap_fifo_iarg_83_dout(ap_fifo_iarg_83_dout),
        .ap_fifo_iarg_83_read(ap_fifo_iarg_83_read),
        .s_axis_fifo_84_aclk(s_axis_fifo_84_aclk),
        .s_axis_fifo_84_aresetn(s_axis_fifo_84_aresetn),
        .s_axis_fifo_84_tlast(s_axis_fifo_84_tlast),
        .s_axis_fifo_84_tvalid(s_axis_fifo_84_tvalid),
        .s_axis_fifo_84_tkeep(s_axis_fifo_84_tkeep),
        .s_axis_fifo_84_tstrb(s_axis_fifo_84_tstrb),
        .s_axis_fifo_84_tdata(s_axis_fifo_84_tdata),
        .s_axis_fifo_84_tready(s_axis_fifo_84_tready),
        .ap_fifo_iarg_84_empty_n(ap_fifo_iarg_84_empty_n),
        .ap_fifo_iarg_84_dout(ap_fifo_iarg_84_dout),
        .ap_fifo_iarg_84_read(ap_fifo_iarg_84_read),
        .s_axis_fifo_85_aclk(s_axis_fifo_85_aclk),
        .s_axis_fifo_85_aresetn(s_axis_fifo_85_aresetn),
        .s_axis_fifo_85_tlast(s_axis_fifo_85_tlast),
        .s_axis_fifo_85_tvalid(s_axis_fifo_85_tvalid),
        .s_axis_fifo_85_tkeep(s_axis_fifo_85_tkeep),
        .s_axis_fifo_85_tstrb(s_axis_fifo_85_tstrb),
        .s_axis_fifo_85_tdata(s_axis_fifo_85_tdata),
        .s_axis_fifo_85_tready(s_axis_fifo_85_tready),
        .ap_fifo_iarg_85_empty_n(ap_fifo_iarg_85_empty_n),
        .ap_fifo_iarg_85_dout(ap_fifo_iarg_85_dout),
        .ap_fifo_iarg_85_read(ap_fifo_iarg_85_read),
        .s_axis_fifo_86_aclk(s_axis_fifo_86_aclk),
        .s_axis_fifo_86_aresetn(s_axis_fifo_86_aresetn),
        .s_axis_fifo_86_tlast(s_axis_fifo_86_tlast),
        .s_axis_fifo_86_tvalid(s_axis_fifo_86_tvalid),
        .s_axis_fifo_86_tkeep(s_axis_fifo_86_tkeep),
        .s_axis_fifo_86_tstrb(s_axis_fifo_86_tstrb),
        .s_axis_fifo_86_tdata(s_axis_fifo_86_tdata),
        .s_axis_fifo_86_tready(s_axis_fifo_86_tready),
        .ap_fifo_iarg_86_empty_n(ap_fifo_iarg_86_empty_n),
        .ap_fifo_iarg_86_dout(ap_fifo_iarg_86_dout),
        .ap_fifo_iarg_86_read(ap_fifo_iarg_86_read),
        .s_axis_fifo_87_aclk(s_axis_fifo_87_aclk),
        .s_axis_fifo_87_aresetn(s_axis_fifo_87_aresetn),
        .s_axis_fifo_87_tlast(s_axis_fifo_87_tlast),
        .s_axis_fifo_87_tvalid(s_axis_fifo_87_tvalid),
        .s_axis_fifo_87_tkeep(s_axis_fifo_87_tkeep),
        .s_axis_fifo_87_tstrb(s_axis_fifo_87_tstrb),
        .s_axis_fifo_87_tdata(s_axis_fifo_87_tdata),
        .s_axis_fifo_87_tready(s_axis_fifo_87_tready),
        .ap_fifo_iarg_87_empty_n(ap_fifo_iarg_87_empty_n),
        .ap_fifo_iarg_87_dout(ap_fifo_iarg_87_dout),
        .ap_fifo_iarg_87_read(ap_fifo_iarg_87_read),
        .s_axis_fifo_88_aclk(s_axis_fifo_88_aclk),
        .s_axis_fifo_88_aresetn(s_axis_fifo_88_aresetn),
        .s_axis_fifo_88_tlast(s_axis_fifo_88_tlast),
        .s_axis_fifo_88_tvalid(s_axis_fifo_88_tvalid),
        .s_axis_fifo_88_tkeep(s_axis_fifo_88_tkeep),
        .s_axis_fifo_88_tstrb(s_axis_fifo_88_tstrb),
        .s_axis_fifo_88_tdata(s_axis_fifo_88_tdata),
        .s_axis_fifo_88_tready(s_axis_fifo_88_tready),
        .ap_fifo_iarg_88_empty_n(ap_fifo_iarg_88_empty_n),
        .ap_fifo_iarg_88_dout(ap_fifo_iarg_88_dout),
        .ap_fifo_iarg_88_read(ap_fifo_iarg_88_read),
        .s_axis_fifo_89_aclk(s_axis_fifo_89_aclk),
        .s_axis_fifo_89_aresetn(s_axis_fifo_89_aresetn),
        .s_axis_fifo_89_tlast(s_axis_fifo_89_tlast),
        .s_axis_fifo_89_tvalid(s_axis_fifo_89_tvalid),
        .s_axis_fifo_89_tkeep(s_axis_fifo_89_tkeep),
        .s_axis_fifo_89_tstrb(s_axis_fifo_89_tstrb),
        .s_axis_fifo_89_tdata(s_axis_fifo_89_tdata),
        .s_axis_fifo_89_tready(s_axis_fifo_89_tready),
        .ap_fifo_iarg_89_empty_n(ap_fifo_iarg_89_empty_n),
        .ap_fifo_iarg_89_dout(ap_fifo_iarg_89_dout),
        .ap_fifo_iarg_89_read(ap_fifo_iarg_89_read),
        .s_axis_fifo_90_aclk(s_axis_fifo_90_aclk),
        .s_axis_fifo_90_aresetn(s_axis_fifo_90_aresetn),
        .s_axis_fifo_90_tlast(s_axis_fifo_90_tlast),
        .s_axis_fifo_90_tvalid(s_axis_fifo_90_tvalid),
        .s_axis_fifo_90_tkeep(s_axis_fifo_90_tkeep),
        .s_axis_fifo_90_tstrb(s_axis_fifo_90_tstrb),
        .s_axis_fifo_90_tdata(s_axis_fifo_90_tdata),
        .s_axis_fifo_90_tready(s_axis_fifo_90_tready),
        .ap_fifo_iarg_90_empty_n(ap_fifo_iarg_90_empty_n),
        .ap_fifo_iarg_90_dout(ap_fifo_iarg_90_dout),
        .ap_fifo_iarg_90_read(ap_fifo_iarg_90_read),
        .s_axis_fifo_91_aclk(s_axis_fifo_91_aclk),
        .s_axis_fifo_91_aresetn(s_axis_fifo_91_aresetn),
        .s_axis_fifo_91_tlast(s_axis_fifo_91_tlast),
        .s_axis_fifo_91_tvalid(s_axis_fifo_91_tvalid),
        .s_axis_fifo_91_tkeep(s_axis_fifo_91_tkeep),
        .s_axis_fifo_91_tstrb(s_axis_fifo_91_tstrb),
        .s_axis_fifo_91_tdata(s_axis_fifo_91_tdata),
        .s_axis_fifo_91_tready(s_axis_fifo_91_tready),
        .ap_fifo_iarg_91_empty_n(ap_fifo_iarg_91_empty_n),
        .ap_fifo_iarg_91_dout(ap_fifo_iarg_91_dout),
        .ap_fifo_iarg_91_read(ap_fifo_iarg_91_read),
        .s_axis_fifo_92_aclk(s_axis_fifo_92_aclk),
        .s_axis_fifo_92_aresetn(s_axis_fifo_92_aresetn),
        .s_axis_fifo_92_tlast(s_axis_fifo_92_tlast),
        .s_axis_fifo_92_tvalid(s_axis_fifo_92_tvalid),
        .s_axis_fifo_92_tkeep(s_axis_fifo_92_tkeep),
        .s_axis_fifo_92_tstrb(s_axis_fifo_92_tstrb),
        .s_axis_fifo_92_tdata(s_axis_fifo_92_tdata),
        .s_axis_fifo_92_tready(s_axis_fifo_92_tready),
        .ap_fifo_iarg_92_empty_n(ap_fifo_iarg_92_empty_n),
        .ap_fifo_iarg_92_dout(ap_fifo_iarg_92_dout),
        .ap_fifo_iarg_92_read(ap_fifo_iarg_92_read),
        .s_axis_fifo_93_aclk(s_axis_fifo_93_aclk),
        .s_axis_fifo_93_aresetn(s_axis_fifo_93_aresetn),
        .s_axis_fifo_93_tlast(s_axis_fifo_93_tlast),
        .s_axis_fifo_93_tvalid(s_axis_fifo_93_tvalid),
        .s_axis_fifo_93_tkeep(s_axis_fifo_93_tkeep),
        .s_axis_fifo_93_tstrb(s_axis_fifo_93_tstrb),
        .s_axis_fifo_93_tdata(s_axis_fifo_93_tdata),
        .s_axis_fifo_93_tready(s_axis_fifo_93_tready),
        .ap_fifo_iarg_93_empty_n(ap_fifo_iarg_93_empty_n),
        .ap_fifo_iarg_93_dout(ap_fifo_iarg_93_dout),
        .ap_fifo_iarg_93_read(ap_fifo_iarg_93_read),
        .s_axis_fifo_94_aclk(s_axis_fifo_94_aclk),
        .s_axis_fifo_94_aresetn(s_axis_fifo_94_aresetn),
        .s_axis_fifo_94_tlast(s_axis_fifo_94_tlast),
        .s_axis_fifo_94_tvalid(s_axis_fifo_94_tvalid),
        .s_axis_fifo_94_tkeep(s_axis_fifo_94_tkeep),
        .s_axis_fifo_94_tstrb(s_axis_fifo_94_tstrb),
        .s_axis_fifo_94_tdata(s_axis_fifo_94_tdata),
        .s_axis_fifo_94_tready(s_axis_fifo_94_tready),
        .ap_fifo_iarg_94_empty_n(ap_fifo_iarg_94_empty_n),
        .ap_fifo_iarg_94_dout(ap_fifo_iarg_94_dout),
        .ap_fifo_iarg_94_read(ap_fifo_iarg_94_read),
        .s_axis_fifo_95_aclk(s_axis_fifo_95_aclk),
        .s_axis_fifo_95_aresetn(s_axis_fifo_95_aresetn),
        .s_axis_fifo_95_tlast(s_axis_fifo_95_tlast),
        .s_axis_fifo_95_tvalid(s_axis_fifo_95_tvalid),
        .s_axis_fifo_95_tkeep(s_axis_fifo_95_tkeep),
        .s_axis_fifo_95_tstrb(s_axis_fifo_95_tstrb),
        .s_axis_fifo_95_tdata(s_axis_fifo_95_tdata),
        .s_axis_fifo_95_tready(s_axis_fifo_95_tready),
        .ap_fifo_iarg_95_empty_n(ap_fifo_iarg_95_empty_n),
        .ap_fifo_iarg_95_dout(ap_fifo_iarg_95_dout),
        .ap_fifo_iarg_95_read(ap_fifo_iarg_95_read),
        .s_axis_fifo_96_aclk(s_axis_fifo_96_aclk),
        .s_axis_fifo_96_aresetn(s_axis_fifo_96_aresetn),
        .s_axis_fifo_96_tlast(s_axis_fifo_96_tlast),
        .s_axis_fifo_96_tvalid(s_axis_fifo_96_tvalid),
        .s_axis_fifo_96_tkeep(s_axis_fifo_96_tkeep),
        .s_axis_fifo_96_tstrb(s_axis_fifo_96_tstrb),
        .s_axis_fifo_96_tdata(s_axis_fifo_96_tdata),
        .s_axis_fifo_96_tready(s_axis_fifo_96_tready),
        .ap_fifo_iarg_96_empty_n(ap_fifo_iarg_96_empty_n),
        .ap_fifo_iarg_96_dout(ap_fifo_iarg_96_dout),
        .ap_fifo_iarg_96_read(ap_fifo_iarg_96_read),
        .s_axis_fifo_97_aclk(s_axis_fifo_97_aclk),
        .s_axis_fifo_97_aresetn(s_axis_fifo_97_aresetn),
        .s_axis_fifo_97_tlast(s_axis_fifo_97_tlast),
        .s_axis_fifo_97_tvalid(s_axis_fifo_97_tvalid),
        .s_axis_fifo_97_tkeep(s_axis_fifo_97_tkeep),
        .s_axis_fifo_97_tstrb(s_axis_fifo_97_tstrb),
        .s_axis_fifo_97_tdata(s_axis_fifo_97_tdata),
        .s_axis_fifo_97_tready(s_axis_fifo_97_tready),
        .ap_fifo_iarg_97_empty_n(ap_fifo_iarg_97_empty_n),
        .ap_fifo_iarg_97_dout(ap_fifo_iarg_97_dout),
        .ap_fifo_iarg_97_read(ap_fifo_iarg_97_read),
        .s_axis_fifo_98_aclk(s_axis_fifo_98_aclk),
        .s_axis_fifo_98_aresetn(s_axis_fifo_98_aresetn),
        .s_axis_fifo_98_tlast(s_axis_fifo_98_tlast),
        .s_axis_fifo_98_tvalid(s_axis_fifo_98_tvalid),
        .s_axis_fifo_98_tkeep(s_axis_fifo_98_tkeep),
        .s_axis_fifo_98_tstrb(s_axis_fifo_98_tstrb),
        .s_axis_fifo_98_tdata(s_axis_fifo_98_tdata),
        .s_axis_fifo_98_tready(s_axis_fifo_98_tready),
        .ap_fifo_iarg_98_empty_n(ap_fifo_iarg_98_empty_n),
        .ap_fifo_iarg_98_dout(ap_fifo_iarg_98_dout),
        .ap_fifo_iarg_98_read(ap_fifo_iarg_98_read),
        .s_axis_fifo_99_aclk(s_axis_fifo_99_aclk),
        .s_axis_fifo_99_aresetn(s_axis_fifo_99_aresetn),
        .s_axis_fifo_99_tlast(s_axis_fifo_99_tlast),
        .s_axis_fifo_99_tvalid(s_axis_fifo_99_tvalid),
        .s_axis_fifo_99_tkeep(s_axis_fifo_99_tkeep),
        .s_axis_fifo_99_tstrb(s_axis_fifo_99_tstrb),
        .s_axis_fifo_99_tdata(s_axis_fifo_99_tdata),
        .s_axis_fifo_99_tready(s_axis_fifo_99_tready),
        .ap_fifo_iarg_99_empty_n(ap_fifo_iarg_99_empty_n),
        .ap_fifo_iarg_99_dout(ap_fifo_iarg_99_dout),
        .ap_fifo_iarg_99_read(ap_fifo_iarg_99_read),
        .s_axis_fifo_100_aclk(s_axis_fifo_100_aclk),
        .s_axis_fifo_100_aresetn(s_axis_fifo_100_aresetn),
        .s_axis_fifo_100_tlast(s_axis_fifo_100_tlast),
        .s_axis_fifo_100_tvalid(s_axis_fifo_100_tvalid),
        .s_axis_fifo_100_tkeep(s_axis_fifo_100_tkeep),
        .s_axis_fifo_100_tstrb(s_axis_fifo_100_tstrb),
        .s_axis_fifo_100_tdata(s_axis_fifo_100_tdata),
        .s_axis_fifo_100_tready(s_axis_fifo_100_tready),
        .ap_fifo_iarg_100_empty_n(ap_fifo_iarg_100_empty_n),
        .ap_fifo_iarg_100_dout(ap_fifo_iarg_100_dout),
        .ap_fifo_iarg_100_read(ap_fifo_iarg_100_read),
        .s_axis_fifo_101_aclk(s_axis_fifo_101_aclk),
        .s_axis_fifo_101_aresetn(s_axis_fifo_101_aresetn),
        .s_axis_fifo_101_tlast(s_axis_fifo_101_tlast),
        .s_axis_fifo_101_tvalid(s_axis_fifo_101_tvalid),
        .s_axis_fifo_101_tkeep(s_axis_fifo_101_tkeep),
        .s_axis_fifo_101_tstrb(s_axis_fifo_101_tstrb),
        .s_axis_fifo_101_tdata(s_axis_fifo_101_tdata),
        .s_axis_fifo_101_tready(s_axis_fifo_101_tready),
        .ap_fifo_iarg_101_empty_n(ap_fifo_iarg_101_empty_n),
        .ap_fifo_iarg_101_dout(ap_fifo_iarg_101_dout),
        .ap_fifo_iarg_101_read(ap_fifo_iarg_101_read),
        .s_axis_fifo_102_aclk(s_axis_fifo_102_aclk),
        .s_axis_fifo_102_aresetn(s_axis_fifo_102_aresetn),
        .s_axis_fifo_102_tlast(s_axis_fifo_102_tlast),
        .s_axis_fifo_102_tvalid(s_axis_fifo_102_tvalid),
        .s_axis_fifo_102_tkeep(s_axis_fifo_102_tkeep),
        .s_axis_fifo_102_tstrb(s_axis_fifo_102_tstrb),
        .s_axis_fifo_102_tdata(s_axis_fifo_102_tdata),
        .s_axis_fifo_102_tready(s_axis_fifo_102_tready),
        .ap_fifo_iarg_102_empty_n(ap_fifo_iarg_102_empty_n),
        .ap_fifo_iarg_102_dout(ap_fifo_iarg_102_dout),
        .ap_fifo_iarg_102_read(ap_fifo_iarg_102_read),
        .s_axis_fifo_103_aclk(s_axis_fifo_103_aclk),
        .s_axis_fifo_103_aresetn(s_axis_fifo_103_aresetn),
        .s_axis_fifo_103_tlast(s_axis_fifo_103_tlast),
        .s_axis_fifo_103_tvalid(s_axis_fifo_103_tvalid),
        .s_axis_fifo_103_tkeep(s_axis_fifo_103_tkeep),
        .s_axis_fifo_103_tstrb(s_axis_fifo_103_tstrb),
        .s_axis_fifo_103_tdata(s_axis_fifo_103_tdata),
        .s_axis_fifo_103_tready(s_axis_fifo_103_tready),
        .ap_fifo_iarg_103_empty_n(ap_fifo_iarg_103_empty_n),
        .ap_fifo_iarg_103_dout(ap_fifo_iarg_103_dout),
        .ap_fifo_iarg_103_read(ap_fifo_iarg_103_read),
        .s_axis_fifo_104_aclk(s_axis_fifo_104_aclk),
        .s_axis_fifo_104_aresetn(s_axis_fifo_104_aresetn),
        .s_axis_fifo_104_tlast(s_axis_fifo_104_tlast),
        .s_axis_fifo_104_tvalid(s_axis_fifo_104_tvalid),
        .s_axis_fifo_104_tkeep(s_axis_fifo_104_tkeep),
        .s_axis_fifo_104_tstrb(s_axis_fifo_104_tstrb),
        .s_axis_fifo_104_tdata(s_axis_fifo_104_tdata),
        .s_axis_fifo_104_tready(s_axis_fifo_104_tready),
        .ap_fifo_iarg_104_empty_n(ap_fifo_iarg_104_empty_n),
        .ap_fifo_iarg_104_dout(ap_fifo_iarg_104_dout),
        .ap_fifo_iarg_104_read(ap_fifo_iarg_104_read),
        .s_axis_fifo_105_aclk(s_axis_fifo_105_aclk),
        .s_axis_fifo_105_aresetn(s_axis_fifo_105_aresetn),
        .s_axis_fifo_105_tlast(s_axis_fifo_105_tlast),
        .s_axis_fifo_105_tvalid(s_axis_fifo_105_tvalid),
        .s_axis_fifo_105_tkeep(s_axis_fifo_105_tkeep),
        .s_axis_fifo_105_tstrb(s_axis_fifo_105_tstrb),
        .s_axis_fifo_105_tdata(s_axis_fifo_105_tdata),
        .s_axis_fifo_105_tready(s_axis_fifo_105_tready),
        .ap_fifo_iarg_105_empty_n(ap_fifo_iarg_105_empty_n),
        .ap_fifo_iarg_105_dout(ap_fifo_iarg_105_dout),
        .ap_fifo_iarg_105_read(ap_fifo_iarg_105_read),
        .s_axis_fifo_106_aclk(s_axis_fifo_106_aclk),
        .s_axis_fifo_106_aresetn(s_axis_fifo_106_aresetn),
        .s_axis_fifo_106_tlast(s_axis_fifo_106_tlast),
        .s_axis_fifo_106_tvalid(s_axis_fifo_106_tvalid),
        .s_axis_fifo_106_tkeep(s_axis_fifo_106_tkeep),
        .s_axis_fifo_106_tstrb(s_axis_fifo_106_tstrb),
        .s_axis_fifo_106_tdata(s_axis_fifo_106_tdata),
        .s_axis_fifo_106_tready(s_axis_fifo_106_tready),
        .ap_fifo_iarg_106_empty_n(ap_fifo_iarg_106_empty_n),
        .ap_fifo_iarg_106_dout(ap_fifo_iarg_106_dout),
        .ap_fifo_iarg_106_read(ap_fifo_iarg_106_read),
        .s_axis_fifo_107_aclk(s_axis_fifo_107_aclk),
        .s_axis_fifo_107_aresetn(s_axis_fifo_107_aresetn),
        .s_axis_fifo_107_tlast(s_axis_fifo_107_tlast),
        .s_axis_fifo_107_tvalid(s_axis_fifo_107_tvalid),
        .s_axis_fifo_107_tkeep(s_axis_fifo_107_tkeep),
        .s_axis_fifo_107_tstrb(s_axis_fifo_107_tstrb),
        .s_axis_fifo_107_tdata(s_axis_fifo_107_tdata),
        .s_axis_fifo_107_tready(s_axis_fifo_107_tready),
        .ap_fifo_iarg_107_empty_n(ap_fifo_iarg_107_empty_n),
        .ap_fifo_iarg_107_dout(ap_fifo_iarg_107_dout),
        .ap_fifo_iarg_107_read(ap_fifo_iarg_107_read),
        .s_axis_fifo_108_aclk(s_axis_fifo_108_aclk),
        .s_axis_fifo_108_aresetn(s_axis_fifo_108_aresetn),
        .s_axis_fifo_108_tlast(s_axis_fifo_108_tlast),
        .s_axis_fifo_108_tvalid(s_axis_fifo_108_tvalid),
        .s_axis_fifo_108_tkeep(s_axis_fifo_108_tkeep),
        .s_axis_fifo_108_tstrb(s_axis_fifo_108_tstrb),
        .s_axis_fifo_108_tdata(s_axis_fifo_108_tdata),
        .s_axis_fifo_108_tready(s_axis_fifo_108_tready),
        .ap_fifo_iarg_108_empty_n(ap_fifo_iarg_108_empty_n),
        .ap_fifo_iarg_108_dout(ap_fifo_iarg_108_dout),
        .ap_fifo_iarg_108_read(ap_fifo_iarg_108_read),
        .s_axis_fifo_109_aclk(s_axis_fifo_109_aclk),
        .s_axis_fifo_109_aresetn(s_axis_fifo_109_aresetn),
        .s_axis_fifo_109_tlast(s_axis_fifo_109_tlast),
        .s_axis_fifo_109_tvalid(s_axis_fifo_109_tvalid),
        .s_axis_fifo_109_tkeep(s_axis_fifo_109_tkeep),
        .s_axis_fifo_109_tstrb(s_axis_fifo_109_tstrb),
        .s_axis_fifo_109_tdata(s_axis_fifo_109_tdata),
        .s_axis_fifo_109_tready(s_axis_fifo_109_tready),
        .ap_fifo_iarg_109_empty_n(ap_fifo_iarg_109_empty_n),
        .ap_fifo_iarg_109_dout(ap_fifo_iarg_109_dout),
        .ap_fifo_iarg_109_read(ap_fifo_iarg_109_read),
        .s_axis_fifo_110_aclk(s_axis_fifo_110_aclk),
        .s_axis_fifo_110_aresetn(s_axis_fifo_110_aresetn),
        .s_axis_fifo_110_tlast(s_axis_fifo_110_tlast),
        .s_axis_fifo_110_tvalid(s_axis_fifo_110_tvalid),
        .s_axis_fifo_110_tkeep(s_axis_fifo_110_tkeep),
        .s_axis_fifo_110_tstrb(s_axis_fifo_110_tstrb),
        .s_axis_fifo_110_tdata(s_axis_fifo_110_tdata),
        .s_axis_fifo_110_tready(s_axis_fifo_110_tready),
        .ap_fifo_iarg_110_empty_n(ap_fifo_iarg_110_empty_n),
        .ap_fifo_iarg_110_dout(ap_fifo_iarg_110_dout),
        .ap_fifo_iarg_110_read(ap_fifo_iarg_110_read),
        .s_axis_fifo_111_aclk(s_axis_fifo_111_aclk),
        .s_axis_fifo_111_aresetn(s_axis_fifo_111_aresetn),
        .s_axis_fifo_111_tlast(s_axis_fifo_111_tlast),
        .s_axis_fifo_111_tvalid(s_axis_fifo_111_tvalid),
        .s_axis_fifo_111_tkeep(s_axis_fifo_111_tkeep),
        .s_axis_fifo_111_tstrb(s_axis_fifo_111_tstrb),
        .s_axis_fifo_111_tdata(s_axis_fifo_111_tdata),
        .s_axis_fifo_111_tready(s_axis_fifo_111_tready),
        .ap_fifo_iarg_111_empty_n(ap_fifo_iarg_111_empty_n),
        .ap_fifo_iarg_111_dout(ap_fifo_iarg_111_dout),
        .ap_fifo_iarg_111_read(ap_fifo_iarg_111_read),
        .s_axis_fifo_112_aclk(s_axis_fifo_112_aclk),
        .s_axis_fifo_112_aresetn(s_axis_fifo_112_aresetn),
        .s_axis_fifo_112_tlast(s_axis_fifo_112_tlast),
        .s_axis_fifo_112_tvalid(s_axis_fifo_112_tvalid),
        .s_axis_fifo_112_tkeep(s_axis_fifo_112_tkeep),
        .s_axis_fifo_112_tstrb(s_axis_fifo_112_tstrb),
        .s_axis_fifo_112_tdata(s_axis_fifo_112_tdata),
        .s_axis_fifo_112_tready(s_axis_fifo_112_tready),
        .ap_fifo_iarg_112_empty_n(ap_fifo_iarg_112_empty_n),
        .ap_fifo_iarg_112_dout(ap_fifo_iarg_112_dout),
        .ap_fifo_iarg_112_read(ap_fifo_iarg_112_read),
        .s_axis_fifo_113_aclk(s_axis_fifo_113_aclk),
        .s_axis_fifo_113_aresetn(s_axis_fifo_113_aresetn),
        .s_axis_fifo_113_tlast(s_axis_fifo_113_tlast),
        .s_axis_fifo_113_tvalid(s_axis_fifo_113_tvalid),
        .s_axis_fifo_113_tkeep(s_axis_fifo_113_tkeep),
        .s_axis_fifo_113_tstrb(s_axis_fifo_113_tstrb),
        .s_axis_fifo_113_tdata(s_axis_fifo_113_tdata),
        .s_axis_fifo_113_tready(s_axis_fifo_113_tready),
        .ap_fifo_iarg_113_empty_n(ap_fifo_iarg_113_empty_n),
        .ap_fifo_iarg_113_dout(ap_fifo_iarg_113_dout),
        .ap_fifo_iarg_113_read(ap_fifo_iarg_113_read),
        .s_axis_fifo_114_aclk(s_axis_fifo_114_aclk),
        .s_axis_fifo_114_aresetn(s_axis_fifo_114_aresetn),
        .s_axis_fifo_114_tlast(s_axis_fifo_114_tlast),
        .s_axis_fifo_114_tvalid(s_axis_fifo_114_tvalid),
        .s_axis_fifo_114_tkeep(s_axis_fifo_114_tkeep),
        .s_axis_fifo_114_tstrb(s_axis_fifo_114_tstrb),
        .s_axis_fifo_114_tdata(s_axis_fifo_114_tdata),
        .s_axis_fifo_114_tready(s_axis_fifo_114_tready),
        .ap_fifo_iarg_114_empty_n(ap_fifo_iarg_114_empty_n),
        .ap_fifo_iarg_114_dout(ap_fifo_iarg_114_dout),
        .ap_fifo_iarg_114_read(ap_fifo_iarg_114_read),
        .s_axis_fifo_115_aclk(s_axis_fifo_115_aclk),
        .s_axis_fifo_115_aresetn(s_axis_fifo_115_aresetn),
        .s_axis_fifo_115_tlast(s_axis_fifo_115_tlast),
        .s_axis_fifo_115_tvalid(s_axis_fifo_115_tvalid),
        .s_axis_fifo_115_tkeep(s_axis_fifo_115_tkeep),
        .s_axis_fifo_115_tstrb(s_axis_fifo_115_tstrb),
        .s_axis_fifo_115_tdata(s_axis_fifo_115_tdata),
        .s_axis_fifo_115_tready(s_axis_fifo_115_tready),
        .ap_fifo_iarg_115_empty_n(ap_fifo_iarg_115_empty_n),
        .ap_fifo_iarg_115_dout(ap_fifo_iarg_115_dout),
        .ap_fifo_iarg_115_read(ap_fifo_iarg_115_read),
        .s_axis_fifo_116_aclk(s_axis_fifo_116_aclk),
        .s_axis_fifo_116_aresetn(s_axis_fifo_116_aresetn),
        .s_axis_fifo_116_tlast(s_axis_fifo_116_tlast),
        .s_axis_fifo_116_tvalid(s_axis_fifo_116_tvalid),
        .s_axis_fifo_116_tkeep(s_axis_fifo_116_tkeep),
        .s_axis_fifo_116_tstrb(s_axis_fifo_116_tstrb),
        .s_axis_fifo_116_tdata(s_axis_fifo_116_tdata),
        .s_axis_fifo_116_tready(s_axis_fifo_116_tready),
        .ap_fifo_iarg_116_empty_n(ap_fifo_iarg_116_empty_n),
        .ap_fifo_iarg_116_dout(ap_fifo_iarg_116_dout),
        .ap_fifo_iarg_116_read(ap_fifo_iarg_116_read),
        .s_axis_fifo_117_aclk(s_axis_fifo_117_aclk),
        .s_axis_fifo_117_aresetn(s_axis_fifo_117_aresetn),
        .s_axis_fifo_117_tlast(s_axis_fifo_117_tlast),
        .s_axis_fifo_117_tvalid(s_axis_fifo_117_tvalid),
        .s_axis_fifo_117_tkeep(s_axis_fifo_117_tkeep),
        .s_axis_fifo_117_tstrb(s_axis_fifo_117_tstrb),
        .s_axis_fifo_117_tdata(s_axis_fifo_117_tdata),
        .s_axis_fifo_117_tready(s_axis_fifo_117_tready),
        .ap_fifo_iarg_117_empty_n(ap_fifo_iarg_117_empty_n),
        .ap_fifo_iarg_117_dout(ap_fifo_iarg_117_dout),
        .ap_fifo_iarg_117_read(ap_fifo_iarg_117_read),
        .s_axis_fifo_118_aclk(s_axis_fifo_118_aclk),
        .s_axis_fifo_118_aresetn(s_axis_fifo_118_aresetn),
        .s_axis_fifo_118_tlast(s_axis_fifo_118_tlast),
        .s_axis_fifo_118_tvalid(s_axis_fifo_118_tvalid),
        .s_axis_fifo_118_tkeep(s_axis_fifo_118_tkeep),
        .s_axis_fifo_118_tstrb(s_axis_fifo_118_tstrb),
        .s_axis_fifo_118_tdata(s_axis_fifo_118_tdata),
        .s_axis_fifo_118_tready(s_axis_fifo_118_tready),
        .ap_fifo_iarg_118_empty_n(ap_fifo_iarg_118_empty_n),
        .ap_fifo_iarg_118_dout(ap_fifo_iarg_118_dout),
        .ap_fifo_iarg_118_read(ap_fifo_iarg_118_read),
        .s_axis_fifo_119_aclk(s_axis_fifo_119_aclk),
        .s_axis_fifo_119_aresetn(s_axis_fifo_119_aresetn),
        .s_axis_fifo_119_tlast(s_axis_fifo_119_tlast),
        .s_axis_fifo_119_tvalid(s_axis_fifo_119_tvalid),
        .s_axis_fifo_119_tkeep(s_axis_fifo_119_tkeep),
        .s_axis_fifo_119_tstrb(s_axis_fifo_119_tstrb),
        .s_axis_fifo_119_tdata(s_axis_fifo_119_tdata),
        .s_axis_fifo_119_tready(s_axis_fifo_119_tready),
        .ap_fifo_iarg_119_empty_n(ap_fifo_iarg_119_empty_n),
        .ap_fifo_iarg_119_dout(ap_fifo_iarg_119_dout),
        .ap_fifo_iarg_119_read(ap_fifo_iarg_119_read),
        .s_axis_fifo_120_aclk(s_axis_fifo_120_aclk),
        .s_axis_fifo_120_aresetn(s_axis_fifo_120_aresetn),
        .s_axis_fifo_120_tlast(s_axis_fifo_120_tlast),
        .s_axis_fifo_120_tvalid(s_axis_fifo_120_tvalid),
        .s_axis_fifo_120_tkeep(s_axis_fifo_120_tkeep),
        .s_axis_fifo_120_tstrb(s_axis_fifo_120_tstrb),
        .s_axis_fifo_120_tdata(s_axis_fifo_120_tdata),
        .s_axis_fifo_120_tready(s_axis_fifo_120_tready),
        .ap_fifo_iarg_120_empty_n(ap_fifo_iarg_120_empty_n),
        .ap_fifo_iarg_120_dout(ap_fifo_iarg_120_dout),
        .ap_fifo_iarg_120_read(ap_fifo_iarg_120_read),
        .s_axis_fifo_121_aclk(s_axis_fifo_121_aclk),
        .s_axis_fifo_121_aresetn(s_axis_fifo_121_aresetn),
        .s_axis_fifo_121_tlast(s_axis_fifo_121_tlast),
        .s_axis_fifo_121_tvalid(s_axis_fifo_121_tvalid),
        .s_axis_fifo_121_tkeep(s_axis_fifo_121_tkeep),
        .s_axis_fifo_121_tstrb(s_axis_fifo_121_tstrb),
        .s_axis_fifo_121_tdata(s_axis_fifo_121_tdata),
        .s_axis_fifo_121_tready(s_axis_fifo_121_tready),
        .ap_fifo_iarg_121_empty_n(ap_fifo_iarg_121_empty_n),
        .ap_fifo_iarg_121_dout(ap_fifo_iarg_121_dout),
        .ap_fifo_iarg_121_read(ap_fifo_iarg_121_read),
        .s_axis_fifo_122_aclk(s_axis_fifo_122_aclk),
        .s_axis_fifo_122_aresetn(s_axis_fifo_122_aresetn),
        .s_axis_fifo_122_tlast(s_axis_fifo_122_tlast),
        .s_axis_fifo_122_tvalid(s_axis_fifo_122_tvalid),
        .s_axis_fifo_122_tkeep(s_axis_fifo_122_tkeep),
        .s_axis_fifo_122_tstrb(s_axis_fifo_122_tstrb),
        .s_axis_fifo_122_tdata(s_axis_fifo_122_tdata),
        .s_axis_fifo_122_tready(s_axis_fifo_122_tready),
        .ap_fifo_iarg_122_empty_n(ap_fifo_iarg_122_empty_n),
        .ap_fifo_iarg_122_dout(ap_fifo_iarg_122_dout),
        .ap_fifo_iarg_122_read(ap_fifo_iarg_122_read),
        .s_axis_fifo_123_aclk(s_axis_fifo_123_aclk),
        .s_axis_fifo_123_aresetn(s_axis_fifo_123_aresetn),
        .s_axis_fifo_123_tlast(s_axis_fifo_123_tlast),
        .s_axis_fifo_123_tvalid(s_axis_fifo_123_tvalid),
        .s_axis_fifo_123_tkeep(s_axis_fifo_123_tkeep),
        .s_axis_fifo_123_tstrb(s_axis_fifo_123_tstrb),
        .s_axis_fifo_123_tdata(s_axis_fifo_123_tdata),
        .s_axis_fifo_123_tready(s_axis_fifo_123_tready),
        .ap_fifo_iarg_123_empty_n(ap_fifo_iarg_123_empty_n),
        .ap_fifo_iarg_123_dout(ap_fifo_iarg_123_dout),
        .ap_fifo_iarg_123_read(ap_fifo_iarg_123_read),
        .s_axis_fifo_124_aclk(s_axis_fifo_124_aclk),
        .s_axis_fifo_124_aresetn(s_axis_fifo_124_aresetn),
        .s_axis_fifo_124_tlast(s_axis_fifo_124_tlast),
        .s_axis_fifo_124_tvalid(s_axis_fifo_124_tvalid),
        .s_axis_fifo_124_tkeep(s_axis_fifo_124_tkeep),
        .s_axis_fifo_124_tstrb(s_axis_fifo_124_tstrb),
        .s_axis_fifo_124_tdata(s_axis_fifo_124_tdata),
        .s_axis_fifo_124_tready(s_axis_fifo_124_tready),
        .ap_fifo_iarg_124_empty_n(ap_fifo_iarg_124_empty_n),
        .ap_fifo_iarg_124_dout(ap_fifo_iarg_124_dout),
        .ap_fifo_iarg_124_read(ap_fifo_iarg_124_read),
        .s_axis_fifo_125_aclk(s_axis_fifo_125_aclk),
        .s_axis_fifo_125_aresetn(s_axis_fifo_125_aresetn),
        .s_axis_fifo_125_tlast(s_axis_fifo_125_tlast),
        .s_axis_fifo_125_tvalid(s_axis_fifo_125_tvalid),
        .s_axis_fifo_125_tkeep(s_axis_fifo_125_tkeep),
        .s_axis_fifo_125_tstrb(s_axis_fifo_125_tstrb),
        .s_axis_fifo_125_tdata(s_axis_fifo_125_tdata),
        .s_axis_fifo_125_tready(s_axis_fifo_125_tready),
        .ap_fifo_iarg_125_empty_n(ap_fifo_iarg_125_empty_n),
        .ap_fifo_iarg_125_dout(ap_fifo_iarg_125_dout),
        .ap_fifo_iarg_125_read(ap_fifo_iarg_125_read),
        .s_axis_fifo_126_aclk(s_axis_fifo_126_aclk),
        .s_axis_fifo_126_aresetn(s_axis_fifo_126_aresetn),
        .s_axis_fifo_126_tlast(s_axis_fifo_126_tlast),
        .s_axis_fifo_126_tvalid(s_axis_fifo_126_tvalid),
        .s_axis_fifo_126_tkeep(s_axis_fifo_126_tkeep),
        .s_axis_fifo_126_tstrb(s_axis_fifo_126_tstrb),
        .s_axis_fifo_126_tdata(s_axis_fifo_126_tdata),
        .s_axis_fifo_126_tready(s_axis_fifo_126_tready),
        .ap_fifo_iarg_126_empty_n(ap_fifo_iarg_126_empty_n),
        .ap_fifo_iarg_126_dout(ap_fifo_iarg_126_dout),
        .ap_fifo_iarg_126_read(ap_fifo_iarg_126_read),
        .s_axis_fifo_127_aclk(s_axis_fifo_127_aclk),
        .s_axis_fifo_127_aresetn(s_axis_fifo_127_aresetn),
        .s_axis_fifo_127_tlast(s_axis_fifo_127_tlast),
        .s_axis_fifo_127_tvalid(s_axis_fifo_127_tvalid),
        .s_axis_fifo_127_tkeep(s_axis_fifo_127_tkeep),
        .s_axis_fifo_127_tstrb(s_axis_fifo_127_tstrb),
        .s_axis_fifo_127_tdata(s_axis_fifo_127_tdata),
        .s_axis_fifo_127_tready(s_axis_fifo_127_tready),
        .ap_fifo_iarg_127_empty_n(ap_fifo_iarg_127_empty_n),
        .ap_fifo_iarg_127_dout(ap_fifo_iarg_127_dout),
        .ap_fifo_iarg_127_read(ap_fifo_iarg_127_read)
    );
        
    out_fifo_args #(
        .C_NUM_OUTPUT_FIFOs(C_NUM_OUTPUT_FIFOs),
        .M_AXIS_FIFO_0_WIDTH(M_AXIS_FIFO_0_WIDTH),
        .M_AXIS_FIFO_1_WIDTH(M_AXIS_FIFO_1_WIDTH),
        .M_AXIS_FIFO_2_WIDTH(M_AXIS_FIFO_2_WIDTH),
        .M_AXIS_FIFO_3_WIDTH(M_AXIS_FIFO_3_WIDTH),
        .M_AXIS_FIFO_4_WIDTH(M_AXIS_FIFO_4_WIDTH),
        .M_AXIS_FIFO_5_WIDTH(M_AXIS_FIFO_5_WIDTH),
        .M_AXIS_FIFO_6_WIDTH(M_AXIS_FIFO_6_WIDTH),
        .M_AXIS_FIFO_7_WIDTH(M_AXIS_FIFO_7_WIDTH),
        .M_AXIS_FIFO_8_WIDTH(M_AXIS_FIFO_8_WIDTH),
        .M_AXIS_FIFO_9_WIDTH(M_AXIS_FIFO_9_WIDTH),
        .M_AXIS_FIFO_10_WIDTH(M_AXIS_FIFO_10_WIDTH),
        .M_AXIS_FIFO_11_WIDTH(M_AXIS_FIFO_11_WIDTH),
        .M_AXIS_FIFO_12_WIDTH(M_AXIS_FIFO_12_WIDTH),
        .M_AXIS_FIFO_13_WIDTH(M_AXIS_FIFO_13_WIDTH),
        .M_AXIS_FIFO_14_WIDTH(M_AXIS_FIFO_14_WIDTH),
        .M_AXIS_FIFO_15_WIDTH(M_AXIS_FIFO_15_WIDTH),
        .M_AXIS_FIFO_16_WIDTH(M_AXIS_FIFO_16_WIDTH),
        .M_AXIS_FIFO_17_WIDTH(M_AXIS_FIFO_17_WIDTH),
        .M_AXIS_FIFO_18_WIDTH(M_AXIS_FIFO_18_WIDTH),
        .M_AXIS_FIFO_19_WIDTH(M_AXIS_FIFO_19_WIDTH),
        .M_AXIS_FIFO_20_WIDTH(M_AXIS_FIFO_20_WIDTH),
        .M_AXIS_FIFO_21_WIDTH(M_AXIS_FIFO_21_WIDTH),
        .M_AXIS_FIFO_22_WIDTH(M_AXIS_FIFO_22_WIDTH),
        .M_AXIS_FIFO_23_WIDTH(M_AXIS_FIFO_23_WIDTH),
        .M_AXIS_FIFO_24_WIDTH(M_AXIS_FIFO_24_WIDTH),
        .M_AXIS_FIFO_25_WIDTH(M_AXIS_FIFO_25_WIDTH),
        .M_AXIS_FIFO_26_WIDTH(M_AXIS_FIFO_26_WIDTH),
        .M_AXIS_FIFO_27_WIDTH(M_AXIS_FIFO_27_WIDTH),
        .M_AXIS_FIFO_28_WIDTH(M_AXIS_FIFO_28_WIDTH),
        .M_AXIS_FIFO_29_WIDTH(M_AXIS_FIFO_29_WIDTH),
        .M_AXIS_FIFO_30_WIDTH(M_AXIS_FIFO_30_WIDTH),
        .M_AXIS_FIFO_31_WIDTH(M_AXIS_FIFO_31_WIDTH),
        .M_AXIS_FIFO_32_WIDTH(M_AXIS_FIFO_32_WIDTH),
        .M_AXIS_FIFO_33_WIDTH(M_AXIS_FIFO_33_WIDTH),
        .M_AXIS_FIFO_34_WIDTH(M_AXIS_FIFO_34_WIDTH),
        .M_AXIS_FIFO_35_WIDTH(M_AXIS_FIFO_35_WIDTH),
        .M_AXIS_FIFO_36_WIDTH(M_AXIS_FIFO_36_WIDTH),
        .M_AXIS_FIFO_37_WIDTH(M_AXIS_FIFO_37_WIDTH),
        .M_AXIS_FIFO_38_WIDTH(M_AXIS_FIFO_38_WIDTH),
        .M_AXIS_FIFO_39_WIDTH(M_AXIS_FIFO_39_WIDTH),
        .M_AXIS_FIFO_40_WIDTH(M_AXIS_FIFO_40_WIDTH),
        .M_AXIS_FIFO_41_WIDTH(M_AXIS_FIFO_41_WIDTH),
        .M_AXIS_FIFO_42_WIDTH(M_AXIS_FIFO_42_WIDTH),
        .M_AXIS_FIFO_43_WIDTH(M_AXIS_FIFO_43_WIDTH),
        .M_AXIS_FIFO_44_WIDTH(M_AXIS_FIFO_44_WIDTH),
        .M_AXIS_FIFO_45_WIDTH(M_AXIS_FIFO_45_WIDTH),
        .M_AXIS_FIFO_46_WIDTH(M_AXIS_FIFO_46_WIDTH),
        .M_AXIS_FIFO_47_WIDTH(M_AXIS_FIFO_47_WIDTH),
        .M_AXIS_FIFO_48_WIDTH(M_AXIS_FIFO_48_WIDTH),
        .M_AXIS_FIFO_49_WIDTH(M_AXIS_FIFO_49_WIDTH),
        .M_AXIS_FIFO_50_WIDTH(M_AXIS_FIFO_50_WIDTH),
        .M_AXIS_FIFO_51_WIDTH(M_AXIS_FIFO_51_WIDTH),
        .M_AXIS_FIFO_52_WIDTH(M_AXIS_FIFO_52_WIDTH),
        .M_AXIS_FIFO_53_WIDTH(M_AXIS_FIFO_53_WIDTH),
        .M_AXIS_FIFO_54_WIDTH(M_AXIS_FIFO_54_WIDTH),
        .M_AXIS_FIFO_55_WIDTH(M_AXIS_FIFO_55_WIDTH),
        .M_AXIS_FIFO_56_WIDTH(M_AXIS_FIFO_56_WIDTH),
        .M_AXIS_FIFO_57_WIDTH(M_AXIS_FIFO_57_WIDTH),
        .M_AXIS_FIFO_58_WIDTH(M_AXIS_FIFO_58_WIDTH),
        .M_AXIS_FIFO_59_WIDTH(M_AXIS_FIFO_59_WIDTH),
        .M_AXIS_FIFO_60_WIDTH(M_AXIS_FIFO_60_WIDTH),
        .M_AXIS_FIFO_61_WIDTH(M_AXIS_FIFO_61_WIDTH),
        .M_AXIS_FIFO_62_WIDTH(M_AXIS_FIFO_62_WIDTH),
        .M_AXIS_FIFO_63_WIDTH(M_AXIS_FIFO_63_WIDTH),
        .M_AXIS_FIFO_64_WIDTH(M_AXIS_FIFO_64_WIDTH),
        .M_AXIS_FIFO_65_WIDTH(M_AXIS_FIFO_65_WIDTH),
        .M_AXIS_FIFO_66_WIDTH(M_AXIS_FIFO_66_WIDTH),
        .M_AXIS_FIFO_67_WIDTH(M_AXIS_FIFO_67_WIDTH),
        .M_AXIS_FIFO_68_WIDTH(M_AXIS_FIFO_68_WIDTH),
        .M_AXIS_FIFO_69_WIDTH(M_AXIS_FIFO_69_WIDTH),
        .M_AXIS_FIFO_70_WIDTH(M_AXIS_FIFO_70_WIDTH),
        .M_AXIS_FIFO_71_WIDTH(M_AXIS_FIFO_71_WIDTH),
        .M_AXIS_FIFO_72_WIDTH(M_AXIS_FIFO_72_WIDTH),
        .M_AXIS_FIFO_73_WIDTH(M_AXIS_FIFO_73_WIDTH),
        .M_AXIS_FIFO_74_WIDTH(M_AXIS_FIFO_74_WIDTH),
        .M_AXIS_FIFO_75_WIDTH(M_AXIS_FIFO_75_WIDTH),
        .M_AXIS_FIFO_76_WIDTH(M_AXIS_FIFO_76_WIDTH),
        .M_AXIS_FIFO_77_WIDTH(M_AXIS_FIFO_77_WIDTH),
        .M_AXIS_FIFO_78_WIDTH(M_AXIS_FIFO_78_WIDTH),
        .M_AXIS_FIFO_79_WIDTH(M_AXIS_FIFO_79_WIDTH),
        .M_AXIS_FIFO_80_WIDTH(M_AXIS_FIFO_80_WIDTH),
        .M_AXIS_FIFO_81_WIDTH(M_AXIS_FIFO_81_WIDTH),
        .M_AXIS_FIFO_82_WIDTH(M_AXIS_FIFO_82_WIDTH),
        .M_AXIS_FIFO_83_WIDTH(M_AXIS_FIFO_83_WIDTH),
        .M_AXIS_FIFO_84_WIDTH(M_AXIS_FIFO_84_WIDTH),
        .M_AXIS_FIFO_85_WIDTH(M_AXIS_FIFO_85_WIDTH),
        .M_AXIS_FIFO_86_WIDTH(M_AXIS_FIFO_86_WIDTH),
        .M_AXIS_FIFO_87_WIDTH(M_AXIS_FIFO_87_WIDTH),
        .M_AXIS_FIFO_88_WIDTH(M_AXIS_FIFO_88_WIDTH),
        .M_AXIS_FIFO_89_WIDTH(M_AXIS_FIFO_89_WIDTH),
        .M_AXIS_FIFO_90_WIDTH(M_AXIS_FIFO_90_WIDTH),
        .M_AXIS_FIFO_91_WIDTH(M_AXIS_FIFO_91_WIDTH),
        .M_AXIS_FIFO_92_WIDTH(M_AXIS_FIFO_92_WIDTH),
        .M_AXIS_FIFO_93_WIDTH(M_AXIS_FIFO_93_WIDTH),
        .M_AXIS_FIFO_94_WIDTH(M_AXIS_FIFO_94_WIDTH),
        .M_AXIS_FIFO_95_WIDTH(M_AXIS_FIFO_95_WIDTH),
        .M_AXIS_FIFO_96_WIDTH(M_AXIS_FIFO_96_WIDTH),
        .M_AXIS_FIFO_97_WIDTH(M_AXIS_FIFO_97_WIDTH),
        .M_AXIS_FIFO_98_WIDTH(M_AXIS_FIFO_98_WIDTH),
        .M_AXIS_FIFO_99_WIDTH(M_AXIS_FIFO_99_WIDTH),
        .M_AXIS_FIFO_100_WIDTH(M_AXIS_FIFO_100_WIDTH),
        .M_AXIS_FIFO_101_WIDTH(M_AXIS_FIFO_101_WIDTH),
        .M_AXIS_FIFO_102_WIDTH(M_AXIS_FIFO_102_WIDTH),
        .M_AXIS_FIFO_103_WIDTH(M_AXIS_FIFO_103_WIDTH),
        .M_AXIS_FIFO_104_WIDTH(M_AXIS_FIFO_104_WIDTH),
        .M_AXIS_FIFO_105_WIDTH(M_AXIS_FIFO_105_WIDTH),
        .M_AXIS_FIFO_106_WIDTH(M_AXIS_FIFO_106_WIDTH),
        .M_AXIS_FIFO_107_WIDTH(M_AXIS_FIFO_107_WIDTH),
        .M_AXIS_FIFO_108_WIDTH(M_AXIS_FIFO_108_WIDTH),
        .M_AXIS_FIFO_109_WIDTH(M_AXIS_FIFO_109_WIDTH),
        .M_AXIS_FIFO_110_WIDTH(M_AXIS_FIFO_110_WIDTH),
        .M_AXIS_FIFO_111_WIDTH(M_AXIS_FIFO_111_WIDTH),
        .M_AXIS_FIFO_112_WIDTH(M_AXIS_FIFO_112_WIDTH),
        .M_AXIS_FIFO_113_WIDTH(M_AXIS_FIFO_113_WIDTH),
        .M_AXIS_FIFO_114_WIDTH(M_AXIS_FIFO_114_WIDTH),
        .M_AXIS_FIFO_115_WIDTH(M_AXIS_FIFO_115_WIDTH),
        .M_AXIS_FIFO_116_WIDTH(M_AXIS_FIFO_116_WIDTH),
        .M_AXIS_FIFO_117_WIDTH(M_AXIS_FIFO_117_WIDTH),
        .M_AXIS_FIFO_118_WIDTH(M_AXIS_FIFO_118_WIDTH),
        .M_AXIS_FIFO_119_WIDTH(M_AXIS_FIFO_119_WIDTH),
        .M_AXIS_FIFO_120_WIDTH(M_AXIS_FIFO_120_WIDTH),
        .M_AXIS_FIFO_121_WIDTH(M_AXIS_FIFO_121_WIDTH),
        .M_AXIS_FIFO_122_WIDTH(M_AXIS_FIFO_122_WIDTH),
        .M_AXIS_FIFO_123_WIDTH(M_AXIS_FIFO_123_WIDTH),
        .M_AXIS_FIFO_124_WIDTH(M_AXIS_FIFO_124_WIDTH),
        .M_AXIS_FIFO_125_WIDTH(M_AXIS_FIFO_125_WIDTH),
        .M_AXIS_FIFO_126_WIDTH(M_AXIS_FIFO_126_WIDTH),
        .M_AXIS_FIFO_127_WIDTH(M_AXIS_FIFO_127_WIDTH),
        .M_AXIS_FIFO_0_DEPTH(M_AXIS_FIFO_0_DEPTH),
        .M_AXIS_FIFO_1_DEPTH(M_AXIS_FIFO_1_DEPTH),
        .M_AXIS_FIFO_2_DEPTH(M_AXIS_FIFO_2_DEPTH),
        .M_AXIS_FIFO_3_DEPTH(M_AXIS_FIFO_3_DEPTH),
        .M_AXIS_FIFO_4_DEPTH(M_AXIS_FIFO_4_DEPTH),
        .M_AXIS_FIFO_5_DEPTH(M_AXIS_FIFO_5_DEPTH),
        .M_AXIS_FIFO_6_DEPTH(M_AXIS_FIFO_6_DEPTH),
        .M_AXIS_FIFO_7_DEPTH(M_AXIS_FIFO_7_DEPTH),
        .M_AXIS_FIFO_8_DEPTH(M_AXIS_FIFO_8_DEPTH),
        .M_AXIS_FIFO_9_DEPTH(M_AXIS_FIFO_9_DEPTH),
        .M_AXIS_FIFO_10_DEPTH(M_AXIS_FIFO_10_DEPTH),
        .M_AXIS_FIFO_11_DEPTH(M_AXIS_FIFO_11_DEPTH),
        .M_AXIS_FIFO_12_DEPTH(M_AXIS_FIFO_12_DEPTH),
        .M_AXIS_FIFO_13_DEPTH(M_AXIS_FIFO_13_DEPTH),
        .M_AXIS_FIFO_14_DEPTH(M_AXIS_FIFO_14_DEPTH),
        .M_AXIS_FIFO_15_DEPTH(M_AXIS_FIFO_15_DEPTH),
        .M_AXIS_FIFO_16_DEPTH(M_AXIS_FIFO_16_DEPTH),
        .M_AXIS_FIFO_17_DEPTH(M_AXIS_FIFO_17_DEPTH),
        .M_AXIS_FIFO_18_DEPTH(M_AXIS_FIFO_18_DEPTH),
        .M_AXIS_FIFO_19_DEPTH(M_AXIS_FIFO_19_DEPTH),
        .M_AXIS_FIFO_20_DEPTH(M_AXIS_FIFO_20_DEPTH),
        .M_AXIS_FIFO_21_DEPTH(M_AXIS_FIFO_21_DEPTH),
        .M_AXIS_FIFO_22_DEPTH(M_AXIS_FIFO_22_DEPTH),
        .M_AXIS_FIFO_23_DEPTH(M_AXIS_FIFO_23_DEPTH),
        .M_AXIS_FIFO_24_DEPTH(M_AXIS_FIFO_24_DEPTH),
        .M_AXIS_FIFO_25_DEPTH(M_AXIS_FIFO_25_DEPTH),
        .M_AXIS_FIFO_26_DEPTH(M_AXIS_FIFO_26_DEPTH),
        .M_AXIS_FIFO_27_DEPTH(M_AXIS_FIFO_27_DEPTH),
        .M_AXIS_FIFO_28_DEPTH(M_AXIS_FIFO_28_DEPTH),
        .M_AXIS_FIFO_29_DEPTH(M_AXIS_FIFO_29_DEPTH),
        .M_AXIS_FIFO_30_DEPTH(M_AXIS_FIFO_30_DEPTH),
        .M_AXIS_FIFO_31_DEPTH(M_AXIS_FIFO_31_DEPTH),
        .M_AXIS_FIFO_32_DEPTH(M_AXIS_FIFO_32_DEPTH),
        .M_AXIS_FIFO_33_DEPTH(M_AXIS_FIFO_33_DEPTH),
        .M_AXIS_FIFO_34_DEPTH(M_AXIS_FIFO_34_DEPTH),
        .M_AXIS_FIFO_35_DEPTH(M_AXIS_FIFO_35_DEPTH),
        .M_AXIS_FIFO_36_DEPTH(M_AXIS_FIFO_36_DEPTH),
        .M_AXIS_FIFO_37_DEPTH(M_AXIS_FIFO_37_DEPTH),
        .M_AXIS_FIFO_38_DEPTH(M_AXIS_FIFO_38_DEPTH),
        .M_AXIS_FIFO_39_DEPTH(M_AXIS_FIFO_39_DEPTH),
        .M_AXIS_FIFO_40_DEPTH(M_AXIS_FIFO_40_DEPTH),
        .M_AXIS_FIFO_41_DEPTH(M_AXIS_FIFO_41_DEPTH),
        .M_AXIS_FIFO_42_DEPTH(M_AXIS_FIFO_42_DEPTH),
        .M_AXIS_FIFO_43_DEPTH(M_AXIS_FIFO_43_DEPTH),
        .M_AXIS_FIFO_44_DEPTH(M_AXIS_FIFO_44_DEPTH),
        .M_AXIS_FIFO_45_DEPTH(M_AXIS_FIFO_45_DEPTH),
        .M_AXIS_FIFO_46_DEPTH(M_AXIS_FIFO_46_DEPTH),
        .M_AXIS_FIFO_47_DEPTH(M_AXIS_FIFO_47_DEPTH),
        .M_AXIS_FIFO_48_DEPTH(M_AXIS_FIFO_48_DEPTH),
        .M_AXIS_FIFO_49_DEPTH(M_AXIS_FIFO_49_DEPTH),
        .M_AXIS_FIFO_50_DEPTH(M_AXIS_FIFO_50_DEPTH),
        .M_AXIS_FIFO_51_DEPTH(M_AXIS_FIFO_51_DEPTH),
        .M_AXIS_FIFO_52_DEPTH(M_AXIS_FIFO_52_DEPTH),
        .M_AXIS_FIFO_53_DEPTH(M_AXIS_FIFO_53_DEPTH),
        .M_AXIS_FIFO_54_DEPTH(M_AXIS_FIFO_54_DEPTH),
        .M_AXIS_FIFO_55_DEPTH(M_AXIS_FIFO_55_DEPTH),
        .M_AXIS_FIFO_56_DEPTH(M_AXIS_FIFO_56_DEPTH),
        .M_AXIS_FIFO_57_DEPTH(M_AXIS_FIFO_57_DEPTH),
        .M_AXIS_FIFO_58_DEPTH(M_AXIS_FIFO_58_DEPTH),
        .M_AXIS_FIFO_59_DEPTH(M_AXIS_FIFO_59_DEPTH),
        .M_AXIS_FIFO_60_DEPTH(M_AXIS_FIFO_60_DEPTH),
        .M_AXIS_FIFO_61_DEPTH(M_AXIS_FIFO_61_DEPTH),
        .M_AXIS_FIFO_62_DEPTH(M_AXIS_FIFO_62_DEPTH),
        .M_AXIS_FIFO_63_DEPTH(M_AXIS_FIFO_63_DEPTH),
        .M_AXIS_FIFO_64_DEPTH(M_AXIS_FIFO_64_DEPTH),
        .M_AXIS_FIFO_65_DEPTH(M_AXIS_FIFO_65_DEPTH),
        .M_AXIS_FIFO_66_DEPTH(M_AXIS_FIFO_66_DEPTH),
        .M_AXIS_FIFO_67_DEPTH(M_AXIS_FIFO_67_DEPTH),
        .M_AXIS_FIFO_68_DEPTH(M_AXIS_FIFO_68_DEPTH),
        .M_AXIS_FIFO_69_DEPTH(M_AXIS_FIFO_69_DEPTH),
        .M_AXIS_FIFO_70_DEPTH(M_AXIS_FIFO_70_DEPTH),
        .M_AXIS_FIFO_71_DEPTH(M_AXIS_FIFO_71_DEPTH),
        .M_AXIS_FIFO_72_DEPTH(M_AXIS_FIFO_72_DEPTH),
        .M_AXIS_FIFO_73_DEPTH(M_AXIS_FIFO_73_DEPTH),
        .M_AXIS_FIFO_74_DEPTH(M_AXIS_FIFO_74_DEPTH),
        .M_AXIS_FIFO_75_DEPTH(M_AXIS_FIFO_75_DEPTH),
        .M_AXIS_FIFO_76_DEPTH(M_AXIS_FIFO_76_DEPTH),
        .M_AXIS_FIFO_77_DEPTH(M_AXIS_FIFO_77_DEPTH),
        .M_AXIS_FIFO_78_DEPTH(M_AXIS_FIFO_78_DEPTH),
        .M_AXIS_FIFO_79_DEPTH(M_AXIS_FIFO_79_DEPTH),
        .M_AXIS_FIFO_80_DEPTH(M_AXIS_FIFO_80_DEPTH),
        .M_AXIS_FIFO_81_DEPTH(M_AXIS_FIFO_81_DEPTH),
        .M_AXIS_FIFO_82_DEPTH(M_AXIS_FIFO_82_DEPTH),
        .M_AXIS_FIFO_83_DEPTH(M_AXIS_FIFO_83_DEPTH),
        .M_AXIS_FIFO_84_DEPTH(M_AXIS_FIFO_84_DEPTH),
        .M_AXIS_FIFO_85_DEPTH(M_AXIS_FIFO_85_DEPTH),
        .M_AXIS_FIFO_86_DEPTH(M_AXIS_FIFO_86_DEPTH),
        .M_AXIS_FIFO_87_DEPTH(M_AXIS_FIFO_87_DEPTH),
        .M_AXIS_FIFO_88_DEPTH(M_AXIS_FIFO_88_DEPTH),
        .M_AXIS_FIFO_89_DEPTH(M_AXIS_FIFO_89_DEPTH),
        .M_AXIS_FIFO_90_DEPTH(M_AXIS_FIFO_90_DEPTH),
        .M_AXIS_FIFO_91_DEPTH(M_AXIS_FIFO_91_DEPTH),
        .M_AXIS_FIFO_92_DEPTH(M_AXIS_FIFO_92_DEPTH),
        .M_AXIS_FIFO_93_DEPTH(M_AXIS_FIFO_93_DEPTH),
        .M_AXIS_FIFO_94_DEPTH(M_AXIS_FIFO_94_DEPTH),
        .M_AXIS_FIFO_95_DEPTH(M_AXIS_FIFO_95_DEPTH),
        .M_AXIS_FIFO_96_DEPTH(M_AXIS_FIFO_96_DEPTH),
        .M_AXIS_FIFO_97_DEPTH(M_AXIS_FIFO_97_DEPTH),
        .M_AXIS_FIFO_98_DEPTH(M_AXIS_FIFO_98_DEPTH),
        .M_AXIS_FIFO_99_DEPTH(M_AXIS_FIFO_99_DEPTH),
        .M_AXIS_FIFO_100_DEPTH(M_AXIS_FIFO_100_DEPTH),
        .M_AXIS_FIFO_101_DEPTH(M_AXIS_FIFO_101_DEPTH),
        .M_AXIS_FIFO_102_DEPTH(M_AXIS_FIFO_102_DEPTH),
        .M_AXIS_FIFO_103_DEPTH(M_AXIS_FIFO_103_DEPTH),
        .M_AXIS_FIFO_104_DEPTH(M_AXIS_FIFO_104_DEPTH),
        .M_AXIS_FIFO_105_DEPTH(M_AXIS_FIFO_105_DEPTH),
        .M_AXIS_FIFO_106_DEPTH(M_AXIS_FIFO_106_DEPTH),
        .M_AXIS_FIFO_107_DEPTH(M_AXIS_FIFO_107_DEPTH),
        .M_AXIS_FIFO_108_DEPTH(M_AXIS_FIFO_108_DEPTH),
        .M_AXIS_FIFO_109_DEPTH(M_AXIS_FIFO_109_DEPTH),
        .M_AXIS_FIFO_110_DEPTH(M_AXIS_FIFO_110_DEPTH),
        .M_AXIS_FIFO_111_DEPTH(M_AXIS_FIFO_111_DEPTH),
        .M_AXIS_FIFO_112_DEPTH(M_AXIS_FIFO_112_DEPTH),
        .M_AXIS_FIFO_113_DEPTH(M_AXIS_FIFO_113_DEPTH),
        .M_AXIS_FIFO_114_DEPTH(M_AXIS_FIFO_114_DEPTH),
        .M_AXIS_FIFO_115_DEPTH(M_AXIS_FIFO_115_DEPTH),
        .M_AXIS_FIFO_116_DEPTH(M_AXIS_FIFO_116_DEPTH),
        .M_AXIS_FIFO_117_DEPTH(M_AXIS_FIFO_117_DEPTH),
        .M_AXIS_FIFO_118_DEPTH(M_AXIS_FIFO_118_DEPTH),
        .M_AXIS_FIFO_119_DEPTH(M_AXIS_FIFO_119_DEPTH),
        .M_AXIS_FIFO_120_DEPTH(M_AXIS_FIFO_120_DEPTH),
        .M_AXIS_FIFO_121_DEPTH(M_AXIS_FIFO_121_DEPTH),
        .M_AXIS_FIFO_122_DEPTH(M_AXIS_FIFO_122_DEPTH),
        .M_AXIS_FIFO_123_DEPTH(M_AXIS_FIFO_123_DEPTH),
        .M_AXIS_FIFO_124_DEPTH(M_AXIS_FIFO_124_DEPTH),
        .M_AXIS_FIFO_125_DEPTH(M_AXIS_FIFO_125_DEPTH),
        .M_AXIS_FIFO_126_DEPTH(M_AXIS_FIFO_126_DEPTH),
        .M_AXIS_FIFO_127_DEPTH(M_AXIS_FIFO_127_DEPTH),
        .M_AXIS_FIFO_0_IS_ASYNC(M_AXIS_FIFO_0_IS_ASYNC),
        .M_AXIS_FIFO_1_IS_ASYNC(M_AXIS_FIFO_1_IS_ASYNC),
        .M_AXIS_FIFO_2_IS_ASYNC(M_AXIS_FIFO_2_IS_ASYNC),
        .M_AXIS_FIFO_3_IS_ASYNC(M_AXIS_FIFO_3_IS_ASYNC),
        .M_AXIS_FIFO_4_IS_ASYNC(M_AXIS_FIFO_4_IS_ASYNC),
        .M_AXIS_FIFO_5_IS_ASYNC(M_AXIS_FIFO_5_IS_ASYNC),
        .M_AXIS_FIFO_6_IS_ASYNC(M_AXIS_FIFO_6_IS_ASYNC),
        .M_AXIS_FIFO_7_IS_ASYNC(M_AXIS_FIFO_7_IS_ASYNC),
        .M_AXIS_FIFO_8_IS_ASYNC(M_AXIS_FIFO_8_IS_ASYNC),
        .M_AXIS_FIFO_9_IS_ASYNC(M_AXIS_FIFO_9_IS_ASYNC),
        .M_AXIS_FIFO_10_IS_ASYNC(M_AXIS_FIFO_10_IS_ASYNC),
        .M_AXIS_FIFO_11_IS_ASYNC(M_AXIS_FIFO_11_IS_ASYNC),
        .M_AXIS_FIFO_12_IS_ASYNC(M_AXIS_FIFO_12_IS_ASYNC),
        .M_AXIS_FIFO_13_IS_ASYNC(M_AXIS_FIFO_13_IS_ASYNC),
        .M_AXIS_FIFO_14_IS_ASYNC(M_AXIS_FIFO_14_IS_ASYNC),
        .M_AXIS_FIFO_15_IS_ASYNC(M_AXIS_FIFO_15_IS_ASYNC),
        .M_AXIS_FIFO_16_IS_ASYNC(M_AXIS_FIFO_16_IS_ASYNC),
        .M_AXIS_FIFO_17_IS_ASYNC(M_AXIS_FIFO_17_IS_ASYNC),
        .M_AXIS_FIFO_18_IS_ASYNC(M_AXIS_FIFO_18_IS_ASYNC),
        .M_AXIS_FIFO_19_IS_ASYNC(M_AXIS_FIFO_19_IS_ASYNC),
        .M_AXIS_FIFO_20_IS_ASYNC(M_AXIS_FIFO_20_IS_ASYNC),
        .M_AXIS_FIFO_21_IS_ASYNC(M_AXIS_FIFO_21_IS_ASYNC),
        .M_AXIS_FIFO_22_IS_ASYNC(M_AXIS_FIFO_22_IS_ASYNC),
        .M_AXIS_FIFO_23_IS_ASYNC(M_AXIS_FIFO_23_IS_ASYNC),
        .M_AXIS_FIFO_24_IS_ASYNC(M_AXIS_FIFO_24_IS_ASYNC),
        .M_AXIS_FIFO_25_IS_ASYNC(M_AXIS_FIFO_25_IS_ASYNC),
        .M_AXIS_FIFO_26_IS_ASYNC(M_AXIS_FIFO_26_IS_ASYNC),
        .M_AXIS_FIFO_27_IS_ASYNC(M_AXIS_FIFO_27_IS_ASYNC),
        .M_AXIS_FIFO_28_IS_ASYNC(M_AXIS_FIFO_28_IS_ASYNC),
        .M_AXIS_FIFO_29_IS_ASYNC(M_AXIS_FIFO_29_IS_ASYNC),
        .M_AXIS_FIFO_30_IS_ASYNC(M_AXIS_FIFO_30_IS_ASYNC),
        .M_AXIS_FIFO_31_IS_ASYNC(M_AXIS_FIFO_31_IS_ASYNC),
        .M_AXIS_FIFO_32_IS_ASYNC(M_AXIS_FIFO_32_IS_ASYNC),
        .M_AXIS_FIFO_33_IS_ASYNC(M_AXIS_FIFO_33_IS_ASYNC),
        .M_AXIS_FIFO_34_IS_ASYNC(M_AXIS_FIFO_34_IS_ASYNC),
        .M_AXIS_FIFO_35_IS_ASYNC(M_AXIS_FIFO_35_IS_ASYNC),
        .M_AXIS_FIFO_36_IS_ASYNC(M_AXIS_FIFO_36_IS_ASYNC),
        .M_AXIS_FIFO_37_IS_ASYNC(M_AXIS_FIFO_37_IS_ASYNC),
        .M_AXIS_FIFO_38_IS_ASYNC(M_AXIS_FIFO_38_IS_ASYNC),
        .M_AXIS_FIFO_39_IS_ASYNC(M_AXIS_FIFO_39_IS_ASYNC),
        .M_AXIS_FIFO_40_IS_ASYNC(M_AXIS_FIFO_40_IS_ASYNC),
        .M_AXIS_FIFO_41_IS_ASYNC(M_AXIS_FIFO_41_IS_ASYNC),
        .M_AXIS_FIFO_42_IS_ASYNC(M_AXIS_FIFO_42_IS_ASYNC),
        .M_AXIS_FIFO_43_IS_ASYNC(M_AXIS_FIFO_43_IS_ASYNC),
        .M_AXIS_FIFO_44_IS_ASYNC(M_AXIS_FIFO_44_IS_ASYNC),
        .M_AXIS_FIFO_45_IS_ASYNC(M_AXIS_FIFO_45_IS_ASYNC),
        .M_AXIS_FIFO_46_IS_ASYNC(M_AXIS_FIFO_46_IS_ASYNC),
        .M_AXIS_FIFO_47_IS_ASYNC(M_AXIS_FIFO_47_IS_ASYNC),
        .M_AXIS_FIFO_48_IS_ASYNC(M_AXIS_FIFO_48_IS_ASYNC),
        .M_AXIS_FIFO_49_IS_ASYNC(M_AXIS_FIFO_49_IS_ASYNC),
        .M_AXIS_FIFO_50_IS_ASYNC(M_AXIS_FIFO_50_IS_ASYNC),
        .M_AXIS_FIFO_51_IS_ASYNC(M_AXIS_FIFO_51_IS_ASYNC),
        .M_AXIS_FIFO_52_IS_ASYNC(M_AXIS_FIFO_52_IS_ASYNC),
        .M_AXIS_FIFO_53_IS_ASYNC(M_AXIS_FIFO_53_IS_ASYNC),
        .M_AXIS_FIFO_54_IS_ASYNC(M_AXIS_FIFO_54_IS_ASYNC),
        .M_AXIS_FIFO_55_IS_ASYNC(M_AXIS_FIFO_55_IS_ASYNC),
        .M_AXIS_FIFO_56_IS_ASYNC(M_AXIS_FIFO_56_IS_ASYNC),
        .M_AXIS_FIFO_57_IS_ASYNC(M_AXIS_FIFO_57_IS_ASYNC),
        .M_AXIS_FIFO_58_IS_ASYNC(M_AXIS_FIFO_58_IS_ASYNC),
        .M_AXIS_FIFO_59_IS_ASYNC(M_AXIS_FIFO_59_IS_ASYNC),
        .M_AXIS_FIFO_60_IS_ASYNC(M_AXIS_FIFO_60_IS_ASYNC),
        .M_AXIS_FIFO_61_IS_ASYNC(M_AXIS_FIFO_61_IS_ASYNC),
        .M_AXIS_FIFO_62_IS_ASYNC(M_AXIS_FIFO_62_IS_ASYNC),
        .M_AXIS_FIFO_63_IS_ASYNC(M_AXIS_FIFO_63_IS_ASYNC),
        .M_AXIS_FIFO_64_IS_ASYNC(M_AXIS_FIFO_64_IS_ASYNC),
        .M_AXIS_FIFO_65_IS_ASYNC(M_AXIS_FIFO_65_IS_ASYNC),
        .M_AXIS_FIFO_66_IS_ASYNC(M_AXIS_FIFO_66_IS_ASYNC),
        .M_AXIS_FIFO_67_IS_ASYNC(M_AXIS_FIFO_67_IS_ASYNC),
        .M_AXIS_FIFO_68_IS_ASYNC(M_AXIS_FIFO_68_IS_ASYNC),
        .M_AXIS_FIFO_69_IS_ASYNC(M_AXIS_FIFO_69_IS_ASYNC),
        .M_AXIS_FIFO_70_IS_ASYNC(M_AXIS_FIFO_70_IS_ASYNC),
        .M_AXIS_FIFO_71_IS_ASYNC(M_AXIS_FIFO_71_IS_ASYNC),
        .M_AXIS_FIFO_72_IS_ASYNC(M_AXIS_FIFO_72_IS_ASYNC),
        .M_AXIS_FIFO_73_IS_ASYNC(M_AXIS_FIFO_73_IS_ASYNC),
        .M_AXIS_FIFO_74_IS_ASYNC(M_AXIS_FIFO_74_IS_ASYNC),
        .M_AXIS_FIFO_75_IS_ASYNC(M_AXIS_FIFO_75_IS_ASYNC),
        .M_AXIS_FIFO_76_IS_ASYNC(M_AXIS_FIFO_76_IS_ASYNC),
        .M_AXIS_FIFO_77_IS_ASYNC(M_AXIS_FIFO_77_IS_ASYNC),
        .M_AXIS_FIFO_78_IS_ASYNC(M_AXIS_FIFO_78_IS_ASYNC),
        .M_AXIS_FIFO_79_IS_ASYNC(M_AXIS_FIFO_79_IS_ASYNC),
        .M_AXIS_FIFO_80_IS_ASYNC(M_AXIS_FIFO_80_IS_ASYNC),
        .M_AXIS_FIFO_81_IS_ASYNC(M_AXIS_FIFO_81_IS_ASYNC),
        .M_AXIS_FIFO_82_IS_ASYNC(M_AXIS_FIFO_82_IS_ASYNC),
        .M_AXIS_FIFO_83_IS_ASYNC(M_AXIS_FIFO_83_IS_ASYNC),
        .M_AXIS_FIFO_84_IS_ASYNC(M_AXIS_FIFO_84_IS_ASYNC),
        .M_AXIS_FIFO_85_IS_ASYNC(M_AXIS_FIFO_85_IS_ASYNC),
        .M_AXIS_FIFO_86_IS_ASYNC(M_AXIS_FIFO_86_IS_ASYNC),
        .M_AXIS_FIFO_87_IS_ASYNC(M_AXIS_FIFO_87_IS_ASYNC),
        .M_AXIS_FIFO_88_IS_ASYNC(M_AXIS_FIFO_88_IS_ASYNC),
        .M_AXIS_FIFO_89_IS_ASYNC(M_AXIS_FIFO_89_IS_ASYNC),
        .M_AXIS_FIFO_90_IS_ASYNC(M_AXIS_FIFO_90_IS_ASYNC),
        .M_AXIS_FIFO_91_IS_ASYNC(M_AXIS_FIFO_91_IS_ASYNC),
        .M_AXIS_FIFO_92_IS_ASYNC(M_AXIS_FIFO_92_IS_ASYNC),
        .M_AXIS_FIFO_93_IS_ASYNC(M_AXIS_FIFO_93_IS_ASYNC),
        .M_AXIS_FIFO_94_IS_ASYNC(M_AXIS_FIFO_94_IS_ASYNC),
        .M_AXIS_FIFO_95_IS_ASYNC(M_AXIS_FIFO_95_IS_ASYNC),
        .M_AXIS_FIFO_96_IS_ASYNC(M_AXIS_FIFO_96_IS_ASYNC),
        .M_AXIS_FIFO_97_IS_ASYNC(M_AXIS_FIFO_97_IS_ASYNC),
        .M_AXIS_FIFO_98_IS_ASYNC(M_AXIS_FIFO_98_IS_ASYNC),
        .M_AXIS_FIFO_99_IS_ASYNC(M_AXIS_FIFO_99_IS_ASYNC),
        .M_AXIS_FIFO_100_IS_ASYNC(M_AXIS_FIFO_100_IS_ASYNC),
        .M_AXIS_FIFO_101_IS_ASYNC(M_AXIS_FIFO_101_IS_ASYNC),
        .M_AXIS_FIFO_102_IS_ASYNC(M_AXIS_FIFO_102_IS_ASYNC),
        .M_AXIS_FIFO_103_IS_ASYNC(M_AXIS_FIFO_103_IS_ASYNC),
        .M_AXIS_FIFO_104_IS_ASYNC(M_AXIS_FIFO_104_IS_ASYNC),
        .M_AXIS_FIFO_105_IS_ASYNC(M_AXIS_FIFO_105_IS_ASYNC),
        .M_AXIS_FIFO_106_IS_ASYNC(M_AXIS_FIFO_106_IS_ASYNC),
        .M_AXIS_FIFO_107_IS_ASYNC(M_AXIS_FIFO_107_IS_ASYNC),
        .M_AXIS_FIFO_108_IS_ASYNC(M_AXIS_FIFO_108_IS_ASYNC),
        .M_AXIS_FIFO_109_IS_ASYNC(M_AXIS_FIFO_109_IS_ASYNC),
        .M_AXIS_FIFO_110_IS_ASYNC(M_AXIS_FIFO_110_IS_ASYNC),
        .M_AXIS_FIFO_111_IS_ASYNC(M_AXIS_FIFO_111_IS_ASYNC),
        .M_AXIS_FIFO_112_IS_ASYNC(M_AXIS_FIFO_112_IS_ASYNC),
        .M_AXIS_FIFO_113_IS_ASYNC(M_AXIS_FIFO_113_IS_ASYNC),
        .M_AXIS_FIFO_114_IS_ASYNC(M_AXIS_FIFO_114_IS_ASYNC),
        .M_AXIS_FIFO_115_IS_ASYNC(M_AXIS_FIFO_115_IS_ASYNC),
        .M_AXIS_FIFO_116_IS_ASYNC(M_AXIS_FIFO_116_IS_ASYNC),
        .M_AXIS_FIFO_117_IS_ASYNC(M_AXIS_FIFO_117_IS_ASYNC),
        .M_AXIS_FIFO_118_IS_ASYNC(M_AXIS_FIFO_118_IS_ASYNC),
        .M_AXIS_FIFO_119_IS_ASYNC(M_AXIS_FIFO_119_IS_ASYNC),
        .M_AXIS_FIFO_120_IS_ASYNC(M_AXIS_FIFO_120_IS_ASYNC),
        .M_AXIS_FIFO_121_IS_ASYNC(M_AXIS_FIFO_121_IS_ASYNC),
        .M_AXIS_FIFO_122_IS_ASYNC(M_AXIS_FIFO_122_IS_ASYNC),
        .M_AXIS_FIFO_123_IS_ASYNC(M_AXIS_FIFO_123_IS_ASYNC),
        .M_AXIS_FIFO_124_IS_ASYNC(M_AXIS_FIFO_124_IS_ASYNC),
        .M_AXIS_FIFO_125_IS_ASYNC(M_AXIS_FIFO_125_IS_ASYNC),
        .M_AXIS_FIFO_126_IS_ASYNC(M_AXIS_FIFO_126_IS_ASYNC),
        .M_AXIS_FIFO_127_IS_ASYNC(M_AXIS_FIFO_127_IS_ASYNC),
        .M_AXIS_FIFO_0_BYTE_WIDTH(M_AXIS_FIFO_0_BYTE_WIDTH),
        .M_AXIS_FIFO_1_BYTE_WIDTH(M_AXIS_FIFO_1_BYTE_WIDTH),
        .M_AXIS_FIFO_2_BYTE_WIDTH(M_AXIS_FIFO_2_BYTE_WIDTH),
        .M_AXIS_FIFO_3_BYTE_WIDTH(M_AXIS_FIFO_3_BYTE_WIDTH),
        .M_AXIS_FIFO_4_BYTE_WIDTH(M_AXIS_FIFO_4_BYTE_WIDTH),
        .M_AXIS_FIFO_5_BYTE_WIDTH(M_AXIS_FIFO_5_BYTE_WIDTH),
        .M_AXIS_FIFO_6_BYTE_WIDTH(M_AXIS_FIFO_6_BYTE_WIDTH),
        .M_AXIS_FIFO_7_BYTE_WIDTH(M_AXIS_FIFO_7_BYTE_WIDTH),
        .M_AXIS_FIFO_8_BYTE_WIDTH(M_AXIS_FIFO_8_BYTE_WIDTH),
        .M_AXIS_FIFO_9_BYTE_WIDTH(M_AXIS_FIFO_9_BYTE_WIDTH),
        .M_AXIS_FIFO_10_BYTE_WIDTH(M_AXIS_FIFO_10_BYTE_WIDTH),
        .M_AXIS_FIFO_11_BYTE_WIDTH(M_AXIS_FIFO_11_BYTE_WIDTH),
        .M_AXIS_FIFO_12_BYTE_WIDTH(M_AXIS_FIFO_12_BYTE_WIDTH),
        .M_AXIS_FIFO_13_BYTE_WIDTH(M_AXIS_FIFO_13_BYTE_WIDTH),
        .M_AXIS_FIFO_14_BYTE_WIDTH(M_AXIS_FIFO_14_BYTE_WIDTH),
        .M_AXIS_FIFO_15_BYTE_WIDTH(M_AXIS_FIFO_15_BYTE_WIDTH),
        .M_AXIS_FIFO_16_BYTE_WIDTH(M_AXIS_FIFO_16_BYTE_WIDTH),
        .M_AXIS_FIFO_17_BYTE_WIDTH(M_AXIS_FIFO_17_BYTE_WIDTH),
        .M_AXIS_FIFO_18_BYTE_WIDTH(M_AXIS_FIFO_18_BYTE_WIDTH),
        .M_AXIS_FIFO_19_BYTE_WIDTH(M_AXIS_FIFO_19_BYTE_WIDTH),
        .M_AXIS_FIFO_20_BYTE_WIDTH(M_AXIS_FIFO_20_BYTE_WIDTH),
        .M_AXIS_FIFO_21_BYTE_WIDTH(M_AXIS_FIFO_21_BYTE_WIDTH),
        .M_AXIS_FIFO_22_BYTE_WIDTH(M_AXIS_FIFO_22_BYTE_WIDTH),
        .M_AXIS_FIFO_23_BYTE_WIDTH(M_AXIS_FIFO_23_BYTE_WIDTH),
        .M_AXIS_FIFO_24_BYTE_WIDTH(M_AXIS_FIFO_24_BYTE_WIDTH),
        .M_AXIS_FIFO_25_BYTE_WIDTH(M_AXIS_FIFO_25_BYTE_WIDTH),
        .M_AXIS_FIFO_26_BYTE_WIDTH(M_AXIS_FIFO_26_BYTE_WIDTH),
        .M_AXIS_FIFO_27_BYTE_WIDTH(M_AXIS_FIFO_27_BYTE_WIDTH),
        .M_AXIS_FIFO_28_BYTE_WIDTH(M_AXIS_FIFO_28_BYTE_WIDTH),
        .M_AXIS_FIFO_29_BYTE_WIDTH(M_AXIS_FIFO_29_BYTE_WIDTH),
        .M_AXIS_FIFO_30_BYTE_WIDTH(M_AXIS_FIFO_30_BYTE_WIDTH),
        .M_AXIS_FIFO_31_BYTE_WIDTH(M_AXIS_FIFO_31_BYTE_WIDTH),
        .M_AXIS_FIFO_32_BYTE_WIDTH(M_AXIS_FIFO_32_BYTE_WIDTH),
        .M_AXIS_FIFO_33_BYTE_WIDTH(M_AXIS_FIFO_33_BYTE_WIDTH),
        .M_AXIS_FIFO_34_BYTE_WIDTH(M_AXIS_FIFO_34_BYTE_WIDTH),
        .M_AXIS_FIFO_35_BYTE_WIDTH(M_AXIS_FIFO_35_BYTE_WIDTH),
        .M_AXIS_FIFO_36_BYTE_WIDTH(M_AXIS_FIFO_36_BYTE_WIDTH),
        .M_AXIS_FIFO_37_BYTE_WIDTH(M_AXIS_FIFO_37_BYTE_WIDTH),
        .M_AXIS_FIFO_38_BYTE_WIDTH(M_AXIS_FIFO_38_BYTE_WIDTH),
        .M_AXIS_FIFO_39_BYTE_WIDTH(M_AXIS_FIFO_39_BYTE_WIDTH),
        .M_AXIS_FIFO_40_BYTE_WIDTH(M_AXIS_FIFO_40_BYTE_WIDTH),
        .M_AXIS_FIFO_41_BYTE_WIDTH(M_AXIS_FIFO_41_BYTE_WIDTH),
        .M_AXIS_FIFO_42_BYTE_WIDTH(M_AXIS_FIFO_42_BYTE_WIDTH),
        .M_AXIS_FIFO_43_BYTE_WIDTH(M_AXIS_FIFO_43_BYTE_WIDTH),
        .M_AXIS_FIFO_44_BYTE_WIDTH(M_AXIS_FIFO_44_BYTE_WIDTH),
        .M_AXIS_FIFO_45_BYTE_WIDTH(M_AXIS_FIFO_45_BYTE_WIDTH),
        .M_AXIS_FIFO_46_BYTE_WIDTH(M_AXIS_FIFO_46_BYTE_WIDTH),
        .M_AXIS_FIFO_47_BYTE_WIDTH(M_AXIS_FIFO_47_BYTE_WIDTH),
        .M_AXIS_FIFO_48_BYTE_WIDTH(M_AXIS_FIFO_48_BYTE_WIDTH),
        .M_AXIS_FIFO_49_BYTE_WIDTH(M_AXIS_FIFO_49_BYTE_WIDTH),
        .M_AXIS_FIFO_50_BYTE_WIDTH(M_AXIS_FIFO_50_BYTE_WIDTH),
        .M_AXIS_FIFO_51_BYTE_WIDTH(M_AXIS_FIFO_51_BYTE_WIDTH),
        .M_AXIS_FIFO_52_BYTE_WIDTH(M_AXIS_FIFO_52_BYTE_WIDTH),
        .M_AXIS_FIFO_53_BYTE_WIDTH(M_AXIS_FIFO_53_BYTE_WIDTH),
        .M_AXIS_FIFO_54_BYTE_WIDTH(M_AXIS_FIFO_54_BYTE_WIDTH),
        .M_AXIS_FIFO_55_BYTE_WIDTH(M_AXIS_FIFO_55_BYTE_WIDTH),
        .M_AXIS_FIFO_56_BYTE_WIDTH(M_AXIS_FIFO_56_BYTE_WIDTH),
        .M_AXIS_FIFO_57_BYTE_WIDTH(M_AXIS_FIFO_57_BYTE_WIDTH),
        .M_AXIS_FIFO_58_BYTE_WIDTH(M_AXIS_FIFO_58_BYTE_WIDTH),
        .M_AXIS_FIFO_59_BYTE_WIDTH(M_AXIS_FIFO_59_BYTE_WIDTH),
        .M_AXIS_FIFO_60_BYTE_WIDTH(M_AXIS_FIFO_60_BYTE_WIDTH),
        .M_AXIS_FIFO_61_BYTE_WIDTH(M_AXIS_FIFO_61_BYTE_WIDTH),
        .M_AXIS_FIFO_62_BYTE_WIDTH(M_AXIS_FIFO_62_BYTE_WIDTH),
        .M_AXIS_FIFO_63_BYTE_WIDTH(M_AXIS_FIFO_63_BYTE_WIDTH),
        .M_AXIS_FIFO_64_BYTE_WIDTH(M_AXIS_FIFO_64_BYTE_WIDTH),
        .M_AXIS_FIFO_65_BYTE_WIDTH(M_AXIS_FIFO_65_BYTE_WIDTH),
        .M_AXIS_FIFO_66_BYTE_WIDTH(M_AXIS_FIFO_66_BYTE_WIDTH),
        .M_AXIS_FIFO_67_BYTE_WIDTH(M_AXIS_FIFO_67_BYTE_WIDTH),
        .M_AXIS_FIFO_68_BYTE_WIDTH(M_AXIS_FIFO_68_BYTE_WIDTH),
        .M_AXIS_FIFO_69_BYTE_WIDTH(M_AXIS_FIFO_69_BYTE_WIDTH),
        .M_AXIS_FIFO_70_BYTE_WIDTH(M_AXIS_FIFO_70_BYTE_WIDTH),
        .M_AXIS_FIFO_71_BYTE_WIDTH(M_AXIS_FIFO_71_BYTE_WIDTH),
        .M_AXIS_FIFO_72_BYTE_WIDTH(M_AXIS_FIFO_72_BYTE_WIDTH),
        .M_AXIS_FIFO_73_BYTE_WIDTH(M_AXIS_FIFO_73_BYTE_WIDTH),
        .M_AXIS_FIFO_74_BYTE_WIDTH(M_AXIS_FIFO_74_BYTE_WIDTH),
        .M_AXIS_FIFO_75_BYTE_WIDTH(M_AXIS_FIFO_75_BYTE_WIDTH),
        .M_AXIS_FIFO_76_BYTE_WIDTH(M_AXIS_FIFO_76_BYTE_WIDTH),
        .M_AXIS_FIFO_77_BYTE_WIDTH(M_AXIS_FIFO_77_BYTE_WIDTH),
        .M_AXIS_FIFO_78_BYTE_WIDTH(M_AXIS_FIFO_78_BYTE_WIDTH),
        .M_AXIS_FIFO_79_BYTE_WIDTH(M_AXIS_FIFO_79_BYTE_WIDTH),
        .M_AXIS_FIFO_80_BYTE_WIDTH(M_AXIS_FIFO_80_BYTE_WIDTH),
        .M_AXIS_FIFO_81_BYTE_WIDTH(M_AXIS_FIFO_81_BYTE_WIDTH),
        .M_AXIS_FIFO_82_BYTE_WIDTH(M_AXIS_FIFO_82_BYTE_WIDTH),
        .M_AXIS_FIFO_83_BYTE_WIDTH(M_AXIS_FIFO_83_BYTE_WIDTH),
        .M_AXIS_FIFO_84_BYTE_WIDTH(M_AXIS_FIFO_84_BYTE_WIDTH),
        .M_AXIS_FIFO_85_BYTE_WIDTH(M_AXIS_FIFO_85_BYTE_WIDTH),
        .M_AXIS_FIFO_86_BYTE_WIDTH(M_AXIS_FIFO_86_BYTE_WIDTH),
        .M_AXIS_FIFO_87_BYTE_WIDTH(M_AXIS_FIFO_87_BYTE_WIDTH),
        .M_AXIS_FIFO_88_BYTE_WIDTH(M_AXIS_FIFO_88_BYTE_WIDTH),
        .M_AXIS_FIFO_89_BYTE_WIDTH(M_AXIS_FIFO_89_BYTE_WIDTH),
        .M_AXIS_FIFO_90_BYTE_WIDTH(M_AXIS_FIFO_90_BYTE_WIDTH),
        .M_AXIS_FIFO_91_BYTE_WIDTH(M_AXIS_FIFO_91_BYTE_WIDTH),
        .M_AXIS_FIFO_92_BYTE_WIDTH(M_AXIS_FIFO_92_BYTE_WIDTH),
        .M_AXIS_FIFO_93_BYTE_WIDTH(M_AXIS_FIFO_93_BYTE_WIDTH),
        .M_AXIS_FIFO_94_BYTE_WIDTH(M_AXIS_FIFO_94_BYTE_WIDTH),
        .M_AXIS_FIFO_95_BYTE_WIDTH(M_AXIS_FIFO_95_BYTE_WIDTH),
        .M_AXIS_FIFO_96_BYTE_WIDTH(M_AXIS_FIFO_96_BYTE_WIDTH),
        .M_AXIS_FIFO_97_BYTE_WIDTH(M_AXIS_FIFO_97_BYTE_WIDTH),
        .M_AXIS_FIFO_98_BYTE_WIDTH(M_AXIS_FIFO_98_BYTE_WIDTH),
        .M_AXIS_FIFO_99_BYTE_WIDTH(M_AXIS_FIFO_99_BYTE_WIDTH),
        .M_AXIS_FIFO_100_BYTE_WIDTH(M_AXIS_FIFO_100_BYTE_WIDTH),
        .M_AXIS_FIFO_101_BYTE_WIDTH(M_AXIS_FIFO_101_BYTE_WIDTH),
        .M_AXIS_FIFO_102_BYTE_WIDTH(M_AXIS_FIFO_102_BYTE_WIDTH),
        .M_AXIS_FIFO_103_BYTE_WIDTH(M_AXIS_FIFO_103_BYTE_WIDTH),
        .M_AXIS_FIFO_104_BYTE_WIDTH(M_AXIS_FIFO_104_BYTE_WIDTH),
        .M_AXIS_FIFO_105_BYTE_WIDTH(M_AXIS_FIFO_105_BYTE_WIDTH),
        .M_AXIS_FIFO_106_BYTE_WIDTH(M_AXIS_FIFO_106_BYTE_WIDTH),
        .M_AXIS_FIFO_107_BYTE_WIDTH(M_AXIS_FIFO_107_BYTE_WIDTH),
        .M_AXIS_FIFO_108_BYTE_WIDTH(M_AXIS_FIFO_108_BYTE_WIDTH),
        .M_AXIS_FIFO_109_BYTE_WIDTH(M_AXIS_FIFO_109_BYTE_WIDTH),
        .M_AXIS_FIFO_110_BYTE_WIDTH(M_AXIS_FIFO_110_BYTE_WIDTH),
        .M_AXIS_FIFO_111_BYTE_WIDTH(M_AXIS_FIFO_111_BYTE_WIDTH),
        .M_AXIS_FIFO_112_BYTE_WIDTH(M_AXIS_FIFO_112_BYTE_WIDTH),
        .M_AXIS_FIFO_113_BYTE_WIDTH(M_AXIS_FIFO_113_BYTE_WIDTH),
        .M_AXIS_FIFO_114_BYTE_WIDTH(M_AXIS_FIFO_114_BYTE_WIDTH),
        .M_AXIS_FIFO_115_BYTE_WIDTH(M_AXIS_FIFO_115_BYTE_WIDTH),
        .M_AXIS_FIFO_116_BYTE_WIDTH(M_AXIS_FIFO_116_BYTE_WIDTH),
        .M_AXIS_FIFO_117_BYTE_WIDTH(M_AXIS_FIFO_117_BYTE_WIDTH),
        .M_AXIS_FIFO_118_BYTE_WIDTH(M_AXIS_FIFO_118_BYTE_WIDTH),
        .M_AXIS_FIFO_119_BYTE_WIDTH(M_AXIS_FIFO_119_BYTE_WIDTH),
        .M_AXIS_FIFO_120_BYTE_WIDTH(M_AXIS_FIFO_120_BYTE_WIDTH),
        .M_AXIS_FIFO_121_BYTE_WIDTH(M_AXIS_FIFO_121_BYTE_WIDTH),
        .M_AXIS_FIFO_122_BYTE_WIDTH(M_AXIS_FIFO_122_BYTE_WIDTH),
        .M_AXIS_FIFO_123_BYTE_WIDTH(M_AXIS_FIFO_123_BYTE_WIDTH),
        .M_AXIS_FIFO_124_BYTE_WIDTH(M_AXIS_FIFO_124_BYTE_WIDTH),
        .M_AXIS_FIFO_125_BYTE_WIDTH(M_AXIS_FIFO_125_BYTE_WIDTH),
        .M_AXIS_FIFO_126_BYTE_WIDTH(M_AXIS_FIFO_126_BYTE_WIDTH),
        .M_AXIS_FIFO_127_BYTE_WIDTH(M_AXIS_FIFO_127_BYTE_WIDTH),
        .M_AXIS_FIFO_0_DMWIDTH(M_AXIS_FIFO_0_DMWIDTH),
        .M_AXIS_FIFO_1_DMWIDTH(M_AXIS_FIFO_1_DMWIDTH),
        .M_AXIS_FIFO_2_DMWIDTH(M_AXIS_FIFO_2_DMWIDTH),
        .M_AXIS_FIFO_3_DMWIDTH(M_AXIS_FIFO_3_DMWIDTH),
        .M_AXIS_FIFO_4_DMWIDTH(M_AXIS_FIFO_4_DMWIDTH),
        .M_AXIS_FIFO_5_DMWIDTH(M_AXIS_FIFO_5_DMWIDTH),
        .M_AXIS_FIFO_6_DMWIDTH(M_AXIS_FIFO_6_DMWIDTH),
        .M_AXIS_FIFO_7_DMWIDTH(M_AXIS_FIFO_7_DMWIDTH),
        .M_AXIS_FIFO_8_DMWIDTH(M_AXIS_FIFO_8_DMWIDTH),
        .M_AXIS_FIFO_9_DMWIDTH(M_AXIS_FIFO_9_DMWIDTH),
        .M_AXIS_FIFO_10_DMWIDTH(M_AXIS_FIFO_10_DMWIDTH),
        .M_AXIS_FIFO_11_DMWIDTH(M_AXIS_FIFO_11_DMWIDTH),
        .M_AXIS_FIFO_12_DMWIDTH(M_AXIS_FIFO_12_DMWIDTH),
        .M_AXIS_FIFO_13_DMWIDTH(M_AXIS_FIFO_13_DMWIDTH),
        .M_AXIS_FIFO_14_DMWIDTH(M_AXIS_FIFO_14_DMWIDTH),
        .M_AXIS_FIFO_15_DMWIDTH(M_AXIS_FIFO_15_DMWIDTH),
        .M_AXIS_FIFO_16_DMWIDTH(M_AXIS_FIFO_16_DMWIDTH),
        .M_AXIS_FIFO_17_DMWIDTH(M_AXIS_FIFO_17_DMWIDTH),
        .M_AXIS_FIFO_18_DMWIDTH(M_AXIS_FIFO_18_DMWIDTH),
        .M_AXIS_FIFO_19_DMWIDTH(M_AXIS_FIFO_19_DMWIDTH),
        .M_AXIS_FIFO_20_DMWIDTH(M_AXIS_FIFO_20_DMWIDTH),
        .M_AXIS_FIFO_21_DMWIDTH(M_AXIS_FIFO_21_DMWIDTH),
        .M_AXIS_FIFO_22_DMWIDTH(M_AXIS_FIFO_22_DMWIDTH),
        .M_AXIS_FIFO_23_DMWIDTH(M_AXIS_FIFO_23_DMWIDTH),
        .M_AXIS_FIFO_24_DMWIDTH(M_AXIS_FIFO_24_DMWIDTH),
        .M_AXIS_FIFO_25_DMWIDTH(M_AXIS_FIFO_25_DMWIDTH),
        .M_AXIS_FIFO_26_DMWIDTH(M_AXIS_FIFO_26_DMWIDTH),
        .M_AXIS_FIFO_27_DMWIDTH(M_AXIS_FIFO_27_DMWIDTH),
        .M_AXIS_FIFO_28_DMWIDTH(M_AXIS_FIFO_28_DMWIDTH),
        .M_AXIS_FIFO_29_DMWIDTH(M_AXIS_FIFO_29_DMWIDTH),
        .M_AXIS_FIFO_30_DMWIDTH(M_AXIS_FIFO_30_DMWIDTH),
        .M_AXIS_FIFO_31_DMWIDTH(M_AXIS_FIFO_31_DMWIDTH),
        .M_AXIS_FIFO_32_DMWIDTH(M_AXIS_FIFO_32_DMWIDTH),
        .M_AXIS_FIFO_33_DMWIDTH(M_AXIS_FIFO_33_DMWIDTH),
        .M_AXIS_FIFO_34_DMWIDTH(M_AXIS_FIFO_34_DMWIDTH),
        .M_AXIS_FIFO_35_DMWIDTH(M_AXIS_FIFO_35_DMWIDTH),
        .M_AXIS_FIFO_36_DMWIDTH(M_AXIS_FIFO_36_DMWIDTH),
        .M_AXIS_FIFO_37_DMWIDTH(M_AXIS_FIFO_37_DMWIDTH),
        .M_AXIS_FIFO_38_DMWIDTH(M_AXIS_FIFO_38_DMWIDTH),
        .M_AXIS_FIFO_39_DMWIDTH(M_AXIS_FIFO_39_DMWIDTH),
        .M_AXIS_FIFO_40_DMWIDTH(M_AXIS_FIFO_40_DMWIDTH),
        .M_AXIS_FIFO_41_DMWIDTH(M_AXIS_FIFO_41_DMWIDTH),
        .M_AXIS_FIFO_42_DMWIDTH(M_AXIS_FIFO_42_DMWIDTH),
        .M_AXIS_FIFO_43_DMWIDTH(M_AXIS_FIFO_43_DMWIDTH),
        .M_AXIS_FIFO_44_DMWIDTH(M_AXIS_FIFO_44_DMWIDTH),
        .M_AXIS_FIFO_45_DMWIDTH(M_AXIS_FIFO_45_DMWIDTH),
        .M_AXIS_FIFO_46_DMWIDTH(M_AXIS_FIFO_46_DMWIDTH),
        .M_AXIS_FIFO_47_DMWIDTH(M_AXIS_FIFO_47_DMWIDTH),
        .M_AXIS_FIFO_48_DMWIDTH(M_AXIS_FIFO_48_DMWIDTH),
        .M_AXIS_FIFO_49_DMWIDTH(M_AXIS_FIFO_49_DMWIDTH),
        .M_AXIS_FIFO_50_DMWIDTH(M_AXIS_FIFO_50_DMWIDTH),
        .M_AXIS_FIFO_51_DMWIDTH(M_AXIS_FIFO_51_DMWIDTH),
        .M_AXIS_FIFO_52_DMWIDTH(M_AXIS_FIFO_52_DMWIDTH),
        .M_AXIS_FIFO_53_DMWIDTH(M_AXIS_FIFO_53_DMWIDTH),
        .M_AXIS_FIFO_54_DMWIDTH(M_AXIS_FIFO_54_DMWIDTH),
        .M_AXIS_FIFO_55_DMWIDTH(M_AXIS_FIFO_55_DMWIDTH),
        .M_AXIS_FIFO_56_DMWIDTH(M_AXIS_FIFO_56_DMWIDTH),
        .M_AXIS_FIFO_57_DMWIDTH(M_AXIS_FIFO_57_DMWIDTH),
        .M_AXIS_FIFO_58_DMWIDTH(M_AXIS_FIFO_58_DMWIDTH),
        .M_AXIS_FIFO_59_DMWIDTH(M_AXIS_FIFO_59_DMWIDTH),
        .M_AXIS_FIFO_60_DMWIDTH(M_AXIS_FIFO_60_DMWIDTH),
        .M_AXIS_FIFO_61_DMWIDTH(M_AXIS_FIFO_61_DMWIDTH),
        .M_AXIS_FIFO_62_DMWIDTH(M_AXIS_FIFO_62_DMWIDTH),
        .M_AXIS_FIFO_63_DMWIDTH(M_AXIS_FIFO_63_DMWIDTH),
        .M_AXIS_FIFO_64_DMWIDTH(M_AXIS_FIFO_64_DMWIDTH),
        .M_AXIS_FIFO_65_DMWIDTH(M_AXIS_FIFO_65_DMWIDTH),
        .M_AXIS_FIFO_66_DMWIDTH(M_AXIS_FIFO_66_DMWIDTH),
        .M_AXIS_FIFO_67_DMWIDTH(M_AXIS_FIFO_67_DMWIDTH),
        .M_AXIS_FIFO_68_DMWIDTH(M_AXIS_FIFO_68_DMWIDTH),
        .M_AXIS_FIFO_69_DMWIDTH(M_AXIS_FIFO_69_DMWIDTH),
        .M_AXIS_FIFO_70_DMWIDTH(M_AXIS_FIFO_70_DMWIDTH),
        .M_AXIS_FIFO_71_DMWIDTH(M_AXIS_FIFO_71_DMWIDTH),
        .M_AXIS_FIFO_72_DMWIDTH(M_AXIS_FIFO_72_DMWIDTH),
        .M_AXIS_FIFO_73_DMWIDTH(M_AXIS_FIFO_73_DMWIDTH),
        .M_AXIS_FIFO_74_DMWIDTH(M_AXIS_FIFO_74_DMWIDTH),
        .M_AXIS_FIFO_75_DMWIDTH(M_AXIS_FIFO_75_DMWIDTH),
        .M_AXIS_FIFO_76_DMWIDTH(M_AXIS_FIFO_76_DMWIDTH),
        .M_AXIS_FIFO_77_DMWIDTH(M_AXIS_FIFO_77_DMWIDTH),
        .M_AXIS_FIFO_78_DMWIDTH(M_AXIS_FIFO_78_DMWIDTH),
        .M_AXIS_FIFO_79_DMWIDTH(M_AXIS_FIFO_79_DMWIDTH),
        .M_AXIS_FIFO_80_DMWIDTH(M_AXIS_FIFO_80_DMWIDTH),
        .M_AXIS_FIFO_81_DMWIDTH(M_AXIS_FIFO_81_DMWIDTH),
        .M_AXIS_FIFO_82_DMWIDTH(M_AXIS_FIFO_82_DMWIDTH),
        .M_AXIS_FIFO_83_DMWIDTH(M_AXIS_FIFO_83_DMWIDTH),
        .M_AXIS_FIFO_84_DMWIDTH(M_AXIS_FIFO_84_DMWIDTH),
        .M_AXIS_FIFO_85_DMWIDTH(M_AXIS_FIFO_85_DMWIDTH),
        .M_AXIS_FIFO_86_DMWIDTH(M_AXIS_FIFO_86_DMWIDTH),
        .M_AXIS_FIFO_87_DMWIDTH(M_AXIS_FIFO_87_DMWIDTH),
        .M_AXIS_FIFO_88_DMWIDTH(M_AXIS_FIFO_88_DMWIDTH),
        .M_AXIS_FIFO_89_DMWIDTH(M_AXIS_FIFO_89_DMWIDTH),
        .M_AXIS_FIFO_90_DMWIDTH(M_AXIS_FIFO_90_DMWIDTH),
        .M_AXIS_FIFO_91_DMWIDTH(M_AXIS_FIFO_91_DMWIDTH),
        .M_AXIS_FIFO_92_DMWIDTH(M_AXIS_FIFO_92_DMWIDTH),
        .M_AXIS_FIFO_93_DMWIDTH(M_AXIS_FIFO_93_DMWIDTH),
        .M_AXIS_FIFO_94_DMWIDTH(M_AXIS_FIFO_94_DMWIDTH),
        .M_AXIS_FIFO_95_DMWIDTH(M_AXIS_FIFO_95_DMWIDTH),
        .M_AXIS_FIFO_96_DMWIDTH(M_AXIS_FIFO_96_DMWIDTH),
        .M_AXIS_FIFO_97_DMWIDTH(M_AXIS_FIFO_97_DMWIDTH),
        .M_AXIS_FIFO_98_DMWIDTH(M_AXIS_FIFO_98_DMWIDTH),
        .M_AXIS_FIFO_99_DMWIDTH(M_AXIS_FIFO_99_DMWIDTH),
        .M_AXIS_FIFO_100_DMWIDTH(M_AXIS_FIFO_100_DMWIDTH),
        .M_AXIS_FIFO_101_DMWIDTH(M_AXIS_FIFO_101_DMWIDTH),
        .M_AXIS_FIFO_102_DMWIDTH(M_AXIS_FIFO_102_DMWIDTH),
        .M_AXIS_FIFO_103_DMWIDTH(M_AXIS_FIFO_103_DMWIDTH),
        .M_AXIS_FIFO_104_DMWIDTH(M_AXIS_FIFO_104_DMWIDTH),
        .M_AXIS_FIFO_105_DMWIDTH(M_AXIS_FIFO_105_DMWIDTH),
        .M_AXIS_FIFO_106_DMWIDTH(M_AXIS_FIFO_106_DMWIDTH),
        .M_AXIS_FIFO_107_DMWIDTH(M_AXIS_FIFO_107_DMWIDTH),
        .M_AXIS_FIFO_108_DMWIDTH(M_AXIS_FIFO_108_DMWIDTH),
        .M_AXIS_FIFO_109_DMWIDTH(M_AXIS_FIFO_109_DMWIDTH),
        .M_AXIS_FIFO_110_DMWIDTH(M_AXIS_FIFO_110_DMWIDTH),
        .M_AXIS_FIFO_111_DMWIDTH(M_AXIS_FIFO_111_DMWIDTH),
        .M_AXIS_FIFO_112_DMWIDTH(M_AXIS_FIFO_112_DMWIDTH),
        .M_AXIS_FIFO_113_DMWIDTH(M_AXIS_FIFO_113_DMWIDTH),
        .M_AXIS_FIFO_114_DMWIDTH(M_AXIS_FIFO_114_DMWIDTH),
        .M_AXIS_FIFO_115_DMWIDTH(M_AXIS_FIFO_115_DMWIDTH),
        .M_AXIS_FIFO_116_DMWIDTH(M_AXIS_FIFO_116_DMWIDTH),
        .M_AXIS_FIFO_117_DMWIDTH(M_AXIS_FIFO_117_DMWIDTH),
        .M_AXIS_FIFO_118_DMWIDTH(M_AXIS_FIFO_118_DMWIDTH),
        .M_AXIS_FIFO_119_DMWIDTH(M_AXIS_FIFO_119_DMWIDTH),
        .M_AXIS_FIFO_120_DMWIDTH(M_AXIS_FIFO_120_DMWIDTH),
        .M_AXIS_FIFO_121_DMWIDTH(M_AXIS_FIFO_121_DMWIDTH),
        .M_AXIS_FIFO_122_DMWIDTH(M_AXIS_FIFO_122_DMWIDTH),
        .M_AXIS_FIFO_123_DMWIDTH(M_AXIS_FIFO_123_DMWIDTH),
        .M_AXIS_FIFO_124_DMWIDTH(M_AXIS_FIFO_124_DMWIDTH),
        .M_AXIS_FIFO_125_DMWIDTH(M_AXIS_FIFO_125_DMWIDTH),
        .M_AXIS_FIFO_126_DMWIDTH(M_AXIS_FIFO_126_DMWIDTH),
        .M_AXIS_FIFO_127_DMWIDTH(M_AXIS_FIFO_127_DMWIDTH)
    ) out_fifo_args_i (
        .acc_clk(acc_aclk),
        .acc_aresetn(acc_aresetn),
        .out_fifo_allow(outfifo_ctrl_allow),
        .m_axis_fifo_0_aclk(m_axis_fifo_0_aclk),
        .m_axis_fifo_0_aresetn(m_axis_fifo_0_aresetn),
        .m_axis_fifo_0_tlast(m_axis_fifo_0_tlast),
        .m_axis_fifo_0_tvalid(m_axis_fifo_0_tvalid),
        .m_axis_fifo_0_tkeep(m_axis_fifo_0_tkeep),
        .m_axis_fifo_0_tstrb(m_axis_fifo_0_tstrb),
        .m_axis_fifo_0_tdata(m_axis_fifo_0_tdata),
        .m_axis_fifo_0_tready(m_axis_fifo_0_tready),
        .ap_fifo_oarg_0_full_n(ap_fifo_oarg_0_full_n),
        .ap_fifo_oarg_0_din(ap_fifo_oarg_0_din),
        .ap_fifo_oarg_0_write(ap_fifo_oarg_0_write),
        .m_axis_fifo_1_aclk(m_axis_fifo_1_aclk),
        .m_axis_fifo_1_aresetn(m_axis_fifo_1_aresetn),
        .m_axis_fifo_1_tlast(m_axis_fifo_1_tlast),
        .m_axis_fifo_1_tvalid(m_axis_fifo_1_tvalid),
        .m_axis_fifo_1_tkeep(m_axis_fifo_1_tkeep),
        .m_axis_fifo_1_tstrb(m_axis_fifo_1_tstrb),
        .m_axis_fifo_1_tdata(m_axis_fifo_1_tdata),
        .m_axis_fifo_1_tready(m_axis_fifo_1_tready),
        .ap_fifo_oarg_1_full_n(ap_fifo_oarg_1_full_n),
        .ap_fifo_oarg_1_din(ap_fifo_oarg_1_din),
        .ap_fifo_oarg_1_write(ap_fifo_oarg_1_write),
        .m_axis_fifo_2_aclk(m_axis_fifo_2_aclk),
        .m_axis_fifo_2_aresetn(m_axis_fifo_2_aresetn),
        .m_axis_fifo_2_tlast(m_axis_fifo_2_tlast),
        .m_axis_fifo_2_tvalid(m_axis_fifo_2_tvalid),
        .m_axis_fifo_2_tkeep(m_axis_fifo_2_tkeep),
        .m_axis_fifo_2_tstrb(m_axis_fifo_2_tstrb),
        .m_axis_fifo_2_tdata(m_axis_fifo_2_tdata),
        .m_axis_fifo_2_tready(m_axis_fifo_2_tready),
        .ap_fifo_oarg_2_full_n(ap_fifo_oarg_2_full_n),
        .ap_fifo_oarg_2_din(ap_fifo_oarg_2_din),
        .ap_fifo_oarg_2_write(ap_fifo_oarg_2_write),
        .m_axis_fifo_3_aclk(m_axis_fifo_3_aclk),
        .m_axis_fifo_3_aresetn(m_axis_fifo_3_aresetn),
        .m_axis_fifo_3_tlast(m_axis_fifo_3_tlast),
        .m_axis_fifo_3_tvalid(m_axis_fifo_3_tvalid),
        .m_axis_fifo_3_tkeep(m_axis_fifo_3_tkeep),
        .m_axis_fifo_3_tstrb(m_axis_fifo_3_tstrb),
        .m_axis_fifo_3_tdata(m_axis_fifo_3_tdata),
        .m_axis_fifo_3_tready(m_axis_fifo_3_tready),
        .ap_fifo_oarg_3_full_n(ap_fifo_oarg_3_full_n),
        .ap_fifo_oarg_3_din(ap_fifo_oarg_3_din),
        .ap_fifo_oarg_3_write(ap_fifo_oarg_3_write),
        .m_axis_fifo_4_aclk(m_axis_fifo_4_aclk),
        .m_axis_fifo_4_aresetn(m_axis_fifo_4_aresetn),
        .m_axis_fifo_4_tlast(m_axis_fifo_4_tlast),
        .m_axis_fifo_4_tvalid(m_axis_fifo_4_tvalid),
        .m_axis_fifo_4_tkeep(m_axis_fifo_4_tkeep),
        .m_axis_fifo_4_tstrb(m_axis_fifo_4_tstrb),
        .m_axis_fifo_4_tdata(m_axis_fifo_4_tdata),
        .m_axis_fifo_4_tready(m_axis_fifo_4_tready),
        .ap_fifo_oarg_4_full_n(ap_fifo_oarg_4_full_n),
        .ap_fifo_oarg_4_din(ap_fifo_oarg_4_din),
        .ap_fifo_oarg_4_write(ap_fifo_oarg_4_write),
        .m_axis_fifo_5_aclk(m_axis_fifo_5_aclk),
        .m_axis_fifo_5_aresetn(m_axis_fifo_5_aresetn),
        .m_axis_fifo_5_tlast(m_axis_fifo_5_tlast),
        .m_axis_fifo_5_tvalid(m_axis_fifo_5_tvalid),
        .m_axis_fifo_5_tkeep(m_axis_fifo_5_tkeep),
        .m_axis_fifo_5_tstrb(m_axis_fifo_5_tstrb),
        .m_axis_fifo_5_tdata(m_axis_fifo_5_tdata),
        .m_axis_fifo_5_tready(m_axis_fifo_5_tready),
        .ap_fifo_oarg_5_full_n(ap_fifo_oarg_5_full_n),
        .ap_fifo_oarg_5_din(ap_fifo_oarg_5_din),
        .ap_fifo_oarg_5_write(ap_fifo_oarg_5_write),
        .m_axis_fifo_6_aclk(m_axis_fifo_6_aclk),
        .m_axis_fifo_6_aresetn(m_axis_fifo_6_aresetn),
        .m_axis_fifo_6_tlast(m_axis_fifo_6_tlast),
        .m_axis_fifo_6_tvalid(m_axis_fifo_6_tvalid),
        .m_axis_fifo_6_tkeep(m_axis_fifo_6_tkeep),
        .m_axis_fifo_6_tstrb(m_axis_fifo_6_tstrb),
        .m_axis_fifo_6_tdata(m_axis_fifo_6_tdata),
        .m_axis_fifo_6_tready(m_axis_fifo_6_tready),
        .ap_fifo_oarg_6_full_n(ap_fifo_oarg_6_full_n),
        .ap_fifo_oarg_6_din(ap_fifo_oarg_6_din),
        .ap_fifo_oarg_6_write(ap_fifo_oarg_6_write),
        .m_axis_fifo_7_aclk(m_axis_fifo_7_aclk),
        .m_axis_fifo_7_aresetn(m_axis_fifo_7_aresetn),
        .m_axis_fifo_7_tlast(m_axis_fifo_7_tlast),
        .m_axis_fifo_7_tvalid(m_axis_fifo_7_tvalid),
        .m_axis_fifo_7_tkeep(m_axis_fifo_7_tkeep),
        .m_axis_fifo_7_tstrb(m_axis_fifo_7_tstrb),
        .m_axis_fifo_7_tdata(m_axis_fifo_7_tdata),
        .m_axis_fifo_7_tready(m_axis_fifo_7_tready),
        .ap_fifo_oarg_7_full_n(ap_fifo_oarg_7_full_n),
        .ap_fifo_oarg_7_din(ap_fifo_oarg_7_din),
        .ap_fifo_oarg_7_write(ap_fifo_oarg_7_write),
        .m_axis_fifo_8_aclk(m_axis_fifo_8_aclk),
        .m_axis_fifo_8_aresetn(m_axis_fifo_8_aresetn),
        .m_axis_fifo_8_tlast(m_axis_fifo_8_tlast),
        .m_axis_fifo_8_tvalid(m_axis_fifo_8_tvalid),
        .m_axis_fifo_8_tkeep(m_axis_fifo_8_tkeep),
        .m_axis_fifo_8_tstrb(m_axis_fifo_8_tstrb),
        .m_axis_fifo_8_tdata(m_axis_fifo_8_tdata),
        .m_axis_fifo_8_tready(m_axis_fifo_8_tready),
        .ap_fifo_oarg_8_full_n(ap_fifo_oarg_8_full_n),
        .ap_fifo_oarg_8_din(ap_fifo_oarg_8_din),
        .ap_fifo_oarg_8_write(ap_fifo_oarg_8_write),
        .m_axis_fifo_9_aclk(m_axis_fifo_9_aclk),
        .m_axis_fifo_9_aresetn(m_axis_fifo_9_aresetn),
        .m_axis_fifo_9_tlast(m_axis_fifo_9_tlast),
        .m_axis_fifo_9_tvalid(m_axis_fifo_9_tvalid),
        .m_axis_fifo_9_tkeep(m_axis_fifo_9_tkeep),
        .m_axis_fifo_9_tstrb(m_axis_fifo_9_tstrb),
        .m_axis_fifo_9_tdata(m_axis_fifo_9_tdata),
        .m_axis_fifo_9_tready(m_axis_fifo_9_tready),
        .ap_fifo_oarg_9_full_n(ap_fifo_oarg_9_full_n),
        .ap_fifo_oarg_9_din(ap_fifo_oarg_9_din),
        .ap_fifo_oarg_9_write(ap_fifo_oarg_9_write),
        .m_axis_fifo_10_aclk(m_axis_fifo_10_aclk),
        .m_axis_fifo_10_aresetn(m_axis_fifo_10_aresetn),
        .m_axis_fifo_10_tlast(m_axis_fifo_10_tlast),
        .m_axis_fifo_10_tvalid(m_axis_fifo_10_tvalid),
        .m_axis_fifo_10_tkeep(m_axis_fifo_10_tkeep),
        .m_axis_fifo_10_tstrb(m_axis_fifo_10_tstrb),
        .m_axis_fifo_10_tdata(m_axis_fifo_10_tdata),
        .m_axis_fifo_10_tready(m_axis_fifo_10_tready),
        .ap_fifo_oarg_10_full_n(ap_fifo_oarg_10_full_n),
        .ap_fifo_oarg_10_din(ap_fifo_oarg_10_din),
        .ap_fifo_oarg_10_write(ap_fifo_oarg_10_write),
        .m_axis_fifo_11_aclk(m_axis_fifo_11_aclk),
        .m_axis_fifo_11_aresetn(m_axis_fifo_11_aresetn),
        .m_axis_fifo_11_tlast(m_axis_fifo_11_tlast),
        .m_axis_fifo_11_tvalid(m_axis_fifo_11_tvalid),
        .m_axis_fifo_11_tkeep(m_axis_fifo_11_tkeep),
        .m_axis_fifo_11_tstrb(m_axis_fifo_11_tstrb),
        .m_axis_fifo_11_tdata(m_axis_fifo_11_tdata),
        .m_axis_fifo_11_tready(m_axis_fifo_11_tready),
        .ap_fifo_oarg_11_full_n(ap_fifo_oarg_11_full_n),
        .ap_fifo_oarg_11_din(ap_fifo_oarg_11_din),
        .ap_fifo_oarg_11_write(ap_fifo_oarg_11_write),
        .m_axis_fifo_12_aclk(m_axis_fifo_12_aclk),
        .m_axis_fifo_12_aresetn(m_axis_fifo_12_aresetn),
        .m_axis_fifo_12_tlast(m_axis_fifo_12_tlast),
        .m_axis_fifo_12_tvalid(m_axis_fifo_12_tvalid),
        .m_axis_fifo_12_tkeep(m_axis_fifo_12_tkeep),
        .m_axis_fifo_12_tstrb(m_axis_fifo_12_tstrb),
        .m_axis_fifo_12_tdata(m_axis_fifo_12_tdata),
        .m_axis_fifo_12_tready(m_axis_fifo_12_tready),
        .ap_fifo_oarg_12_full_n(ap_fifo_oarg_12_full_n),
        .ap_fifo_oarg_12_din(ap_fifo_oarg_12_din),
        .ap_fifo_oarg_12_write(ap_fifo_oarg_12_write),
        .m_axis_fifo_13_aclk(m_axis_fifo_13_aclk),
        .m_axis_fifo_13_aresetn(m_axis_fifo_13_aresetn),
        .m_axis_fifo_13_tlast(m_axis_fifo_13_tlast),
        .m_axis_fifo_13_tvalid(m_axis_fifo_13_tvalid),
        .m_axis_fifo_13_tkeep(m_axis_fifo_13_tkeep),
        .m_axis_fifo_13_tstrb(m_axis_fifo_13_tstrb),
        .m_axis_fifo_13_tdata(m_axis_fifo_13_tdata),
        .m_axis_fifo_13_tready(m_axis_fifo_13_tready),
        .ap_fifo_oarg_13_full_n(ap_fifo_oarg_13_full_n),
        .ap_fifo_oarg_13_din(ap_fifo_oarg_13_din),
        .ap_fifo_oarg_13_write(ap_fifo_oarg_13_write),
        .m_axis_fifo_14_aclk(m_axis_fifo_14_aclk),
        .m_axis_fifo_14_aresetn(m_axis_fifo_14_aresetn),
        .m_axis_fifo_14_tlast(m_axis_fifo_14_tlast),
        .m_axis_fifo_14_tvalid(m_axis_fifo_14_tvalid),
        .m_axis_fifo_14_tkeep(m_axis_fifo_14_tkeep),
        .m_axis_fifo_14_tstrb(m_axis_fifo_14_tstrb),
        .m_axis_fifo_14_tdata(m_axis_fifo_14_tdata),
        .m_axis_fifo_14_tready(m_axis_fifo_14_tready),
        .ap_fifo_oarg_14_full_n(ap_fifo_oarg_14_full_n),
        .ap_fifo_oarg_14_din(ap_fifo_oarg_14_din),
        .ap_fifo_oarg_14_write(ap_fifo_oarg_14_write),
        .m_axis_fifo_15_aclk(m_axis_fifo_15_aclk),
        .m_axis_fifo_15_aresetn(m_axis_fifo_15_aresetn),
        .m_axis_fifo_15_tlast(m_axis_fifo_15_tlast),
        .m_axis_fifo_15_tvalid(m_axis_fifo_15_tvalid),
        .m_axis_fifo_15_tkeep(m_axis_fifo_15_tkeep),
        .m_axis_fifo_15_tstrb(m_axis_fifo_15_tstrb),
        .m_axis_fifo_15_tdata(m_axis_fifo_15_tdata),
        .m_axis_fifo_15_tready(m_axis_fifo_15_tready),
        .ap_fifo_oarg_15_full_n(ap_fifo_oarg_15_full_n),
        .ap_fifo_oarg_15_din(ap_fifo_oarg_15_din),
        .ap_fifo_oarg_15_write(ap_fifo_oarg_15_write),
        .m_axis_fifo_16_aclk(m_axis_fifo_16_aclk),
        .m_axis_fifo_16_aresetn(m_axis_fifo_16_aresetn),
        .m_axis_fifo_16_tlast(m_axis_fifo_16_tlast),
        .m_axis_fifo_16_tvalid(m_axis_fifo_16_tvalid),
        .m_axis_fifo_16_tkeep(m_axis_fifo_16_tkeep),
        .m_axis_fifo_16_tstrb(m_axis_fifo_16_tstrb),
        .m_axis_fifo_16_tdata(m_axis_fifo_16_tdata),
        .m_axis_fifo_16_tready(m_axis_fifo_16_tready),
        .ap_fifo_oarg_16_full_n(ap_fifo_oarg_16_full_n),
        .ap_fifo_oarg_16_din(ap_fifo_oarg_16_din),
        .ap_fifo_oarg_16_write(ap_fifo_oarg_16_write),
        .m_axis_fifo_17_aclk(m_axis_fifo_17_aclk),
        .m_axis_fifo_17_aresetn(m_axis_fifo_17_aresetn),
        .m_axis_fifo_17_tlast(m_axis_fifo_17_tlast),
        .m_axis_fifo_17_tvalid(m_axis_fifo_17_tvalid),
        .m_axis_fifo_17_tkeep(m_axis_fifo_17_tkeep),
        .m_axis_fifo_17_tstrb(m_axis_fifo_17_tstrb),
        .m_axis_fifo_17_tdata(m_axis_fifo_17_tdata),
        .m_axis_fifo_17_tready(m_axis_fifo_17_tready),
        .ap_fifo_oarg_17_full_n(ap_fifo_oarg_17_full_n),
        .ap_fifo_oarg_17_din(ap_fifo_oarg_17_din),
        .ap_fifo_oarg_17_write(ap_fifo_oarg_17_write),
        .m_axis_fifo_18_aclk(m_axis_fifo_18_aclk),
        .m_axis_fifo_18_aresetn(m_axis_fifo_18_aresetn),
        .m_axis_fifo_18_tlast(m_axis_fifo_18_tlast),
        .m_axis_fifo_18_tvalid(m_axis_fifo_18_tvalid),
        .m_axis_fifo_18_tkeep(m_axis_fifo_18_tkeep),
        .m_axis_fifo_18_tstrb(m_axis_fifo_18_tstrb),
        .m_axis_fifo_18_tdata(m_axis_fifo_18_tdata),
        .m_axis_fifo_18_tready(m_axis_fifo_18_tready),
        .ap_fifo_oarg_18_full_n(ap_fifo_oarg_18_full_n),
        .ap_fifo_oarg_18_din(ap_fifo_oarg_18_din),
        .ap_fifo_oarg_18_write(ap_fifo_oarg_18_write),
        .m_axis_fifo_19_aclk(m_axis_fifo_19_aclk),
        .m_axis_fifo_19_aresetn(m_axis_fifo_19_aresetn),
        .m_axis_fifo_19_tlast(m_axis_fifo_19_tlast),
        .m_axis_fifo_19_tvalid(m_axis_fifo_19_tvalid),
        .m_axis_fifo_19_tkeep(m_axis_fifo_19_tkeep),
        .m_axis_fifo_19_tstrb(m_axis_fifo_19_tstrb),
        .m_axis_fifo_19_tdata(m_axis_fifo_19_tdata),
        .m_axis_fifo_19_tready(m_axis_fifo_19_tready),
        .ap_fifo_oarg_19_full_n(ap_fifo_oarg_19_full_n),
        .ap_fifo_oarg_19_din(ap_fifo_oarg_19_din),
        .ap_fifo_oarg_19_write(ap_fifo_oarg_19_write),
        .m_axis_fifo_20_aclk(m_axis_fifo_20_aclk),
        .m_axis_fifo_20_aresetn(m_axis_fifo_20_aresetn),
        .m_axis_fifo_20_tlast(m_axis_fifo_20_tlast),
        .m_axis_fifo_20_tvalid(m_axis_fifo_20_tvalid),
        .m_axis_fifo_20_tkeep(m_axis_fifo_20_tkeep),
        .m_axis_fifo_20_tstrb(m_axis_fifo_20_tstrb),
        .m_axis_fifo_20_tdata(m_axis_fifo_20_tdata),
        .m_axis_fifo_20_tready(m_axis_fifo_20_tready),
        .ap_fifo_oarg_20_full_n(ap_fifo_oarg_20_full_n),
        .ap_fifo_oarg_20_din(ap_fifo_oarg_20_din),
        .ap_fifo_oarg_20_write(ap_fifo_oarg_20_write),
        .m_axis_fifo_21_aclk(m_axis_fifo_21_aclk),
        .m_axis_fifo_21_aresetn(m_axis_fifo_21_aresetn),
        .m_axis_fifo_21_tlast(m_axis_fifo_21_tlast),
        .m_axis_fifo_21_tvalid(m_axis_fifo_21_tvalid),
        .m_axis_fifo_21_tkeep(m_axis_fifo_21_tkeep),
        .m_axis_fifo_21_tstrb(m_axis_fifo_21_tstrb),
        .m_axis_fifo_21_tdata(m_axis_fifo_21_tdata),
        .m_axis_fifo_21_tready(m_axis_fifo_21_tready),
        .ap_fifo_oarg_21_full_n(ap_fifo_oarg_21_full_n),
        .ap_fifo_oarg_21_din(ap_fifo_oarg_21_din),
        .ap_fifo_oarg_21_write(ap_fifo_oarg_21_write),
        .m_axis_fifo_22_aclk(m_axis_fifo_22_aclk),
        .m_axis_fifo_22_aresetn(m_axis_fifo_22_aresetn),
        .m_axis_fifo_22_tlast(m_axis_fifo_22_tlast),
        .m_axis_fifo_22_tvalid(m_axis_fifo_22_tvalid),
        .m_axis_fifo_22_tkeep(m_axis_fifo_22_tkeep),
        .m_axis_fifo_22_tstrb(m_axis_fifo_22_tstrb),
        .m_axis_fifo_22_tdata(m_axis_fifo_22_tdata),
        .m_axis_fifo_22_tready(m_axis_fifo_22_tready),
        .ap_fifo_oarg_22_full_n(ap_fifo_oarg_22_full_n),
        .ap_fifo_oarg_22_din(ap_fifo_oarg_22_din),
        .ap_fifo_oarg_22_write(ap_fifo_oarg_22_write),
        .m_axis_fifo_23_aclk(m_axis_fifo_23_aclk),
        .m_axis_fifo_23_aresetn(m_axis_fifo_23_aresetn),
        .m_axis_fifo_23_tlast(m_axis_fifo_23_tlast),
        .m_axis_fifo_23_tvalid(m_axis_fifo_23_tvalid),
        .m_axis_fifo_23_tkeep(m_axis_fifo_23_tkeep),
        .m_axis_fifo_23_tstrb(m_axis_fifo_23_tstrb),
        .m_axis_fifo_23_tdata(m_axis_fifo_23_tdata),
        .m_axis_fifo_23_tready(m_axis_fifo_23_tready),
        .ap_fifo_oarg_23_full_n(ap_fifo_oarg_23_full_n),
        .ap_fifo_oarg_23_din(ap_fifo_oarg_23_din),
        .ap_fifo_oarg_23_write(ap_fifo_oarg_23_write),
        .m_axis_fifo_24_aclk(m_axis_fifo_24_aclk),
        .m_axis_fifo_24_aresetn(m_axis_fifo_24_aresetn),
        .m_axis_fifo_24_tlast(m_axis_fifo_24_tlast),
        .m_axis_fifo_24_tvalid(m_axis_fifo_24_tvalid),
        .m_axis_fifo_24_tkeep(m_axis_fifo_24_tkeep),
        .m_axis_fifo_24_tstrb(m_axis_fifo_24_tstrb),
        .m_axis_fifo_24_tdata(m_axis_fifo_24_tdata),
        .m_axis_fifo_24_tready(m_axis_fifo_24_tready),
        .ap_fifo_oarg_24_full_n(ap_fifo_oarg_24_full_n),
        .ap_fifo_oarg_24_din(ap_fifo_oarg_24_din),
        .ap_fifo_oarg_24_write(ap_fifo_oarg_24_write),
        .m_axis_fifo_25_aclk(m_axis_fifo_25_aclk),
        .m_axis_fifo_25_aresetn(m_axis_fifo_25_aresetn),
        .m_axis_fifo_25_tlast(m_axis_fifo_25_tlast),
        .m_axis_fifo_25_tvalid(m_axis_fifo_25_tvalid),
        .m_axis_fifo_25_tkeep(m_axis_fifo_25_tkeep),
        .m_axis_fifo_25_tstrb(m_axis_fifo_25_tstrb),
        .m_axis_fifo_25_tdata(m_axis_fifo_25_tdata),
        .m_axis_fifo_25_tready(m_axis_fifo_25_tready),
        .ap_fifo_oarg_25_full_n(ap_fifo_oarg_25_full_n),
        .ap_fifo_oarg_25_din(ap_fifo_oarg_25_din),
        .ap_fifo_oarg_25_write(ap_fifo_oarg_25_write),
        .m_axis_fifo_26_aclk(m_axis_fifo_26_aclk),
        .m_axis_fifo_26_aresetn(m_axis_fifo_26_aresetn),
        .m_axis_fifo_26_tlast(m_axis_fifo_26_tlast),
        .m_axis_fifo_26_tvalid(m_axis_fifo_26_tvalid),
        .m_axis_fifo_26_tkeep(m_axis_fifo_26_tkeep),
        .m_axis_fifo_26_tstrb(m_axis_fifo_26_tstrb),
        .m_axis_fifo_26_tdata(m_axis_fifo_26_tdata),
        .m_axis_fifo_26_tready(m_axis_fifo_26_tready),
        .ap_fifo_oarg_26_full_n(ap_fifo_oarg_26_full_n),
        .ap_fifo_oarg_26_din(ap_fifo_oarg_26_din),
        .ap_fifo_oarg_26_write(ap_fifo_oarg_26_write),
        .m_axis_fifo_27_aclk(m_axis_fifo_27_aclk),
        .m_axis_fifo_27_aresetn(m_axis_fifo_27_aresetn),
        .m_axis_fifo_27_tlast(m_axis_fifo_27_tlast),
        .m_axis_fifo_27_tvalid(m_axis_fifo_27_tvalid),
        .m_axis_fifo_27_tkeep(m_axis_fifo_27_tkeep),
        .m_axis_fifo_27_tstrb(m_axis_fifo_27_tstrb),
        .m_axis_fifo_27_tdata(m_axis_fifo_27_tdata),
        .m_axis_fifo_27_tready(m_axis_fifo_27_tready),
        .ap_fifo_oarg_27_full_n(ap_fifo_oarg_27_full_n),
        .ap_fifo_oarg_27_din(ap_fifo_oarg_27_din),
        .ap_fifo_oarg_27_write(ap_fifo_oarg_27_write),
        .m_axis_fifo_28_aclk(m_axis_fifo_28_aclk),
        .m_axis_fifo_28_aresetn(m_axis_fifo_28_aresetn),
        .m_axis_fifo_28_tlast(m_axis_fifo_28_tlast),
        .m_axis_fifo_28_tvalid(m_axis_fifo_28_tvalid),
        .m_axis_fifo_28_tkeep(m_axis_fifo_28_tkeep),
        .m_axis_fifo_28_tstrb(m_axis_fifo_28_tstrb),
        .m_axis_fifo_28_tdata(m_axis_fifo_28_tdata),
        .m_axis_fifo_28_tready(m_axis_fifo_28_tready),
        .ap_fifo_oarg_28_full_n(ap_fifo_oarg_28_full_n),
        .ap_fifo_oarg_28_din(ap_fifo_oarg_28_din),
        .ap_fifo_oarg_28_write(ap_fifo_oarg_28_write),
        .m_axis_fifo_29_aclk(m_axis_fifo_29_aclk),
        .m_axis_fifo_29_aresetn(m_axis_fifo_29_aresetn),
        .m_axis_fifo_29_tlast(m_axis_fifo_29_tlast),
        .m_axis_fifo_29_tvalid(m_axis_fifo_29_tvalid),
        .m_axis_fifo_29_tkeep(m_axis_fifo_29_tkeep),
        .m_axis_fifo_29_tstrb(m_axis_fifo_29_tstrb),
        .m_axis_fifo_29_tdata(m_axis_fifo_29_tdata),
        .m_axis_fifo_29_tready(m_axis_fifo_29_tready),
        .ap_fifo_oarg_29_full_n(ap_fifo_oarg_29_full_n),
        .ap_fifo_oarg_29_din(ap_fifo_oarg_29_din),
        .ap_fifo_oarg_29_write(ap_fifo_oarg_29_write),
        .m_axis_fifo_30_aclk(m_axis_fifo_30_aclk),
        .m_axis_fifo_30_aresetn(m_axis_fifo_30_aresetn),
        .m_axis_fifo_30_tlast(m_axis_fifo_30_tlast),
        .m_axis_fifo_30_tvalid(m_axis_fifo_30_tvalid),
        .m_axis_fifo_30_tkeep(m_axis_fifo_30_tkeep),
        .m_axis_fifo_30_tstrb(m_axis_fifo_30_tstrb),
        .m_axis_fifo_30_tdata(m_axis_fifo_30_tdata),
        .m_axis_fifo_30_tready(m_axis_fifo_30_tready),
        .ap_fifo_oarg_30_full_n(ap_fifo_oarg_30_full_n),
        .ap_fifo_oarg_30_din(ap_fifo_oarg_30_din),
        .ap_fifo_oarg_30_write(ap_fifo_oarg_30_write),
        .m_axis_fifo_31_aclk(m_axis_fifo_31_aclk),
        .m_axis_fifo_31_aresetn(m_axis_fifo_31_aresetn),
        .m_axis_fifo_31_tlast(m_axis_fifo_31_tlast),
        .m_axis_fifo_31_tvalid(m_axis_fifo_31_tvalid),
        .m_axis_fifo_31_tkeep(m_axis_fifo_31_tkeep),
        .m_axis_fifo_31_tstrb(m_axis_fifo_31_tstrb),
        .m_axis_fifo_31_tdata(m_axis_fifo_31_tdata),
        .m_axis_fifo_31_tready(m_axis_fifo_31_tready),
        .ap_fifo_oarg_31_full_n(ap_fifo_oarg_31_full_n),
        .ap_fifo_oarg_31_din(ap_fifo_oarg_31_din),
        .ap_fifo_oarg_31_write(ap_fifo_oarg_31_write),
        .m_axis_fifo_32_aclk(m_axis_fifo_32_aclk),
        .m_axis_fifo_32_aresetn(m_axis_fifo_32_aresetn),
        .m_axis_fifo_32_tlast(m_axis_fifo_32_tlast),
        .m_axis_fifo_32_tvalid(m_axis_fifo_32_tvalid),
        .m_axis_fifo_32_tkeep(m_axis_fifo_32_tkeep),
        .m_axis_fifo_32_tstrb(m_axis_fifo_32_tstrb),
        .m_axis_fifo_32_tdata(m_axis_fifo_32_tdata),
        .m_axis_fifo_32_tready(m_axis_fifo_32_tready),
        .ap_fifo_oarg_32_full_n(ap_fifo_oarg_32_full_n),
        .ap_fifo_oarg_32_din(ap_fifo_oarg_32_din),
        .ap_fifo_oarg_32_write(ap_fifo_oarg_32_write),
        .m_axis_fifo_33_aclk(m_axis_fifo_33_aclk),
        .m_axis_fifo_33_aresetn(m_axis_fifo_33_aresetn),
        .m_axis_fifo_33_tlast(m_axis_fifo_33_tlast),
        .m_axis_fifo_33_tvalid(m_axis_fifo_33_tvalid),
        .m_axis_fifo_33_tkeep(m_axis_fifo_33_tkeep),
        .m_axis_fifo_33_tstrb(m_axis_fifo_33_tstrb),
        .m_axis_fifo_33_tdata(m_axis_fifo_33_tdata),
        .m_axis_fifo_33_tready(m_axis_fifo_33_tready),
        .ap_fifo_oarg_33_full_n(ap_fifo_oarg_33_full_n),
        .ap_fifo_oarg_33_din(ap_fifo_oarg_33_din),
        .ap_fifo_oarg_33_write(ap_fifo_oarg_33_write),
        .m_axis_fifo_34_aclk(m_axis_fifo_34_aclk),
        .m_axis_fifo_34_aresetn(m_axis_fifo_34_aresetn),
        .m_axis_fifo_34_tlast(m_axis_fifo_34_tlast),
        .m_axis_fifo_34_tvalid(m_axis_fifo_34_tvalid),
        .m_axis_fifo_34_tkeep(m_axis_fifo_34_tkeep),
        .m_axis_fifo_34_tstrb(m_axis_fifo_34_tstrb),
        .m_axis_fifo_34_tdata(m_axis_fifo_34_tdata),
        .m_axis_fifo_34_tready(m_axis_fifo_34_tready),
        .ap_fifo_oarg_34_full_n(ap_fifo_oarg_34_full_n),
        .ap_fifo_oarg_34_din(ap_fifo_oarg_34_din),
        .ap_fifo_oarg_34_write(ap_fifo_oarg_34_write),
        .m_axis_fifo_35_aclk(m_axis_fifo_35_aclk),
        .m_axis_fifo_35_aresetn(m_axis_fifo_35_aresetn),
        .m_axis_fifo_35_tlast(m_axis_fifo_35_tlast),
        .m_axis_fifo_35_tvalid(m_axis_fifo_35_tvalid),
        .m_axis_fifo_35_tkeep(m_axis_fifo_35_tkeep),
        .m_axis_fifo_35_tstrb(m_axis_fifo_35_tstrb),
        .m_axis_fifo_35_tdata(m_axis_fifo_35_tdata),
        .m_axis_fifo_35_tready(m_axis_fifo_35_tready),
        .ap_fifo_oarg_35_full_n(ap_fifo_oarg_35_full_n),
        .ap_fifo_oarg_35_din(ap_fifo_oarg_35_din),
        .ap_fifo_oarg_35_write(ap_fifo_oarg_35_write),
        .m_axis_fifo_36_aclk(m_axis_fifo_36_aclk),
        .m_axis_fifo_36_aresetn(m_axis_fifo_36_aresetn),
        .m_axis_fifo_36_tlast(m_axis_fifo_36_tlast),
        .m_axis_fifo_36_tvalid(m_axis_fifo_36_tvalid),
        .m_axis_fifo_36_tkeep(m_axis_fifo_36_tkeep),
        .m_axis_fifo_36_tstrb(m_axis_fifo_36_tstrb),
        .m_axis_fifo_36_tdata(m_axis_fifo_36_tdata),
        .m_axis_fifo_36_tready(m_axis_fifo_36_tready),
        .ap_fifo_oarg_36_full_n(ap_fifo_oarg_36_full_n),
        .ap_fifo_oarg_36_din(ap_fifo_oarg_36_din),
        .ap_fifo_oarg_36_write(ap_fifo_oarg_36_write),
        .m_axis_fifo_37_aclk(m_axis_fifo_37_aclk),
        .m_axis_fifo_37_aresetn(m_axis_fifo_37_aresetn),
        .m_axis_fifo_37_tlast(m_axis_fifo_37_tlast),
        .m_axis_fifo_37_tvalid(m_axis_fifo_37_tvalid),
        .m_axis_fifo_37_tkeep(m_axis_fifo_37_tkeep),
        .m_axis_fifo_37_tstrb(m_axis_fifo_37_tstrb),
        .m_axis_fifo_37_tdata(m_axis_fifo_37_tdata),
        .m_axis_fifo_37_tready(m_axis_fifo_37_tready),
        .ap_fifo_oarg_37_full_n(ap_fifo_oarg_37_full_n),
        .ap_fifo_oarg_37_din(ap_fifo_oarg_37_din),
        .ap_fifo_oarg_37_write(ap_fifo_oarg_37_write),
        .m_axis_fifo_38_aclk(m_axis_fifo_38_aclk),
        .m_axis_fifo_38_aresetn(m_axis_fifo_38_aresetn),
        .m_axis_fifo_38_tlast(m_axis_fifo_38_tlast),
        .m_axis_fifo_38_tvalid(m_axis_fifo_38_tvalid),
        .m_axis_fifo_38_tkeep(m_axis_fifo_38_tkeep),
        .m_axis_fifo_38_tstrb(m_axis_fifo_38_tstrb),
        .m_axis_fifo_38_tdata(m_axis_fifo_38_tdata),
        .m_axis_fifo_38_tready(m_axis_fifo_38_tready),
        .ap_fifo_oarg_38_full_n(ap_fifo_oarg_38_full_n),
        .ap_fifo_oarg_38_din(ap_fifo_oarg_38_din),
        .ap_fifo_oarg_38_write(ap_fifo_oarg_38_write),
        .m_axis_fifo_39_aclk(m_axis_fifo_39_aclk),
        .m_axis_fifo_39_aresetn(m_axis_fifo_39_aresetn),
        .m_axis_fifo_39_tlast(m_axis_fifo_39_tlast),
        .m_axis_fifo_39_tvalid(m_axis_fifo_39_tvalid),
        .m_axis_fifo_39_tkeep(m_axis_fifo_39_tkeep),
        .m_axis_fifo_39_tstrb(m_axis_fifo_39_tstrb),
        .m_axis_fifo_39_tdata(m_axis_fifo_39_tdata),
        .m_axis_fifo_39_tready(m_axis_fifo_39_tready),
        .ap_fifo_oarg_39_full_n(ap_fifo_oarg_39_full_n),
        .ap_fifo_oarg_39_din(ap_fifo_oarg_39_din),
        .ap_fifo_oarg_39_write(ap_fifo_oarg_39_write),
        .m_axis_fifo_40_aclk(m_axis_fifo_40_aclk),
        .m_axis_fifo_40_aresetn(m_axis_fifo_40_aresetn),
        .m_axis_fifo_40_tlast(m_axis_fifo_40_tlast),
        .m_axis_fifo_40_tvalid(m_axis_fifo_40_tvalid),
        .m_axis_fifo_40_tkeep(m_axis_fifo_40_tkeep),
        .m_axis_fifo_40_tstrb(m_axis_fifo_40_tstrb),
        .m_axis_fifo_40_tdata(m_axis_fifo_40_tdata),
        .m_axis_fifo_40_tready(m_axis_fifo_40_tready),
        .ap_fifo_oarg_40_full_n(ap_fifo_oarg_40_full_n),
        .ap_fifo_oarg_40_din(ap_fifo_oarg_40_din),
        .ap_fifo_oarg_40_write(ap_fifo_oarg_40_write),
        .m_axis_fifo_41_aclk(m_axis_fifo_41_aclk),
        .m_axis_fifo_41_aresetn(m_axis_fifo_41_aresetn),
        .m_axis_fifo_41_tlast(m_axis_fifo_41_tlast),
        .m_axis_fifo_41_tvalid(m_axis_fifo_41_tvalid),
        .m_axis_fifo_41_tkeep(m_axis_fifo_41_tkeep),
        .m_axis_fifo_41_tstrb(m_axis_fifo_41_tstrb),
        .m_axis_fifo_41_tdata(m_axis_fifo_41_tdata),
        .m_axis_fifo_41_tready(m_axis_fifo_41_tready),
        .ap_fifo_oarg_41_full_n(ap_fifo_oarg_41_full_n),
        .ap_fifo_oarg_41_din(ap_fifo_oarg_41_din),
        .ap_fifo_oarg_41_write(ap_fifo_oarg_41_write),
        .m_axis_fifo_42_aclk(m_axis_fifo_42_aclk),
        .m_axis_fifo_42_aresetn(m_axis_fifo_42_aresetn),
        .m_axis_fifo_42_tlast(m_axis_fifo_42_tlast),
        .m_axis_fifo_42_tvalid(m_axis_fifo_42_tvalid),
        .m_axis_fifo_42_tkeep(m_axis_fifo_42_tkeep),
        .m_axis_fifo_42_tstrb(m_axis_fifo_42_tstrb),
        .m_axis_fifo_42_tdata(m_axis_fifo_42_tdata),
        .m_axis_fifo_42_tready(m_axis_fifo_42_tready),
        .ap_fifo_oarg_42_full_n(ap_fifo_oarg_42_full_n),
        .ap_fifo_oarg_42_din(ap_fifo_oarg_42_din),
        .ap_fifo_oarg_42_write(ap_fifo_oarg_42_write),
        .m_axis_fifo_43_aclk(m_axis_fifo_43_aclk),
        .m_axis_fifo_43_aresetn(m_axis_fifo_43_aresetn),
        .m_axis_fifo_43_tlast(m_axis_fifo_43_tlast),
        .m_axis_fifo_43_tvalid(m_axis_fifo_43_tvalid),
        .m_axis_fifo_43_tkeep(m_axis_fifo_43_tkeep),
        .m_axis_fifo_43_tstrb(m_axis_fifo_43_tstrb),
        .m_axis_fifo_43_tdata(m_axis_fifo_43_tdata),
        .m_axis_fifo_43_tready(m_axis_fifo_43_tready),
        .ap_fifo_oarg_43_full_n(ap_fifo_oarg_43_full_n),
        .ap_fifo_oarg_43_din(ap_fifo_oarg_43_din),
        .ap_fifo_oarg_43_write(ap_fifo_oarg_43_write),
        .m_axis_fifo_44_aclk(m_axis_fifo_44_aclk),
        .m_axis_fifo_44_aresetn(m_axis_fifo_44_aresetn),
        .m_axis_fifo_44_tlast(m_axis_fifo_44_tlast),
        .m_axis_fifo_44_tvalid(m_axis_fifo_44_tvalid),
        .m_axis_fifo_44_tkeep(m_axis_fifo_44_tkeep),
        .m_axis_fifo_44_tstrb(m_axis_fifo_44_tstrb),
        .m_axis_fifo_44_tdata(m_axis_fifo_44_tdata),
        .m_axis_fifo_44_tready(m_axis_fifo_44_tready),
        .ap_fifo_oarg_44_full_n(ap_fifo_oarg_44_full_n),
        .ap_fifo_oarg_44_din(ap_fifo_oarg_44_din),
        .ap_fifo_oarg_44_write(ap_fifo_oarg_44_write),
        .m_axis_fifo_45_aclk(m_axis_fifo_45_aclk),
        .m_axis_fifo_45_aresetn(m_axis_fifo_45_aresetn),
        .m_axis_fifo_45_tlast(m_axis_fifo_45_tlast),
        .m_axis_fifo_45_tvalid(m_axis_fifo_45_tvalid),
        .m_axis_fifo_45_tkeep(m_axis_fifo_45_tkeep),
        .m_axis_fifo_45_tstrb(m_axis_fifo_45_tstrb),
        .m_axis_fifo_45_tdata(m_axis_fifo_45_tdata),
        .m_axis_fifo_45_tready(m_axis_fifo_45_tready),
        .ap_fifo_oarg_45_full_n(ap_fifo_oarg_45_full_n),
        .ap_fifo_oarg_45_din(ap_fifo_oarg_45_din),
        .ap_fifo_oarg_45_write(ap_fifo_oarg_45_write),
        .m_axis_fifo_46_aclk(m_axis_fifo_46_aclk),
        .m_axis_fifo_46_aresetn(m_axis_fifo_46_aresetn),
        .m_axis_fifo_46_tlast(m_axis_fifo_46_tlast),
        .m_axis_fifo_46_tvalid(m_axis_fifo_46_tvalid),
        .m_axis_fifo_46_tkeep(m_axis_fifo_46_tkeep),
        .m_axis_fifo_46_tstrb(m_axis_fifo_46_tstrb),
        .m_axis_fifo_46_tdata(m_axis_fifo_46_tdata),
        .m_axis_fifo_46_tready(m_axis_fifo_46_tready),
        .ap_fifo_oarg_46_full_n(ap_fifo_oarg_46_full_n),
        .ap_fifo_oarg_46_din(ap_fifo_oarg_46_din),
        .ap_fifo_oarg_46_write(ap_fifo_oarg_46_write),
        .m_axis_fifo_47_aclk(m_axis_fifo_47_aclk),
        .m_axis_fifo_47_aresetn(m_axis_fifo_47_aresetn),
        .m_axis_fifo_47_tlast(m_axis_fifo_47_tlast),
        .m_axis_fifo_47_tvalid(m_axis_fifo_47_tvalid),
        .m_axis_fifo_47_tkeep(m_axis_fifo_47_tkeep),
        .m_axis_fifo_47_tstrb(m_axis_fifo_47_tstrb),
        .m_axis_fifo_47_tdata(m_axis_fifo_47_tdata),
        .m_axis_fifo_47_tready(m_axis_fifo_47_tready),
        .ap_fifo_oarg_47_full_n(ap_fifo_oarg_47_full_n),
        .ap_fifo_oarg_47_din(ap_fifo_oarg_47_din),
        .ap_fifo_oarg_47_write(ap_fifo_oarg_47_write),
        .m_axis_fifo_48_aclk(m_axis_fifo_48_aclk),
        .m_axis_fifo_48_aresetn(m_axis_fifo_48_aresetn),
        .m_axis_fifo_48_tlast(m_axis_fifo_48_tlast),
        .m_axis_fifo_48_tvalid(m_axis_fifo_48_tvalid),
        .m_axis_fifo_48_tkeep(m_axis_fifo_48_tkeep),
        .m_axis_fifo_48_tstrb(m_axis_fifo_48_tstrb),
        .m_axis_fifo_48_tdata(m_axis_fifo_48_tdata),
        .m_axis_fifo_48_tready(m_axis_fifo_48_tready),
        .ap_fifo_oarg_48_full_n(ap_fifo_oarg_48_full_n),
        .ap_fifo_oarg_48_din(ap_fifo_oarg_48_din),
        .ap_fifo_oarg_48_write(ap_fifo_oarg_48_write),
        .m_axis_fifo_49_aclk(m_axis_fifo_49_aclk),
        .m_axis_fifo_49_aresetn(m_axis_fifo_49_aresetn),
        .m_axis_fifo_49_tlast(m_axis_fifo_49_tlast),
        .m_axis_fifo_49_tvalid(m_axis_fifo_49_tvalid),
        .m_axis_fifo_49_tkeep(m_axis_fifo_49_tkeep),
        .m_axis_fifo_49_tstrb(m_axis_fifo_49_tstrb),
        .m_axis_fifo_49_tdata(m_axis_fifo_49_tdata),
        .m_axis_fifo_49_tready(m_axis_fifo_49_tready),
        .ap_fifo_oarg_49_full_n(ap_fifo_oarg_49_full_n),
        .ap_fifo_oarg_49_din(ap_fifo_oarg_49_din),
        .ap_fifo_oarg_49_write(ap_fifo_oarg_49_write),
        .m_axis_fifo_50_aclk(m_axis_fifo_50_aclk),
        .m_axis_fifo_50_aresetn(m_axis_fifo_50_aresetn),
        .m_axis_fifo_50_tlast(m_axis_fifo_50_tlast),
        .m_axis_fifo_50_tvalid(m_axis_fifo_50_tvalid),
        .m_axis_fifo_50_tkeep(m_axis_fifo_50_tkeep),
        .m_axis_fifo_50_tstrb(m_axis_fifo_50_tstrb),
        .m_axis_fifo_50_tdata(m_axis_fifo_50_tdata),
        .m_axis_fifo_50_tready(m_axis_fifo_50_tready),
        .ap_fifo_oarg_50_full_n(ap_fifo_oarg_50_full_n),
        .ap_fifo_oarg_50_din(ap_fifo_oarg_50_din),
        .ap_fifo_oarg_50_write(ap_fifo_oarg_50_write),
        .m_axis_fifo_51_aclk(m_axis_fifo_51_aclk),
        .m_axis_fifo_51_aresetn(m_axis_fifo_51_aresetn),
        .m_axis_fifo_51_tlast(m_axis_fifo_51_tlast),
        .m_axis_fifo_51_tvalid(m_axis_fifo_51_tvalid),
        .m_axis_fifo_51_tkeep(m_axis_fifo_51_tkeep),
        .m_axis_fifo_51_tstrb(m_axis_fifo_51_tstrb),
        .m_axis_fifo_51_tdata(m_axis_fifo_51_tdata),
        .m_axis_fifo_51_tready(m_axis_fifo_51_tready),
        .ap_fifo_oarg_51_full_n(ap_fifo_oarg_51_full_n),
        .ap_fifo_oarg_51_din(ap_fifo_oarg_51_din),
        .ap_fifo_oarg_51_write(ap_fifo_oarg_51_write),
        .m_axis_fifo_52_aclk(m_axis_fifo_52_aclk),
        .m_axis_fifo_52_aresetn(m_axis_fifo_52_aresetn),
        .m_axis_fifo_52_tlast(m_axis_fifo_52_tlast),
        .m_axis_fifo_52_tvalid(m_axis_fifo_52_tvalid),
        .m_axis_fifo_52_tkeep(m_axis_fifo_52_tkeep),
        .m_axis_fifo_52_tstrb(m_axis_fifo_52_tstrb),
        .m_axis_fifo_52_tdata(m_axis_fifo_52_tdata),
        .m_axis_fifo_52_tready(m_axis_fifo_52_tready),
        .ap_fifo_oarg_52_full_n(ap_fifo_oarg_52_full_n),
        .ap_fifo_oarg_52_din(ap_fifo_oarg_52_din),
        .ap_fifo_oarg_52_write(ap_fifo_oarg_52_write),
        .m_axis_fifo_53_aclk(m_axis_fifo_53_aclk),
        .m_axis_fifo_53_aresetn(m_axis_fifo_53_aresetn),
        .m_axis_fifo_53_tlast(m_axis_fifo_53_tlast),
        .m_axis_fifo_53_tvalid(m_axis_fifo_53_tvalid),
        .m_axis_fifo_53_tkeep(m_axis_fifo_53_tkeep),
        .m_axis_fifo_53_tstrb(m_axis_fifo_53_tstrb),
        .m_axis_fifo_53_tdata(m_axis_fifo_53_tdata),
        .m_axis_fifo_53_tready(m_axis_fifo_53_tready),
        .ap_fifo_oarg_53_full_n(ap_fifo_oarg_53_full_n),
        .ap_fifo_oarg_53_din(ap_fifo_oarg_53_din),
        .ap_fifo_oarg_53_write(ap_fifo_oarg_53_write),
        .m_axis_fifo_54_aclk(m_axis_fifo_54_aclk),
        .m_axis_fifo_54_aresetn(m_axis_fifo_54_aresetn),
        .m_axis_fifo_54_tlast(m_axis_fifo_54_tlast),
        .m_axis_fifo_54_tvalid(m_axis_fifo_54_tvalid),
        .m_axis_fifo_54_tkeep(m_axis_fifo_54_tkeep),
        .m_axis_fifo_54_tstrb(m_axis_fifo_54_tstrb),
        .m_axis_fifo_54_tdata(m_axis_fifo_54_tdata),
        .m_axis_fifo_54_tready(m_axis_fifo_54_tready),
        .ap_fifo_oarg_54_full_n(ap_fifo_oarg_54_full_n),
        .ap_fifo_oarg_54_din(ap_fifo_oarg_54_din),
        .ap_fifo_oarg_54_write(ap_fifo_oarg_54_write),
        .m_axis_fifo_55_aclk(m_axis_fifo_55_aclk),
        .m_axis_fifo_55_aresetn(m_axis_fifo_55_aresetn),
        .m_axis_fifo_55_tlast(m_axis_fifo_55_tlast),
        .m_axis_fifo_55_tvalid(m_axis_fifo_55_tvalid),
        .m_axis_fifo_55_tkeep(m_axis_fifo_55_tkeep),
        .m_axis_fifo_55_tstrb(m_axis_fifo_55_tstrb),
        .m_axis_fifo_55_tdata(m_axis_fifo_55_tdata),
        .m_axis_fifo_55_tready(m_axis_fifo_55_tready),
        .ap_fifo_oarg_55_full_n(ap_fifo_oarg_55_full_n),
        .ap_fifo_oarg_55_din(ap_fifo_oarg_55_din),
        .ap_fifo_oarg_55_write(ap_fifo_oarg_55_write),
        .m_axis_fifo_56_aclk(m_axis_fifo_56_aclk),
        .m_axis_fifo_56_aresetn(m_axis_fifo_56_aresetn),
        .m_axis_fifo_56_tlast(m_axis_fifo_56_tlast),
        .m_axis_fifo_56_tvalid(m_axis_fifo_56_tvalid),
        .m_axis_fifo_56_tkeep(m_axis_fifo_56_tkeep),
        .m_axis_fifo_56_tstrb(m_axis_fifo_56_tstrb),
        .m_axis_fifo_56_tdata(m_axis_fifo_56_tdata),
        .m_axis_fifo_56_tready(m_axis_fifo_56_tready),
        .ap_fifo_oarg_56_full_n(ap_fifo_oarg_56_full_n),
        .ap_fifo_oarg_56_din(ap_fifo_oarg_56_din),
        .ap_fifo_oarg_56_write(ap_fifo_oarg_56_write),
        .m_axis_fifo_57_aclk(m_axis_fifo_57_aclk),
        .m_axis_fifo_57_aresetn(m_axis_fifo_57_aresetn),
        .m_axis_fifo_57_tlast(m_axis_fifo_57_tlast),
        .m_axis_fifo_57_tvalid(m_axis_fifo_57_tvalid),
        .m_axis_fifo_57_tkeep(m_axis_fifo_57_tkeep),
        .m_axis_fifo_57_tstrb(m_axis_fifo_57_tstrb),
        .m_axis_fifo_57_tdata(m_axis_fifo_57_tdata),
        .m_axis_fifo_57_tready(m_axis_fifo_57_tready),
        .ap_fifo_oarg_57_full_n(ap_fifo_oarg_57_full_n),
        .ap_fifo_oarg_57_din(ap_fifo_oarg_57_din),
        .ap_fifo_oarg_57_write(ap_fifo_oarg_57_write),
        .m_axis_fifo_58_aclk(m_axis_fifo_58_aclk),
        .m_axis_fifo_58_aresetn(m_axis_fifo_58_aresetn),
        .m_axis_fifo_58_tlast(m_axis_fifo_58_tlast),
        .m_axis_fifo_58_tvalid(m_axis_fifo_58_tvalid),
        .m_axis_fifo_58_tkeep(m_axis_fifo_58_tkeep),
        .m_axis_fifo_58_tstrb(m_axis_fifo_58_tstrb),
        .m_axis_fifo_58_tdata(m_axis_fifo_58_tdata),
        .m_axis_fifo_58_tready(m_axis_fifo_58_tready),
        .ap_fifo_oarg_58_full_n(ap_fifo_oarg_58_full_n),
        .ap_fifo_oarg_58_din(ap_fifo_oarg_58_din),
        .ap_fifo_oarg_58_write(ap_fifo_oarg_58_write),
        .m_axis_fifo_59_aclk(m_axis_fifo_59_aclk),
        .m_axis_fifo_59_aresetn(m_axis_fifo_59_aresetn),
        .m_axis_fifo_59_tlast(m_axis_fifo_59_tlast),
        .m_axis_fifo_59_tvalid(m_axis_fifo_59_tvalid),
        .m_axis_fifo_59_tkeep(m_axis_fifo_59_tkeep),
        .m_axis_fifo_59_tstrb(m_axis_fifo_59_tstrb),
        .m_axis_fifo_59_tdata(m_axis_fifo_59_tdata),
        .m_axis_fifo_59_tready(m_axis_fifo_59_tready),
        .ap_fifo_oarg_59_full_n(ap_fifo_oarg_59_full_n),
        .ap_fifo_oarg_59_din(ap_fifo_oarg_59_din),
        .ap_fifo_oarg_59_write(ap_fifo_oarg_59_write),
        .m_axis_fifo_60_aclk(m_axis_fifo_60_aclk),
        .m_axis_fifo_60_aresetn(m_axis_fifo_60_aresetn),
        .m_axis_fifo_60_tlast(m_axis_fifo_60_tlast),
        .m_axis_fifo_60_tvalid(m_axis_fifo_60_tvalid),
        .m_axis_fifo_60_tkeep(m_axis_fifo_60_tkeep),
        .m_axis_fifo_60_tstrb(m_axis_fifo_60_tstrb),
        .m_axis_fifo_60_tdata(m_axis_fifo_60_tdata),
        .m_axis_fifo_60_tready(m_axis_fifo_60_tready),
        .ap_fifo_oarg_60_full_n(ap_fifo_oarg_60_full_n),
        .ap_fifo_oarg_60_din(ap_fifo_oarg_60_din),
        .ap_fifo_oarg_60_write(ap_fifo_oarg_60_write),
        .m_axis_fifo_61_aclk(m_axis_fifo_61_aclk),
        .m_axis_fifo_61_aresetn(m_axis_fifo_61_aresetn),
        .m_axis_fifo_61_tlast(m_axis_fifo_61_tlast),
        .m_axis_fifo_61_tvalid(m_axis_fifo_61_tvalid),
        .m_axis_fifo_61_tkeep(m_axis_fifo_61_tkeep),
        .m_axis_fifo_61_tstrb(m_axis_fifo_61_tstrb),
        .m_axis_fifo_61_tdata(m_axis_fifo_61_tdata),
        .m_axis_fifo_61_tready(m_axis_fifo_61_tready),
        .ap_fifo_oarg_61_full_n(ap_fifo_oarg_61_full_n),
        .ap_fifo_oarg_61_din(ap_fifo_oarg_61_din),
        .ap_fifo_oarg_61_write(ap_fifo_oarg_61_write),
        .m_axis_fifo_62_aclk(m_axis_fifo_62_aclk),
        .m_axis_fifo_62_aresetn(m_axis_fifo_62_aresetn),
        .m_axis_fifo_62_tlast(m_axis_fifo_62_tlast),
        .m_axis_fifo_62_tvalid(m_axis_fifo_62_tvalid),
        .m_axis_fifo_62_tkeep(m_axis_fifo_62_tkeep),
        .m_axis_fifo_62_tstrb(m_axis_fifo_62_tstrb),
        .m_axis_fifo_62_tdata(m_axis_fifo_62_tdata),
        .m_axis_fifo_62_tready(m_axis_fifo_62_tready),
        .ap_fifo_oarg_62_full_n(ap_fifo_oarg_62_full_n),
        .ap_fifo_oarg_62_din(ap_fifo_oarg_62_din),
        .ap_fifo_oarg_62_write(ap_fifo_oarg_62_write),
        .m_axis_fifo_63_aclk(m_axis_fifo_63_aclk),
        .m_axis_fifo_63_aresetn(m_axis_fifo_63_aresetn),
        .m_axis_fifo_63_tlast(m_axis_fifo_63_tlast),
        .m_axis_fifo_63_tvalid(m_axis_fifo_63_tvalid),
        .m_axis_fifo_63_tkeep(m_axis_fifo_63_tkeep),
        .m_axis_fifo_63_tstrb(m_axis_fifo_63_tstrb),
        .m_axis_fifo_63_tdata(m_axis_fifo_63_tdata),
        .m_axis_fifo_63_tready(m_axis_fifo_63_tready),
        .ap_fifo_oarg_63_full_n(ap_fifo_oarg_63_full_n),
        .ap_fifo_oarg_63_din(ap_fifo_oarg_63_din),
        .ap_fifo_oarg_63_write(ap_fifo_oarg_63_write),
        .m_axis_fifo_64_aclk(m_axis_fifo_64_aclk),
        .m_axis_fifo_64_aresetn(m_axis_fifo_64_aresetn),
        .m_axis_fifo_64_tlast(m_axis_fifo_64_tlast),
        .m_axis_fifo_64_tvalid(m_axis_fifo_64_tvalid),
        .m_axis_fifo_64_tkeep(m_axis_fifo_64_tkeep),
        .m_axis_fifo_64_tstrb(m_axis_fifo_64_tstrb),
        .m_axis_fifo_64_tdata(m_axis_fifo_64_tdata),
        .m_axis_fifo_64_tready(m_axis_fifo_64_tready),
        .ap_fifo_oarg_64_full_n(ap_fifo_oarg_64_full_n),
        .ap_fifo_oarg_64_din(ap_fifo_oarg_64_din),
        .ap_fifo_oarg_64_write(ap_fifo_oarg_64_write),
        .m_axis_fifo_65_aclk(m_axis_fifo_65_aclk),
        .m_axis_fifo_65_aresetn(m_axis_fifo_65_aresetn),
        .m_axis_fifo_65_tlast(m_axis_fifo_65_tlast),
        .m_axis_fifo_65_tvalid(m_axis_fifo_65_tvalid),
        .m_axis_fifo_65_tkeep(m_axis_fifo_65_tkeep),
        .m_axis_fifo_65_tstrb(m_axis_fifo_65_tstrb),
        .m_axis_fifo_65_tdata(m_axis_fifo_65_tdata),
        .m_axis_fifo_65_tready(m_axis_fifo_65_tready),
        .ap_fifo_oarg_65_full_n(ap_fifo_oarg_65_full_n),
        .ap_fifo_oarg_65_din(ap_fifo_oarg_65_din),
        .ap_fifo_oarg_65_write(ap_fifo_oarg_65_write),
        .m_axis_fifo_66_aclk(m_axis_fifo_66_aclk),
        .m_axis_fifo_66_aresetn(m_axis_fifo_66_aresetn),
        .m_axis_fifo_66_tlast(m_axis_fifo_66_tlast),
        .m_axis_fifo_66_tvalid(m_axis_fifo_66_tvalid),
        .m_axis_fifo_66_tkeep(m_axis_fifo_66_tkeep),
        .m_axis_fifo_66_tstrb(m_axis_fifo_66_tstrb),
        .m_axis_fifo_66_tdata(m_axis_fifo_66_tdata),
        .m_axis_fifo_66_tready(m_axis_fifo_66_tready),
        .ap_fifo_oarg_66_full_n(ap_fifo_oarg_66_full_n),
        .ap_fifo_oarg_66_din(ap_fifo_oarg_66_din),
        .ap_fifo_oarg_66_write(ap_fifo_oarg_66_write),
        .m_axis_fifo_67_aclk(m_axis_fifo_67_aclk),
        .m_axis_fifo_67_aresetn(m_axis_fifo_67_aresetn),
        .m_axis_fifo_67_tlast(m_axis_fifo_67_tlast),
        .m_axis_fifo_67_tvalid(m_axis_fifo_67_tvalid),
        .m_axis_fifo_67_tkeep(m_axis_fifo_67_tkeep),
        .m_axis_fifo_67_tstrb(m_axis_fifo_67_tstrb),
        .m_axis_fifo_67_tdata(m_axis_fifo_67_tdata),
        .m_axis_fifo_67_tready(m_axis_fifo_67_tready),
        .ap_fifo_oarg_67_full_n(ap_fifo_oarg_67_full_n),
        .ap_fifo_oarg_67_din(ap_fifo_oarg_67_din),
        .ap_fifo_oarg_67_write(ap_fifo_oarg_67_write),
        .m_axis_fifo_68_aclk(m_axis_fifo_68_aclk),
        .m_axis_fifo_68_aresetn(m_axis_fifo_68_aresetn),
        .m_axis_fifo_68_tlast(m_axis_fifo_68_tlast),
        .m_axis_fifo_68_tvalid(m_axis_fifo_68_tvalid),
        .m_axis_fifo_68_tkeep(m_axis_fifo_68_tkeep),
        .m_axis_fifo_68_tstrb(m_axis_fifo_68_tstrb),
        .m_axis_fifo_68_tdata(m_axis_fifo_68_tdata),
        .m_axis_fifo_68_tready(m_axis_fifo_68_tready),
        .ap_fifo_oarg_68_full_n(ap_fifo_oarg_68_full_n),
        .ap_fifo_oarg_68_din(ap_fifo_oarg_68_din),
        .ap_fifo_oarg_68_write(ap_fifo_oarg_68_write),
        .m_axis_fifo_69_aclk(m_axis_fifo_69_aclk),
        .m_axis_fifo_69_aresetn(m_axis_fifo_69_aresetn),
        .m_axis_fifo_69_tlast(m_axis_fifo_69_tlast),
        .m_axis_fifo_69_tvalid(m_axis_fifo_69_tvalid),
        .m_axis_fifo_69_tkeep(m_axis_fifo_69_tkeep),
        .m_axis_fifo_69_tstrb(m_axis_fifo_69_tstrb),
        .m_axis_fifo_69_tdata(m_axis_fifo_69_tdata),
        .m_axis_fifo_69_tready(m_axis_fifo_69_tready),
        .ap_fifo_oarg_69_full_n(ap_fifo_oarg_69_full_n),
        .ap_fifo_oarg_69_din(ap_fifo_oarg_69_din),
        .ap_fifo_oarg_69_write(ap_fifo_oarg_69_write),
        .m_axis_fifo_70_aclk(m_axis_fifo_70_aclk),
        .m_axis_fifo_70_aresetn(m_axis_fifo_70_aresetn),
        .m_axis_fifo_70_tlast(m_axis_fifo_70_tlast),
        .m_axis_fifo_70_tvalid(m_axis_fifo_70_tvalid),
        .m_axis_fifo_70_tkeep(m_axis_fifo_70_tkeep),
        .m_axis_fifo_70_tstrb(m_axis_fifo_70_tstrb),
        .m_axis_fifo_70_tdata(m_axis_fifo_70_tdata),
        .m_axis_fifo_70_tready(m_axis_fifo_70_tready),
        .ap_fifo_oarg_70_full_n(ap_fifo_oarg_70_full_n),
        .ap_fifo_oarg_70_din(ap_fifo_oarg_70_din),
        .ap_fifo_oarg_70_write(ap_fifo_oarg_70_write),
        .m_axis_fifo_71_aclk(m_axis_fifo_71_aclk),
        .m_axis_fifo_71_aresetn(m_axis_fifo_71_aresetn),
        .m_axis_fifo_71_tlast(m_axis_fifo_71_tlast),
        .m_axis_fifo_71_tvalid(m_axis_fifo_71_tvalid),
        .m_axis_fifo_71_tkeep(m_axis_fifo_71_tkeep),
        .m_axis_fifo_71_tstrb(m_axis_fifo_71_tstrb),
        .m_axis_fifo_71_tdata(m_axis_fifo_71_tdata),
        .m_axis_fifo_71_tready(m_axis_fifo_71_tready),
        .ap_fifo_oarg_71_full_n(ap_fifo_oarg_71_full_n),
        .ap_fifo_oarg_71_din(ap_fifo_oarg_71_din),
        .ap_fifo_oarg_71_write(ap_fifo_oarg_71_write),
        .m_axis_fifo_72_aclk(m_axis_fifo_72_aclk),
        .m_axis_fifo_72_aresetn(m_axis_fifo_72_aresetn),
        .m_axis_fifo_72_tlast(m_axis_fifo_72_tlast),
        .m_axis_fifo_72_tvalid(m_axis_fifo_72_tvalid),
        .m_axis_fifo_72_tkeep(m_axis_fifo_72_tkeep),
        .m_axis_fifo_72_tstrb(m_axis_fifo_72_tstrb),
        .m_axis_fifo_72_tdata(m_axis_fifo_72_tdata),
        .m_axis_fifo_72_tready(m_axis_fifo_72_tready),
        .ap_fifo_oarg_72_full_n(ap_fifo_oarg_72_full_n),
        .ap_fifo_oarg_72_din(ap_fifo_oarg_72_din),
        .ap_fifo_oarg_72_write(ap_fifo_oarg_72_write),
        .m_axis_fifo_73_aclk(m_axis_fifo_73_aclk),
        .m_axis_fifo_73_aresetn(m_axis_fifo_73_aresetn),
        .m_axis_fifo_73_tlast(m_axis_fifo_73_tlast),
        .m_axis_fifo_73_tvalid(m_axis_fifo_73_tvalid),
        .m_axis_fifo_73_tkeep(m_axis_fifo_73_tkeep),
        .m_axis_fifo_73_tstrb(m_axis_fifo_73_tstrb),
        .m_axis_fifo_73_tdata(m_axis_fifo_73_tdata),
        .m_axis_fifo_73_tready(m_axis_fifo_73_tready),
        .ap_fifo_oarg_73_full_n(ap_fifo_oarg_73_full_n),
        .ap_fifo_oarg_73_din(ap_fifo_oarg_73_din),
        .ap_fifo_oarg_73_write(ap_fifo_oarg_73_write),
        .m_axis_fifo_74_aclk(m_axis_fifo_74_aclk),
        .m_axis_fifo_74_aresetn(m_axis_fifo_74_aresetn),
        .m_axis_fifo_74_tlast(m_axis_fifo_74_tlast),
        .m_axis_fifo_74_tvalid(m_axis_fifo_74_tvalid),
        .m_axis_fifo_74_tkeep(m_axis_fifo_74_tkeep),
        .m_axis_fifo_74_tstrb(m_axis_fifo_74_tstrb),
        .m_axis_fifo_74_tdata(m_axis_fifo_74_tdata),
        .m_axis_fifo_74_tready(m_axis_fifo_74_tready),
        .ap_fifo_oarg_74_full_n(ap_fifo_oarg_74_full_n),
        .ap_fifo_oarg_74_din(ap_fifo_oarg_74_din),
        .ap_fifo_oarg_74_write(ap_fifo_oarg_74_write),
        .m_axis_fifo_75_aclk(m_axis_fifo_75_aclk),
        .m_axis_fifo_75_aresetn(m_axis_fifo_75_aresetn),
        .m_axis_fifo_75_tlast(m_axis_fifo_75_tlast),
        .m_axis_fifo_75_tvalid(m_axis_fifo_75_tvalid),
        .m_axis_fifo_75_tkeep(m_axis_fifo_75_tkeep),
        .m_axis_fifo_75_tstrb(m_axis_fifo_75_tstrb),
        .m_axis_fifo_75_tdata(m_axis_fifo_75_tdata),
        .m_axis_fifo_75_tready(m_axis_fifo_75_tready),
        .ap_fifo_oarg_75_full_n(ap_fifo_oarg_75_full_n),
        .ap_fifo_oarg_75_din(ap_fifo_oarg_75_din),
        .ap_fifo_oarg_75_write(ap_fifo_oarg_75_write),
        .m_axis_fifo_76_aclk(m_axis_fifo_76_aclk),
        .m_axis_fifo_76_aresetn(m_axis_fifo_76_aresetn),
        .m_axis_fifo_76_tlast(m_axis_fifo_76_tlast),
        .m_axis_fifo_76_tvalid(m_axis_fifo_76_tvalid),
        .m_axis_fifo_76_tkeep(m_axis_fifo_76_tkeep),
        .m_axis_fifo_76_tstrb(m_axis_fifo_76_tstrb),
        .m_axis_fifo_76_tdata(m_axis_fifo_76_tdata),
        .m_axis_fifo_76_tready(m_axis_fifo_76_tready),
        .ap_fifo_oarg_76_full_n(ap_fifo_oarg_76_full_n),
        .ap_fifo_oarg_76_din(ap_fifo_oarg_76_din),
        .ap_fifo_oarg_76_write(ap_fifo_oarg_76_write),
        .m_axis_fifo_77_aclk(m_axis_fifo_77_aclk),
        .m_axis_fifo_77_aresetn(m_axis_fifo_77_aresetn),
        .m_axis_fifo_77_tlast(m_axis_fifo_77_tlast),
        .m_axis_fifo_77_tvalid(m_axis_fifo_77_tvalid),
        .m_axis_fifo_77_tkeep(m_axis_fifo_77_tkeep),
        .m_axis_fifo_77_tstrb(m_axis_fifo_77_tstrb),
        .m_axis_fifo_77_tdata(m_axis_fifo_77_tdata),
        .m_axis_fifo_77_tready(m_axis_fifo_77_tready),
        .ap_fifo_oarg_77_full_n(ap_fifo_oarg_77_full_n),
        .ap_fifo_oarg_77_din(ap_fifo_oarg_77_din),
        .ap_fifo_oarg_77_write(ap_fifo_oarg_77_write),
        .m_axis_fifo_78_aclk(m_axis_fifo_78_aclk),
        .m_axis_fifo_78_aresetn(m_axis_fifo_78_aresetn),
        .m_axis_fifo_78_tlast(m_axis_fifo_78_tlast),
        .m_axis_fifo_78_tvalid(m_axis_fifo_78_tvalid),
        .m_axis_fifo_78_tkeep(m_axis_fifo_78_tkeep),
        .m_axis_fifo_78_tstrb(m_axis_fifo_78_tstrb),
        .m_axis_fifo_78_tdata(m_axis_fifo_78_tdata),
        .m_axis_fifo_78_tready(m_axis_fifo_78_tready),
        .ap_fifo_oarg_78_full_n(ap_fifo_oarg_78_full_n),
        .ap_fifo_oarg_78_din(ap_fifo_oarg_78_din),
        .ap_fifo_oarg_78_write(ap_fifo_oarg_78_write),
        .m_axis_fifo_79_aclk(m_axis_fifo_79_aclk),
        .m_axis_fifo_79_aresetn(m_axis_fifo_79_aresetn),
        .m_axis_fifo_79_tlast(m_axis_fifo_79_tlast),
        .m_axis_fifo_79_tvalid(m_axis_fifo_79_tvalid),
        .m_axis_fifo_79_tkeep(m_axis_fifo_79_tkeep),
        .m_axis_fifo_79_tstrb(m_axis_fifo_79_tstrb),
        .m_axis_fifo_79_tdata(m_axis_fifo_79_tdata),
        .m_axis_fifo_79_tready(m_axis_fifo_79_tready),
        .ap_fifo_oarg_79_full_n(ap_fifo_oarg_79_full_n),
        .ap_fifo_oarg_79_din(ap_fifo_oarg_79_din),
        .ap_fifo_oarg_79_write(ap_fifo_oarg_79_write),
        .m_axis_fifo_80_aclk(m_axis_fifo_80_aclk),
        .m_axis_fifo_80_aresetn(m_axis_fifo_80_aresetn),
        .m_axis_fifo_80_tlast(m_axis_fifo_80_tlast),
        .m_axis_fifo_80_tvalid(m_axis_fifo_80_tvalid),
        .m_axis_fifo_80_tkeep(m_axis_fifo_80_tkeep),
        .m_axis_fifo_80_tstrb(m_axis_fifo_80_tstrb),
        .m_axis_fifo_80_tdata(m_axis_fifo_80_tdata),
        .m_axis_fifo_80_tready(m_axis_fifo_80_tready),
        .ap_fifo_oarg_80_full_n(ap_fifo_oarg_80_full_n),
        .ap_fifo_oarg_80_din(ap_fifo_oarg_80_din),
        .ap_fifo_oarg_80_write(ap_fifo_oarg_80_write),
        .m_axis_fifo_81_aclk(m_axis_fifo_81_aclk),
        .m_axis_fifo_81_aresetn(m_axis_fifo_81_aresetn),
        .m_axis_fifo_81_tlast(m_axis_fifo_81_tlast),
        .m_axis_fifo_81_tvalid(m_axis_fifo_81_tvalid),
        .m_axis_fifo_81_tkeep(m_axis_fifo_81_tkeep),
        .m_axis_fifo_81_tstrb(m_axis_fifo_81_tstrb),
        .m_axis_fifo_81_tdata(m_axis_fifo_81_tdata),
        .m_axis_fifo_81_tready(m_axis_fifo_81_tready),
        .ap_fifo_oarg_81_full_n(ap_fifo_oarg_81_full_n),
        .ap_fifo_oarg_81_din(ap_fifo_oarg_81_din),
        .ap_fifo_oarg_81_write(ap_fifo_oarg_81_write),
        .m_axis_fifo_82_aclk(m_axis_fifo_82_aclk),
        .m_axis_fifo_82_aresetn(m_axis_fifo_82_aresetn),
        .m_axis_fifo_82_tlast(m_axis_fifo_82_tlast),
        .m_axis_fifo_82_tvalid(m_axis_fifo_82_tvalid),
        .m_axis_fifo_82_tkeep(m_axis_fifo_82_tkeep),
        .m_axis_fifo_82_tstrb(m_axis_fifo_82_tstrb),
        .m_axis_fifo_82_tdata(m_axis_fifo_82_tdata),
        .m_axis_fifo_82_tready(m_axis_fifo_82_tready),
        .ap_fifo_oarg_82_full_n(ap_fifo_oarg_82_full_n),
        .ap_fifo_oarg_82_din(ap_fifo_oarg_82_din),
        .ap_fifo_oarg_82_write(ap_fifo_oarg_82_write),
        .m_axis_fifo_83_aclk(m_axis_fifo_83_aclk),
        .m_axis_fifo_83_aresetn(m_axis_fifo_83_aresetn),
        .m_axis_fifo_83_tlast(m_axis_fifo_83_tlast),
        .m_axis_fifo_83_tvalid(m_axis_fifo_83_tvalid),
        .m_axis_fifo_83_tkeep(m_axis_fifo_83_tkeep),
        .m_axis_fifo_83_tstrb(m_axis_fifo_83_tstrb),
        .m_axis_fifo_83_tdata(m_axis_fifo_83_tdata),
        .m_axis_fifo_83_tready(m_axis_fifo_83_tready),
        .ap_fifo_oarg_83_full_n(ap_fifo_oarg_83_full_n),
        .ap_fifo_oarg_83_din(ap_fifo_oarg_83_din),
        .ap_fifo_oarg_83_write(ap_fifo_oarg_83_write),
        .m_axis_fifo_84_aclk(m_axis_fifo_84_aclk),
        .m_axis_fifo_84_aresetn(m_axis_fifo_84_aresetn),
        .m_axis_fifo_84_tlast(m_axis_fifo_84_tlast),
        .m_axis_fifo_84_tvalid(m_axis_fifo_84_tvalid),
        .m_axis_fifo_84_tkeep(m_axis_fifo_84_tkeep),
        .m_axis_fifo_84_tstrb(m_axis_fifo_84_tstrb),
        .m_axis_fifo_84_tdata(m_axis_fifo_84_tdata),
        .m_axis_fifo_84_tready(m_axis_fifo_84_tready),
        .ap_fifo_oarg_84_full_n(ap_fifo_oarg_84_full_n),
        .ap_fifo_oarg_84_din(ap_fifo_oarg_84_din),
        .ap_fifo_oarg_84_write(ap_fifo_oarg_84_write),
        .m_axis_fifo_85_aclk(m_axis_fifo_85_aclk),
        .m_axis_fifo_85_aresetn(m_axis_fifo_85_aresetn),
        .m_axis_fifo_85_tlast(m_axis_fifo_85_tlast),
        .m_axis_fifo_85_tvalid(m_axis_fifo_85_tvalid),
        .m_axis_fifo_85_tkeep(m_axis_fifo_85_tkeep),
        .m_axis_fifo_85_tstrb(m_axis_fifo_85_tstrb),
        .m_axis_fifo_85_tdata(m_axis_fifo_85_tdata),
        .m_axis_fifo_85_tready(m_axis_fifo_85_tready),
        .ap_fifo_oarg_85_full_n(ap_fifo_oarg_85_full_n),
        .ap_fifo_oarg_85_din(ap_fifo_oarg_85_din),
        .ap_fifo_oarg_85_write(ap_fifo_oarg_85_write),
        .m_axis_fifo_86_aclk(m_axis_fifo_86_aclk),
        .m_axis_fifo_86_aresetn(m_axis_fifo_86_aresetn),
        .m_axis_fifo_86_tlast(m_axis_fifo_86_tlast),
        .m_axis_fifo_86_tvalid(m_axis_fifo_86_tvalid),
        .m_axis_fifo_86_tkeep(m_axis_fifo_86_tkeep),
        .m_axis_fifo_86_tstrb(m_axis_fifo_86_tstrb),
        .m_axis_fifo_86_tdata(m_axis_fifo_86_tdata),
        .m_axis_fifo_86_tready(m_axis_fifo_86_tready),
        .ap_fifo_oarg_86_full_n(ap_fifo_oarg_86_full_n),
        .ap_fifo_oarg_86_din(ap_fifo_oarg_86_din),
        .ap_fifo_oarg_86_write(ap_fifo_oarg_86_write),
        .m_axis_fifo_87_aclk(m_axis_fifo_87_aclk),
        .m_axis_fifo_87_aresetn(m_axis_fifo_87_aresetn),
        .m_axis_fifo_87_tlast(m_axis_fifo_87_tlast),
        .m_axis_fifo_87_tvalid(m_axis_fifo_87_tvalid),
        .m_axis_fifo_87_tkeep(m_axis_fifo_87_tkeep),
        .m_axis_fifo_87_tstrb(m_axis_fifo_87_tstrb),
        .m_axis_fifo_87_tdata(m_axis_fifo_87_tdata),
        .m_axis_fifo_87_tready(m_axis_fifo_87_tready),
        .ap_fifo_oarg_87_full_n(ap_fifo_oarg_87_full_n),
        .ap_fifo_oarg_87_din(ap_fifo_oarg_87_din),
        .ap_fifo_oarg_87_write(ap_fifo_oarg_87_write),
        .m_axis_fifo_88_aclk(m_axis_fifo_88_aclk),
        .m_axis_fifo_88_aresetn(m_axis_fifo_88_aresetn),
        .m_axis_fifo_88_tlast(m_axis_fifo_88_tlast),
        .m_axis_fifo_88_tvalid(m_axis_fifo_88_tvalid),
        .m_axis_fifo_88_tkeep(m_axis_fifo_88_tkeep),
        .m_axis_fifo_88_tstrb(m_axis_fifo_88_tstrb),
        .m_axis_fifo_88_tdata(m_axis_fifo_88_tdata),
        .m_axis_fifo_88_tready(m_axis_fifo_88_tready),
        .ap_fifo_oarg_88_full_n(ap_fifo_oarg_88_full_n),
        .ap_fifo_oarg_88_din(ap_fifo_oarg_88_din),
        .ap_fifo_oarg_88_write(ap_fifo_oarg_88_write),
        .m_axis_fifo_89_aclk(m_axis_fifo_89_aclk),
        .m_axis_fifo_89_aresetn(m_axis_fifo_89_aresetn),
        .m_axis_fifo_89_tlast(m_axis_fifo_89_tlast),
        .m_axis_fifo_89_tvalid(m_axis_fifo_89_tvalid),
        .m_axis_fifo_89_tkeep(m_axis_fifo_89_tkeep),
        .m_axis_fifo_89_tstrb(m_axis_fifo_89_tstrb),
        .m_axis_fifo_89_tdata(m_axis_fifo_89_tdata),
        .m_axis_fifo_89_tready(m_axis_fifo_89_tready),
        .ap_fifo_oarg_89_full_n(ap_fifo_oarg_89_full_n),
        .ap_fifo_oarg_89_din(ap_fifo_oarg_89_din),
        .ap_fifo_oarg_89_write(ap_fifo_oarg_89_write),
        .m_axis_fifo_90_aclk(m_axis_fifo_90_aclk),
        .m_axis_fifo_90_aresetn(m_axis_fifo_90_aresetn),
        .m_axis_fifo_90_tlast(m_axis_fifo_90_tlast),
        .m_axis_fifo_90_tvalid(m_axis_fifo_90_tvalid),
        .m_axis_fifo_90_tkeep(m_axis_fifo_90_tkeep),
        .m_axis_fifo_90_tstrb(m_axis_fifo_90_tstrb),
        .m_axis_fifo_90_tdata(m_axis_fifo_90_tdata),
        .m_axis_fifo_90_tready(m_axis_fifo_90_tready),
        .ap_fifo_oarg_90_full_n(ap_fifo_oarg_90_full_n),
        .ap_fifo_oarg_90_din(ap_fifo_oarg_90_din),
        .ap_fifo_oarg_90_write(ap_fifo_oarg_90_write),
        .m_axis_fifo_91_aclk(m_axis_fifo_91_aclk),
        .m_axis_fifo_91_aresetn(m_axis_fifo_91_aresetn),
        .m_axis_fifo_91_tlast(m_axis_fifo_91_tlast),
        .m_axis_fifo_91_tvalid(m_axis_fifo_91_tvalid),
        .m_axis_fifo_91_tkeep(m_axis_fifo_91_tkeep),
        .m_axis_fifo_91_tstrb(m_axis_fifo_91_tstrb),
        .m_axis_fifo_91_tdata(m_axis_fifo_91_tdata),
        .m_axis_fifo_91_tready(m_axis_fifo_91_tready),
        .ap_fifo_oarg_91_full_n(ap_fifo_oarg_91_full_n),
        .ap_fifo_oarg_91_din(ap_fifo_oarg_91_din),
        .ap_fifo_oarg_91_write(ap_fifo_oarg_91_write),
        .m_axis_fifo_92_aclk(m_axis_fifo_92_aclk),
        .m_axis_fifo_92_aresetn(m_axis_fifo_92_aresetn),
        .m_axis_fifo_92_tlast(m_axis_fifo_92_tlast),
        .m_axis_fifo_92_tvalid(m_axis_fifo_92_tvalid),
        .m_axis_fifo_92_tkeep(m_axis_fifo_92_tkeep),
        .m_axis_fifo_92_tstrb(m_axis_fifo_92_tstrb),
        .m_axis_fifo_92_tdata(m_axis_fifo_92_tdata),
        .m_axis_fifo_92_tready(m_axis_fifo_92_tready),
        .ap_fifo_oarg_92_full_n(ap_fifo_oarg_92_full_n),
        .ap_fifo_oarg_92_din(ap_fifo_oarg_92_din),
        .ap_fifo_oarg_92_write(ap_fifo_oarg_92_write),
        .m_axis_fifo_93_aclk(m_axis_fifo_93_aclk),
        .m_axis_fifo_93_aresetn(m_axis_fifo_93_aresetn),
        .m_axis_fifo_93_tlast(m_axis_fifo_93_tlast),
        .m_axis_fifo_93_tvalid(m_axis_fifo_93_tvalid),
        .m_axis_fifo_93_tkeep(m_axis_fifo_93_tkeep),
        .m_axis_fifo_93_tstrb(m_axis_fifo_93_tstrb),
        .m_axis_fifo_93_tdata(m_axis_fifo_93_tdata),
        .m_axis_fifo_93_tready(m_axis_fifo_93_tready),
        .ap_fifo_oarg_93_full_n(ap_fifo_oarg_93_full_n),
        .ap_fifo_oarg_93_din(ap_fifo_oarg_93_din),
        .ap_fifo_oarg_93_write(ap_fifo_oarg_93_write),
        .m_axis_fifo_94_aclk(m_axis_fifo_94_aclk),
        .m_axis_fifo_94_aresetn(m_axis_fifo_94_aresetn),
        .m_axis_fifo_94_tlast(m_axis_fifo_94_tlast),
        .m_axis_fifo_94_tvalid(m_axis_fifo_94_tvalid),
        .m_axis_fifo_94_tkeep(m_axis_fifo_94_tkeep),
        .m_axis_fifo_94_tstrb(m_axis_fifo_94_tstrb),
        .m_axis_fifo_94_tdata(m_axis_fifo_94_tdata),
        .m_axis_fifo_94_tready(m_axis_fifo_94_tready),
        .ap_fifo_oarg_94_full_n(ap_fifo_oarg_94_full_n),
        .ap_fifo_oarg_94_din(ap_fifo_oarg_94_din),
        .ap_fifo_oarg_94_write(ap_fifo_oarg_94_write),
        .m_axis_fifo_95_aclk(m_axis_fifo_95_aclk),
        .m_axis_fifo_95_aresetn(m_axis_fifo_95_aresetn),
        .m_axis_fifo_95_tlast(m_axis_fifo_95_tlast),
        .m_axis_fifo_95_tvalid(m_axis_fifo_95_tvalid),
        .m_axis_fifo_95_tkeep(m_axis_fifo_95_tkeep),
        .m_axis_fifo_95_tstrb(m_axis_fifo_95_tstrb),
        .m_axis_fifo_95_tdata(m_axis_fifo_95_tdata),
        .m_axis_fifo_95_tready(m_axis_fifo_95_tready),
        .ap_fifo_oarg_95_full_n(ap_fifo_oarg_95_full_n),
        .ap_fifo_oarg_95_din(ap_fifo_oarg_95_din),
        .ap_fifo_oarg_95_write(ap_fifo_oarg_95_write),
        .m_axis_fifo_96_aclk(m_axis_fifo_96_aclk),
        .m_axis_fifo_96_aresetn(m_axis_fifo_96_aresetn),
        .m_axis_fifo_96_tlast(m_axis_fifo_96_tlast),
        .m_axis_fifo_96_tvalid(m_axis_fifo_96_tvalid),
        .m_axis_fifo_96_tkeep(m_axis_fifo_96_tkeep),
        .m_axis_fifo_96_tstrb(m_axis_fifo_96_tstrb),
        .m_axis_fifo_96_tdata(m_axis_fifo_96_tdata),
        .m_axis_fifo_96_tready(m_axis_fifo_96_tready),
        .ap_fifo_oarg_96_full_n(ap_fifo_oarg_96_full_n),
        .ap_fifo_oarg_96_din(ap_fifo_oarg_96_din),
        .ap_fifo_oarg_96_write(ap_fifo_oarg_96_write),
        .m_axis_fifo_97_aclk(m_axis_fifo_97_aclk),
        .m_axis_fifo_97_aresetn(m_axis_fifo_97_aresetn),
        .m_axis_fifo_97_tlast(m_axis_fifo_97_tlast),
        .m_axis_fifo_97_tvalid(m_axis_fifo_97_tvalid),
        .m_axis_fifo_97_tkeep(m_axis_fifo_97_tkeep),
        .m_axis_fifo_97_tstrb(m_axis_fifo_97_tstrb),
        .m_axis_fifo_97_tdata(m_axis_fifo_97_tdata),
        .m_axis_fifo_97_tready(m_axis_fifo_97_tready),
        .ap_fifo_oarg_97_full_n(ap_fifo_oarg_97_full_n),
        .ap_fifo_oarg_97_din(ap_fifo_oarg_97_din),
        .ap_fifo_oarg_97_write(ap_fifo_oarg_97_write),
        .m_axis_fifo_98_aclk(m_axis_fifo_98_aclk),
        .m_axis_fifo_98_aresetn(m_axis_fifo_98_aresetn),
        .m_axis_fifo_98_tlast(m_axis_fifo_98_tlast),
        .m_axis_fifo_98_tvalid(m_axis_fifo_98_tvalid),
        .m_axis_fifo_98_tkeep(m_axis_fifo_98_tkeep),
        .m_axis_fifo_98_tstrb(m_axis_fifo_98_tstrb),
        .m_axis_fifo_98_tdata(m_axis_fifo_98_tdata),
        .m_axis_fifo_98_tready(m_axis_fifo_98_tready),
        .ap_fifo_oarg_98_full_n(ap_fifo_oarg_98_full_n),
        .ap_fifo_oarg_98_din(ap_fifo_oarg_98_din),
        .ap_fifo_oarg_98_write(ap_fifo_oarg_98_write),
        .m_axis_fifo_99_aclk(m_axis_fifo_99_aclk),
        .m_axis_fifo_99_aresetn(m_axis_fifo_99_aresetn),
        .m_axis_fifo_99_tlast(m_axis_fifo_99_tlast),
        .m_axis_fifo_99_tvalid(m_axis_fifo_99_tvalid),
        .m_axis_fifo_99_tkeep(m_axis_fifo_99_tkeep),
        .m_axis_fifo_99_tstrb(m_axis_fifo_99_tstrb),
        .m_axis_fifo_99_tdata(m_axis_fifo_99_tdata),
        .m_axis_fifo_99_tready(m_axis_fifo_99_tready),
        .ap_fifo_oarg_99_full_n(ap_fifo_oarg_99_full_n),
        .ap_fifo_oarg_99_din(ap_fifo_oarg_99_din),
        .ap_fifo_oarg_99_write(ap_fifo_oarg_99_write),
        .m_axis_fifo_100_aclk(m_axis_fifo_100_aclk),
        .m_axis_fifo_100_aresetn(m_axis_fifo_100_aresetn),
        .m_axis_fifo_100_tlast(m_axis_fifo_100_tlast),
        .m_axis_fifo_100_tvalid(m_axis_fifo_100_tvalid),
        .m_axis_fifo_100_tkeep(m_axis_fifo_100_tkeep),
        .m_axis_fifo_100_tstrb(m_axis_fifo_100_tstrb),
        .m_axis_fifo_100_tdata(m_axis_fifo_100_tdata),
        .m_axis_fifo_100_tready(m_axis_fifo_100_tready),
        .ap_fifo_oarg_100_full_n(ap_fifo_oarg_100_full_n),
        .ap_fifo_oarg_100_din(ap_fifo_oarg_100_din),
        .ap_fifo_oarg_100_write(ap_fifo_oarg_100_write),
        .m_axis_fifo_101_aclk(m_axis_fifo_101_aclk),
        .m_axis_fifo_101_aresetn(m_axis_fifo_101_aresetn),
        .m_axis_fifo_101_tlast(m_axis_fifo_101_tlast),
        .m_axis_fifo_101_tvalid(m_axis_fifo_101_tvalid),
        .m_axis_fifo_101_tkeep(m_axis_fifo_101_tkeep),
        .m_axis_fifo_101_tstrb(m_axis_fifo_101_tstrb),
        .m_axis_fifo_101_tdata(m_axis_fifo_101_tdata),
        .m_axis_fifo_101_tready(m_axis_fifo_101_tready),
        .ap_fifo_oarg_101_full_n(ap_fifo_oarg_101_full_n),
        .ap_fifo_oarg_101_din(ap_fifo_oarg_101_din),
        .ap_fifo_oarg_101_write(ap_fifo_oarg_101_write),
        .m_axis_fifo_102_aclk(m_axis_fifo_102_aclk),
        .m_axis_fifo_102_aresetn(m_axis_fifo_102_aresetn),
        .m_axis_fifo_102_tlast(m_axis_fifo_102_tlast),
        .m_axis_fifo_102_tvalid(m_axis_fifo_102_tvalid),
        .m_axis_fifo_102_tkeep(m_axis_fifo_102_tkeep),
        .m_axis_fifo_102_tstrb(m_axis_fifo_102_tstrb),
        .m_axis_fifo_102_tdata(m_axis_fifo_102_tdata),
        .m_axis_fifo_102_tready(m_axis_fifo_102_tready),
        .ap_fifo_oarg_102_full_n(ap_fifo_oarg_102_full_n),
        .ap_fifo_oarg_102_din(ap_fifo_oarg_102_din),
        .ap_fifo_oarg_102_write(ap_fifo_oarg_102_write),
        .m_axis_fifo_103_aclk(m_axis_fifo_103_aclk),
        .m_axis_fifo_103_aresetn(m_axis_fifo_103_aresetn),
        .m_axis_fifo_103_tlast(m_axis_fifo_103_tlast),
        .m_axis_fifo_103_tvalid(m_axis_fifo_103_tvalid),
        .m_axis_fifo_103_tkeep(m_axis_fifo_103_tkeep),
        .m_axis_fifo_103_tstrb(m_axis_fifo_103_tstrb),
        .m_axis_fifo_103_tdata(m_axis_fifo_103_tdata),
        .m_axis_fifo_103_tready(m_axis_fifo_103_tready),
        .ap_fifo_oarg_103_full_n(ap_fifo_oarg_103_full_n),
        .ap_fifo_oarg_103_din(ap_fifo_oarg_103_din),
        .ap_fifo_oarg_103_write(ap_fifo_oarg_103_write),
        .m_axis_fifo_104_aclk(m_axis_fifo_104_aclk),
        .m_axis_fifo_104_aresetn(m_axis_fifo_104_aresetn),
        .m_axis_fifo_104_tlast(m_axis_fifo_104_tlast),
        .m_axis_fifo_104_tvalid(m_axis_fifo_104_tvalid),
        .m_axis_fifo_104_tkeep(m_axis_fifo_104_tkeep),
        .m_axis_fifo_104_tstrb(m_axis_fifo_104_tstrb),
        .m_axis_fifo_104_tdata(m_axis_fifo_104_tdata),
        .m_axis_fifo_104_tready(m_axis_fifo_104_tready),
        .ap_fifo_oarg_104_full_n(ap_fifo_oarg_104_full_n),
        .ap_fifo_oarg_104_din(ap_fifo_oarg_104_din),
        .ap_fifo_oarg_104_write(ap_fifo_oarg_104_write),
        .m_axis_fifo_105_aclk(m_axis_fifo_105_aclk),
        .m_axis_fifo_105_aresetn(m_axis_fifo_105_aresetn),
        .m_axis_fifo_105_tlast(m_axis_fifo_105_tlast),
        .m_axis_fifo_105_tvalid(m_axis_fifo_105_tvalid),
        .m_axis_fifo_105_tkeep(m_axis_fifo_105_tkeep),
        .m_axis_fifo_105_tstrb(m_axis_fifo_105_tstrb),
        .m_axis_fifo_105_tdata(m_axis_fifo_105_tdata),
        .m_axis_fifo_105_tready(m_axis_fifo_105_tready),
        .ap_fifo_oarg_105_full_n(ap_fifo_oarg_105_full_n),
        .ap_fifo_oarg_105_din(ap_fifo_oarg_105_din),
        .ap_fifo_oarg_105_write(ap_fifo_oarg_105_write),
        .m_axis_fifo_106_aclk(m_axis_fifo_106_aclk),
        .m_axis_fifo_106_aresetn(m_axis_fifo_106_aresetn),
        .m_axis_fifo_106_tlast(m_axis_fifo_106_tlast),
        .m_axis_fifo_106_tvalid(m_axis_fifo_106_tvalid),
        .m_axis_fifo_106_tkeep(m_axis_fifo_106_tkeep),
        .m_axis_fifo_106_tstrb(m_axis_fifo_106_tstrb),
        .m_axis_fifo_106_tdata(m_axis_fifo_106_tdata),
        .m_axis_fifo_106_tready(m_axis_fifo_106_tready),
        .ap_fifo_oarg_106_full_n(ap_fifo_oarg_106_full_n),
        .ap_fifo_oarg_106_din(ap_fifo_oarg_106_din),
        .ap_fifo_oarg_106_write(ap_fifo_oarg_106_write),
        .m_axis_fifo_107_aclk(m_axis_fifo_107_aclk),
        .m_axis_fifo_107_aresetn(m_axis_fifo_107_aresetn),
        .m_axis_fifo_107_tlast(m_axis_fifo_107_tlast),
        .m_axis_fifo_107_tvalid(m_axis_fifo_107_tvalid),
        .m_axis_fifo_107_tkeep(m_axis_fifo_107_tkeep),
        .m_axis_fifo_107_tstrb(m_axis_fifo_107_tstrb),
        .m_axis_fifo_107_tdata(m_axis_fifo_107_tdata),
        .m_axis_fifo_107_tready(m_axis_fifo_107_tready),
        .ap_fifo_oarg_107_full_n(ap_fifo_oarg_107_full_n),
        .ap_fifo_oarg_107_din(ap_fifo_oarg_107_din),
        .ap_fifo_oarg_107_write(ap_fifo_oarg_107_write),
        .m_axis_fifo_108_aclk(m_axis_fifo_108_aclk),
        .m_axis_fifo_108_aresetn(m_axis_fifo_108_aresetn),
        .m_axis_fifo_108_tlast(m_axis_fifo_108_tlast),
        .m_axis_fifo_108_tvalid(m_axis_fifo_108_tvalid),
        .m_axis_fifo_108_tkeep(m_axis_fifo_108_tkeep),
        .m_axis_fifo_108_tstrb(m_axis_fifo_108_tstrb),
        .m_axis_fifo_108_tdata(m_axis_fifo_108_tdata),
        .m_axis_fifo_108_tready(m_axis_fifo_108_tready),
        .ap_fifo_oarg_108_full_n(ap_fifo_oarg_108_full_n),
        .ap_fifo_oarg_108_din(ap_fifo_oarg_108_din),
        .ap_fifo_oarg_108_write(ap_fifo_oarg_108_write),
        .m_axis_fifo_109_aclk(m_axis_fifo_109_aclk),
        .m_axis_fifo_109_aresetn(m_axis_fifo_109_aresetn),
        .m_axis_fifo_109_tlast(m_axis_fifo_109_tlast),
        .m_axis_fifo_109_tvalid(m_axis_fifo_109_tvalid),
        .m_axis_fifo_109_tkeep(m_axis_fifo_109_tkeep),
        .m_axis_fifo_109_tstrb(m_axis_fifo_109_tstrb),
        .m_axis_fifo_109_tdata(m_axis_fifo_109_tdata),
        .m_axis_fifo_109_tready(m_axis_fifo_109_tready),
        .ap_fifo_oarg_109_full_n(ap_fifo_oarg_109_full_n),
        .ap_fifo_oarg_109_din(ap_fifo_oarg_109_din),
        .ap_fifo_oarg_109_write(ap_fifo_oarg_109_write),
        .m_axis_fifo_110_aclk(m_axis_fifo_110_aclk),
        .m_axis_fifo_110_aresetn(m_axis_fifo_110_aresetn),
        .m_axis_fifo_110_tlast(m_axis_fifo_110_tlast),
        .m_axis_fifo_110_tvalid(m_axis_fifo_110_tvalid),
        .m_axis_fifo_110_tkeep(m_axis_fifo_110_tkeep),
        .m_axis_fifo_110_tstrb(m_axis_fifo_110_tstrb),
        .m_axis_fifo_110_tdata(m_axis_fifo_110_tdata),
        .m_axis_fifo_110_tready(m_axis_fifo_110_tready),
        .ap_fifo_oarg_110_full_n(ap_fifo_oarg_110_full_n),
        .ap_fifo_oarg_110_din(ap_fifo_oarg_110_din),
        .ap_fifo_oarg_110_write(ap_fifo_oarg_110_write),
        .m_axis_fifo_111_aclk(m_axis_fifo_111_aclk),
        .m_axis_fifo_111_aresetn(m_axis_fifo_111_aresetn),
        .m_axis_fifo_111_tlast(m_axis_fifo_111_tlast),
        .m_axis_fifo_111_tvalid(m_axis_fifo_111_tvalid),
        .m_axis_fifo_111_tkeep(m_axis_fifo_111_tkeep),
        .m_axis_fifo_111_tstrb(m_axis_fifo_111_tstrb),
        .m_axis_fifo_111_tdata(m_axis_fifo_111_tdata),
        .m_axis_fifo_111_tready(m_axis_fifo_111_tready),
        .ap_fifo_oarg_111_full_n(ap_fifo_oarg_111_full_n),
        .ap_fifo_oarg_111_din(ap_fifo_oarg_111_din),
        .ap_fifo_oarg_111_write(ap_fifo_oarg_111_write),
        .m_axis_fifo_112_aclk(m_axis_fifo_112_aclk),
        .m_axis_fifo_112_aresetn(m_axis_fifo_112_aresetn),
        .m_axis_fifo_112_tlast(m_axis_fifo_112_tlast),
        .m_axis_fifo_112_tvalid(m_axis_fifo_112_tvalid),
        .m_axis_fifo_112_tkeep(m_axis_fifo_112_tkeep),
        .m_axis_fifo_112_tstrb(m_axis_fifo_112_tstrb),
        .m_axis_fifo_112_tdata(m_axis_fifo_112_tdata),
        .m_axis_fifo_112_tready(m_axis_fifo_112_tready),
        .ap_fifo_oarg_112_full_n(ap_fifo_oarg_112_full_n),
        .ap_fifo_oarg_112_din(ap_fifo_oarg_112_din),
        .ap_fifo_oarg_112_write(ap_fifo_oarg_112_write),
        .m_axis_fifo_113_aclk(m_axis_fifo_113_aclk),
        .m_axis_fifo_113_aresetn(m_axis_fifo_113_aresetn),
        .m_axis_fifo_113_tlast(m_axis_fifo_113_tlast),
        .m_axis_fifo_113_tvalid(m_axis_fifo_113_tvalid),
        .m_axis_fifo_113_tkeep(m_axis_fifo_113_tkeep),
        .m_axis_fifo_113_tstrb(m_axis_fifo_113_tstrb),
        .m_axis_fifo_113_tdata(m_axis_fifo_113_tdata),
        .m_axis_fifo_113_tready(m_axis_fifo_113_tready),
        .ap_fifo_oarg_113_full_n(ap_fifo_oarg_113_full_n),
        .ap_fifo_oarg_113_din(ap_fifo_oarg_113_din),
        .ap_fifo_oarg_113_write(ap_fifo_oarg_113_write),
        .m_axis_fifo_114_aclk(m_axis_fifo_114_aclk),
        .m_axis_fifo_114_aresetn(m_axis_fifo_114_aresetn),
        .m_axis_fifo_114_tlast(m_axis_fifo_114_tlast),
        .m_axis_fifo_114_tvalid(m_axis_fifo_114_tvalid),
        .m_axis_fifo_114_tkeep(m_axis_fifo_114_tkeep),
        .m_axis_fifo_114_tstrb(m_axis_fifo_114_tstrb),
        .m_axis_fifo_114_tdata(m_axis_fifo_114_tdata),
        .m_axis_fifo_114_tready(m_axis_fifo_114_tready),
        .ap_fifo_oarg_114_full_n(ap_fifo_oarg_114_full_n),
        .ap_fifo_oarg_114_din(ap_fifo_oarg_114_din),
        .ap_fifo_oarg_114_write(ap_fifo_oarg_114_write),
        .m_axis_fifo_115_aclk(m_axis_fifo_115_aclk),
        .m_axis_fifo_115_aresetn(m_axis_fifo_115_aresetn),
        .m_axis_fifo_115_tlast(m_axis_fifo_115_tlast),
        .m_axis_fifo_115_tvalid(m_axis_fifo_115_tvalid),
        .m_axis_fifo_115_tkeep(m_axis_fifo_115_tkeep),
        .m_axis_fifo_115_tstrb(m_axis_fifo_115_tstrb),
        .m_axis_fifo_115_tdata(m_axis_fifo_115_tdata),
        .m_axis_fifo_115_tready(m_axis_fifo_115_tready),
        .ap_fifo_oarg_115_full_n(ap_fifo_oarg_115_full_n),
        .ap_fifo_oarg_115_din(ap_fifo_oarg_115_din),
        .ap_fifo_oarg_115_write(ap_fifo_oarg_115_write),
        .m_axis_fifo_116_aclk(m_axis_fifo_116_aclk),
        .m_axis_fifo_116_aresetn(m_axis_fifo_116_aresetn),
        .m_axis_fifo_116_tlast(m_axis_fifo_116_tlast),
        .m_axis_fifo_116_tvalid(m_axis_fifo_116_tvalid),
        .m_axis_fifo_116_tkeep(m_axis_fifo_116_tkeep),
        .m_axis_fifo_116_tstrb(m_axis_fifo_116_tstrb),
        .m_axis_fifo_116_tdata(m_axis_fifo_116_tdata),
        .m_axis_fifo_116_tready(m_axis_fifo_116_tready),
        .ap_fifo_oarg_116_full_n(ap_fifo_oarg_116_full_n),
        .ap_fifo_oarg_116_din(ap_fifo_oarg_116_din),
        .ap_fifo_oarg_116_write(ap_fifo_oarg_116_write),
        .m_axis_fifo_117_aclk(m_axis_fifo_117_aclk),
        .m_axis_fifo_117_aresetn(m_axis_fifo_117_aresetn),
        .m_axis_fifo_117_tlast(m_axis_fifo_117_tlast),
        .m_axis_fifo_117_tvalid(m_axis_fifo_117_tvalid),
        .m_axis_fifo_117_tkeep(m_axis_fifo_117_tkeep),
        .m_axis_fifo_117_tstrb(m_axis_fifo_117_tstrb),
        .m_axis_fifo_117_tdata(m_axis_fifo_117_tdata),
        .m_axis_fifo_117_tready(m_axis_fifo_117_tready),
        .ap_fifo_oarg_117_full_n(ap_fifo_oarg_117_full_n),
        .ap_fifo_oarg_117_din(ap_fifo_oarg_117_din),
        .ap_fifo_oarg_117_write(ap_fifo_oarg_117_write),
        .m_axis_fifo_118_aclk(m_axis_fifo_118_aclk),
        .m_axis_fifo_118_aresetn(m_axis_fifo_118_aresetn),
        .m_axis_fifo_118_tlast(m_axis_fifo_118_tlast),
        .m_axis_fifo_118_tvalid(m_axis_fifo_118_tvalid),
        .m_axis_fifo_118_tkeep(m_axis_fifo_118_tkeep),
        .m_axis_fifo_118_tstrb(m_axis_fifo_118_tstrb),
        .m_axis_fifo_118_tdata(m_axis_fifo_118_tdata),
        .m_axis_fifo_118_tready(m_axis_fifo_118_tready),
        .ap_fifo_oarg_118_full_n(ap_fifo_oarg_118_full_n),
        .ap_fifo_oarg_118_din(ap_fifo_oarg_118_din),
        .ap_fifo_oarg_118_write(ap_fifo_oarg_118_write),
        .m_axis_fifo_119_aclk(m_axis_fifo_119_aclk),
        .m_axis_fifo_119_aresetn(m_axis_fifo_119_aresetn),
        .m_axis_fifo_119_tlast(m_axis_fifo_119_tlast),
        .m_axis_fifo_119_tvalid(m_axis_fifo_119_tvalid),
        .m_axis_fifo_119_tkeep(m_axis_fifo_119_tkeep),
        .m_axis_fifo_119_tstrb(m_axis_fifo_119_tstrb),
        .m_axis_fifo_119_tdata(m_axis_fifo_119_tdata),
        .m_axis_fifo_119_tready(m_axis_fifo_119_tready),
        .ap_fifo_oarg_119_full_n(ap_fifo_oarg_119_full_n),
        .ap_fifo_oarg_119_din(ap_fifo_oarg_119_din),
        .ap_fifo_oarg_119_write(ap_fifo_oarg_119_write),
        .m_axis_fifo_120_aclk(m_axis_fifo_120_aclk),
        .m_axis_fifo_120_aresetn(m_axis_fifo_120_aresetn),
        .m_axis_fifo_120_tlast(m_axis_fifo_120_tlast),
        .m_axis_fifo_120_tvalid(m_axis_fifo_120_tvalid),
        .m_axis_fifo_120_tkeep(m_axis_fifo_120_tkeep),
        .m_axis_fifo_120_tstrb(m_axis_fifo_120_tstrb),
        .m_axis_fifo_120_tdata(m_axis_fifo_120_tdata),
        .m_axis_fifo_120_tready(m_axis_fifo_120_tready),
        .ap_fifo_oarg_120_full_n(ap_fifo_oarg_120_full_n),
        .ap_fifo_oarg_120_din(ap_fifo_oarg_120_din),
        .ap_fifo_oarg_120_write(ap_fifo_oarg_120_write),
        .m_axis_fifo_121_aclk(m_axis_fifo_121_aclk),
        .m_axis_fifo_121_aresetn(m_axis_fifo_121_aresetn),
        .m_axis_fifo_121_tlast(m_axis_fifo_121_tlast),
        .m_axis_fifo_121_tvalid(m_axis_fifo_121_tvalid),
        .m_axis_fifo_121_tkeep(m_axis_fifo_121_tkeep),
        .m_axis_fifo_121_tstrb(m_axis_fifo_121_tstrb),
        .m_axis_fifo_121_tdata(m_axis_fifo_121_tdata),
        .m_axis_fifo_121_tready(m_axis_fifo_121_tready),
        .ap_fifo_oarg_121_full_n(ap_fifo_oarg_121_full_n),
        .ap_fifo_oarg_121_din(ap_fifo_oarg_121_din),
        .ap_fifo_oarg_121_write(ap_fifo_oarg_121_write),
        .m_axis_fifo_122_aclk(m_axis_fifo_122_aclk),
        .m_axis_fifo_122_aresetn(m_axis_fifo_122_aresetn),
        .m_axis_fifo_122_tlast(m_axis_fifo_122_tlast),
        .m_axis_fifo_122_tvalid(m_axis_fifo_122_tvalid),
        .m_axis_fifo_122_tkeep(m_axis_fifo_122_tkeep),
        .m_axis_fifo_122_tstrb(m_axis_fifo_122_tstrb),
        .m_axis_fifo_122_tdata(m_axis_fifo_122_tdata),
        .m_axis_fifo_122_tready(m_axis_fifo_122_tready),
        .ap_fifo_oarg_122_full_n(ap_fifo_oarg_122_full_n),
        .ap_fifo_oarg_122_din(ap_fifo_oarg_122_din),
        .ap_fifo_oarg_122_write(ap_fifo_oarg_122_write),
        .m_axis_fifo_123_aclk(m_axis_fifo_123_aclk),
        .m_axis_fifo_123_aresetn(m_axis_fifo_123_aresetn),
        .m_axis_fifo_123_tlast(m_axis_fifo_123_tlast),
        .m_axis_fifo_123_tvalid(m_axis_fifo_123_tvalid),
        .m_axis_fifo_123_tkeep(m_axis_fifo_123_tkeep),
        .m_axis_fifo_123_tstrb(m_axis_fifo_123_tstrb),
        .m_axis_fifo_123_tdata(m_axis_fifo_123_tdata),
        .m_axis_fifo_123_tready(m_axis_fifo_123_tready),
        .ap_fifo_oarg_123_full_n(ap_fifo_oarg_123_full_n),
        .ap_fifo_oarg_123_din(ap_fifo_oarg_123_din),
        .ap_fifo_oarg_123_write(ap_fifo_oarg_123_write),
        .m_axis_fifo_124_aclk(m_axis_fifo_124_aclk),
        .m_axis_fifo_124_aresetn(m_axis_fifo_124_aresetn),
        .m_axis_fifo_124_tlast(m_axis_fifo_124_tlast),
        .m_axis_fifo_124_tvalid(m_axis_fifo_124_tvalid),
        .m_axis_fifo_124_tkeep(m_axis_fifo_124_tkeep),
        .m_axis_fifo_124_tstrb(m_axis_fifo_124_tstrb),
        .m_axis_fifo_124_tdata(m_axis_fifo_124_tdata),
        .m_axis_fifo_124_tready(m_axis_fifo_124_tready),
        .ap_fifo_oarg_124_full_n(ap_fifo_oarg_124_full_n),
        .ap_fifo_oarg_124_din(ap_fifo_oarg_124_din),
        .ap_fifo_oarg_124_write(ap_fifo_oarg_124_write),
        .m_axis_fifo_125_aclk(m_axis_fifo_125_aclk),
        .m_axis_fifo_125_aresetn(m_axis_fifo_125_aresetn),
        .m_axis_fifo_125_tlast(m_axis_fifo_125_tlast),
        .m_axis_fifo_125_tvalid(m_axis_fifo_125_tvalid),
        .m_axis_fifo_125_tkeep(m_axis_fifo_125_tkeep),
        .m_axis_fifo_125_tstrb(m_axis_fifo_125_tstrb),
        .m_axis_fifo_125_tdata(m_axis_fifo_125_tdata),
        .m_axis_fifo_125_tready(m_axis_fifo_125_tready),
        .ap_fifo_oarg_125_full_n(ap_fifo_oarg_125_full_n),
        .ap_fifo_oarg_125_din(ap_fifo_oarg_125_din),
        .ap_fifo_oarg_125_write(ap_fifo_oarg_125_write),
        .m_axis_fifo_126_aclk(m_axis_fifo_126_aclk),
        .m_axis_fifo_126_aresetn(m_axis_fifo_126_aresetn),
        .m_axis_fifo_126_tlast(m_axis_fifo_126_tlast),
        .m_axis_fifo_126_tvalid(m_axis_fifo_126_tvalid),
        .m_axis_fifo_126_tkeep(m_axis_fifo_126_tkeep),
        .m_axis_fifo_126_tstrb(m_axis_fifo_126_tstrb),
        .m_axis_fifo_126_tdata(m_axis_fifo_126_tdata),
        .m_axis_fifo_126_tready(m_axis_fifo_126_tready),
        .ap_fifo_oarg_126_full_n(ap_fifo_oarg_126_full_n),
        .ap_fifo_oarg_126_din(ap_fifo_oarg_126_din),
        .ap_fifo_oarg_126_write(ap_fifo_oarg_126_write),
        .m_axis_fifo_127_aclk(m_axis_fifo_127_aclk),
        .m_axis_fifo_127_aresetn(m_axis_fifo_127_aresetn),
        .m_axis_fifo_127_tlast(m_axis_fifo_127_tlast),
        .m_axis_fifo_127_tvalid(m_axis_fifo_127_tvalid),
        .m_axis_fifo_127_tkeep(m_axis_fifo_127_tkeep),
        .m_axis_fifo_127_tstrb(m_axis_fifo_127_tstrb),
        .m_axis_fifo_127_tdata(m_axis_fifo_127_tdata),
        .m_axis_fifo_127_tready(m_axis_fifo_127_tready),
        .ap_fifo_oarg_127_full_n(ap_fifo_oarg_127_full_n),
        .ap_fifo_oarg_127_din(ap_fifo_oarg_127_din),
        .ap_fifo_oarg_127_write(ap_fifo_oarg_127_write)
    );
    
    
    in_axis_args #(
        .C_NUM_INPUT_AXISs(C_NUM_INPUT_AXISs),
        .S_AXIS_IARG_0_WIDTH(S_AXIS_IARG_0_WIDTH),
        .S_AXIS_IARG_1_WIDTH(S_AXIS_IARG_1_WIDTH),
        .S_AXIS_IARG_2_WIDTH(S_AXIS_IARG_2_WIDTH),
        .S_AXIS_IARG_3_WIDTH(S_AXIS_IARG_3_WIDTH),
        .S_AXIS_IARG_4_WIDTH(S_AXIS_IARG_4_WIDTH),
        .S_AXIS_IARG_5_WIDTH(S_AXIS_IARG_5_WIDTH),
        .S_AXIS_IARG_6_WIDTH(S_AXIS_IARG_6_WIDTH),
        .S_AXIS_IARG_7_WIDTH(S_AXIS_IARG_7_WIDTH),
        .S_AXIS_IARG_8_WIDTH(S_AXIS_IARG_8_WIDTH),
        .S_AXIS_IARG_9_WIDTH(S_AXIS_IARG_9_WIDTH),
        .S_AXIS_IARG_10_WIDTH(S_AXIS_IARG_10_WIDTH),
        .S_AXIS_IARG_11_WIDTH(S_AXIS_IARG_11_WIDTH),
        .S_AXIS_IARG_12_WIDTH(S_AXIS_IARG_12_WIDTH),
        .S_AXIS_IARG_13_WIDTH(S_AXIS_IARG_13_WIDTH),
        .S_AXIS_IARG_14_WIDTH(S_AXIS_IARG_14_WIDTH),
        .S_AXIS_IARG_15_WIDTH(S_AXIS_IARG_15_WIDTH),
        .S_AXIS_IARG_16_WIDTH(S_AXIS_IARG_16_WIDTH),
        .S_AXIS_IARG_17_WIDTH(S_AXIS_IARG_17_WIDTH),
        .S_AXIS_IARG_18_WIDTH(S_AXIS_IARG_18_WIDTH),
        .S_AXIS_IARG_19_WIDTH(S_AXIS_IARG_19_WIDTH),
        .S_AXIS_IARG_20_WIDTH(S_AXIS_IARG_20_WIDTH),
        .S_AXIS_IARG_21_WIDTH(S_AXIS_IARG_21_WIDTH),
        .S_AXIS_IARG_22_WIDTH(S_AXIS_IARG_22_WIDTH),
        .S_AXIS_IARG_23_WIDTH(S_AXIS_IARG_23_WIDTH),
        .S_AXIS_IARG_24_WIDTH(S_AXIS_IARG_24_WIDTH),
        .S_AXIS_IARG_25_WIDTH(S_AXIS_IARG_25_WIDTH),
        .S_AXIS_IARG_26_WIDTH(S_AXIS_IARG_26_WIDTH),
        .S_AXIS_IARG_27_WIDTH(S_AXIS_IARG_27_WIDTH),
        .S_AXIS_IARG_28_WIDTH(S_AXIS_IARG_28_WIDTH),
        .S_AXIS_IARG_29_WIDTH(S_AXIS_IARG_29_WIDTH),
        .S_AXIS_IARG_30_WIDTH(S_AXIS_IARG_30_WIDTH),
        .S_AXIS_IARG_31_WIDTH(S_AXIS_IARG_31_WIDTH),
        .S_AXIS_IARG_32_WIDTH(S_AXIS_IARG_32_WIDTH),
        .S_AXIS_IARG_33_WIDTH(S_AXIS_IARG_33_WIDTH),
        .S_AXIS_IARG_34_WIDTH(S_AXIS_IARG_34_WIDTH),
        .S_AXIS_IARG_35_WIDTH(S_AXIS_IARG_35_WIDTH),
        .S_AXIS_IARG_36_WIDTH(S_AXIS_IARG_36_WIDTH),
        .S_AXIS_IARG_37_WIDTH(S_AXIS_IARG_37_WIDTH),
        .S_AXIS_IARG_38_WIDTH(S_AXIS_IARG_38_WIDTH),
        .S_AXIS_IARG_39_WIDTH(S_AXIS_IARG_39_WIDTH),
        .S_AXIS_IARG_40_WIDTH(S_AXIS_IARG_40_WIDTH),
        .S_AXIS_IARG_41_WIDTH(S_AXIS_IARG_41_WIDTH),
        .S_AXIS_IARG_42_WIDTH(S_AXIS_IARG_42_WIDTH),
        .S_AXIS_IARG_43_WIDTH(S_AXIS_IARG_43_WIDTH),
        .S_AXIS_IARG_44_WIDTH(S_AXIS_IARG_44_WIDTH),
        .S_AXIS_IARG_45_WIDTH(S_AXIS_IARG_45_WIDTH),
        .S_AXIS_IARG_46_WIDTH(S_AXIS_IARG_46_WIDTH),
        .S_AXIS_IARG_47_WIDTH(S_AXIS_IARG_47_WIDTH),
        .S_AXIS_IARG_48_WIDTH(S_AXIS_IARG_48_WIDTH),
        .S_AXIS_IARG_49_WIDTH(S_AXIS_IARG_49_WIDTH),
        .S_AXIS_IARG_50_WIDTH(S_AXIS_IARG_50_WIDTH),
        .S_AXIS_IARG_51_WIDTH(S_AXIS_IARG_51_WIDTH),
        .S_AXIS_IARG_52_WIDTH(S_AXIS_IARG_52_WIDTH),
        .S_AXIS_IARG_53_WIDTH(S_AXIS_IARG_53_WIDTH),
        .S_AXIS_IARG_54_WIDTH(S_AXIS_IARG_54_WIDTH),
        .S_AXIS_IARG_55_WIDTH(S_AXIS_IARG_55_WIDTH),
        .S_AXIS_IARG_56_WIDTH(S_AXIS_IARG_56_WIDTH),
        .S_AXIS_IARG_57_WIDTH(S_AXIS_IARG_57_WIDTH),
        .S_AXIS_IARG_58_WIDTH(S_AXIS_IARG_58_WIDTH),
        .S_AXIS_IARG_59_WIDTH(S_AXIS_IARG_59_WIDTH),
        .S_AXIS_IARG_60_WIDTH(S_AXIS_IARG_60_WIDTH),
        .S_AXIS_IARG_61_WIDTH(S_AXIS_IARG_61_WIDTH),
        .S_AXIS_IARG_62_WIDTH(S_AXIS_IARG_62_WIDTH),
        .S_AXIS_IARG_63_WIDTH(S_AXIS_IARG_63_WIDTH),
        .S_AXIS_IARG_64_WIDTH(S_AXIS_IARG_64_WIDTH),
        .S_AXIS_IARG_65_WIDTH(S_AXIS_IARG_65_WIDTH),
        .S_AXIS_IARG_66_WIDTH(S_AXIS_IARG_66_WIDTH),
        .S_AXIS_IARG_67_WIDTH(S_AXIS_IARG_67_WIDTH),
        .S_AXIS_IARG_68_WIDTH(S_AXIS_IARG_68_WIDTH),
        .S_AXIS_IARG_69_WIDTH(S_AXIS_IARG_69_WIDTH),
        .S_AXIS_IARG_70_WIDTH(S_AXIS_IARG_70_WIDTH),
        .S_AXIS_IARG_71_WIDTH(S_AXIS_IARG_71_WIDTH),
        .S_AXIS_IARG_72_WIDTH(S_AXIS_IARG_72_WIDTH),
        .S_AXIS_IARG_73_WIDTH(S_AXIS_IARG_73_WIDTH),
        .S_AXIS_IARG_74_WIDTH(S_AXIS_IARG_74_WIDTH),
        .S_AXIS_IARG_75_WIDTH(S_AXIS_IARG_75_WIDTH),
        .S_AXIS_IARG_76_WIDTH(S_AXIS_IARG_76_WIDTH),
        .S_AXIS_IARG_77_WIDTH(S_AXIS_IARG_77_WIDTH),
        .S_AXIS_IARG_78_WIDTH(S_AXIS_IARG_78_WIDTH),
        .S_AXIS_IARG_79_WIDTH(S_AXIS_IARG_79_WIDTH),
        .S_AXIS_IARG_80_WIDTH(S_AXIS_IARG_80_WIDTH),
        .S_AXIS_IARG_81_WIDTH(S_AXIS_IARG_81_WIDTH),
        .S_AXIS_IARG_82_WIDTH(S_AXIS_IARG_82_WIDTH),
        .S_AXIS_IARG_83_WIDTH(S_AXIS_IARG_83_WIDTH),
        .S_AXIS_IARG_84_WIDTH(S_AXIS_IARG_84_WIDTH),
        .S_AXIS_IARG_85_WIDTH(S_AXIS_IARG_85_WIDTH),
        .S_AXIS_IARG_86_WIDTH(S_AXIS_IARG_86_WIDTH),
        .S_AXIS_IARG_87_WIDTH(S_AXIS_IARG_87_WIDTH),
        .S_AXIS_IARG_88_WIDTH(S_AXIS_IARG_88_WIDTH),
        .S_AXIS_IARG_89_WIDTH(S_AXIS_IARG_89_WIDTH),
        .S_AXIS_IARG_90_WIDTH(S_AXIS_IARG_90_WIDTH),
        .S_AXIS_IARG_91_WIDTH(S_AXIS_IARG_91_WIDTH),
        .S_AXIS_IARG_92_WIDTH(S_AXIS_IARG_92_WIDTH),
        .S_AXIS_IARG_93_WIDTH(S_AXIS_IARG_93_WIDTH),
        .S_AXIS_IARG_94_WIDTH(S_AXIS_IARG_94_WIDTH),
        .S_AXIS_IARG_95_WIDTH(S_AXIS_IARG_95_WIDTH),
        .S_AXIS_IARG_96_WIDTH(S_AXIS_IARG_96_WIDTH),
        .S_AXIS_IARG_97_WIDTH(S_AXIS_IARG_97_WIDTH),
        .S_AXIS_IARG_98_WIDTH(S_AXIS_IARG_98_WIDTH),
        .S_AXIS_IARG_99_WIDTH(S_AXIS_IARG_99_WIDTH),
        .S_AXIS_IARG_100_WIDTH(S_AXIS_IARG_100_WIDTH),
        .S_AXIS_IARG_101_WIDTH(S_AXIS_IARG_101_WIDTH),
        .S_AXIS_IARG_102_WIDTH(S_AXIS_IARG_102_WIDTH),
        .S_AXIS_IARG_103_WIDTH(S_AXIS_IARG_103_WIDTH),
        .S_AXIS_IARG_104_WIDTH(S_AXIS_IARG_104_WIDTH),
        .S_AXIS_IARG_105_WIDTH(S_AXIS_IARG_105_WIDTH),
        .S_AXIS_IARG_106_WIDTH(S_AXIS_IARG_106_WIDTH),
        .S_AXIS_IARG_107_WIDTH(S_AXIS_IARG_107_WIDTH),
        .S_AXIS_IARG_108_WIDTH(S_AXIS_IARG_108_WIDTH),
        .S_AXIS_IARG_109_WIDTH(S_AXIS_IARG_109_WIDTH),
        .S_AXIS_IARG_110_WIDTH(S_AXIS_IARG_110_WIDTH),
        .S_AXIS_IARG_111_WIDTH(S_AXIS_IARG_111_WIDTH),
        .S_AXIS_IARG_112_WIDTH(S_AXIS_IARG_112_WIDTH),
        .S_AXIS_IARG_113_WIDTH(S_AXIS_IARG_113_WIDTH),
        .S_AXIS_IARG_114_WIDTH(S_AXIS_IARG_114_WIDTH),
        .S_AXIS_IARG_115_WIDTH(S_AXIS_IARG_115_WIDTH),
        .S_AXIS_IARG_116_WIDTH(S_AXIS_IARG_116_WIDTH),
        .S_AXIS_IARG_117_WIDTH(S_AXIS_IARG_117_WIDTH),
        .S_AXIS_IARG_118_WIDTH(S_AXIS_IARG_118_WIDTH),
        .S_AXIS_IARG_119_WIDTH(S_AXIS_IARG_119_WIDTH),
        .S_AXIS_IARG_120_WIDTH(S_AXIS_IARG_120_WIDTH),
        .S_AXIS_IARG_121_WIDTH(S_AXIS_IARG_121_WIDTH),
        .S_AXIS_IARG_122_WIDTH(S_AXIS_IARG_122_WIDTH),
        .S_AXIS_IARG_123_WIDTH(S_AXIS_IARG_123_WIDTH),
        .S_AXIS_IARG_124_WIDTH(S_AXIS_IARG_124_WIDTH),
        .S_AXIS_IARG_125_WIDTH(S_AXIS_IARG_125_WIDTH),
        .S_AXIS_IARG_126_WIDTH(S_AXIS_IARG_126_WIDTH),
        .S_AXIS_IARG_127_WIDTH(S_AXIS_IARG_127_WIDTH),
        .S_AXIS_IARG_0_DEPTH(S_AXIS_IARG_0_DEPTH),
        .S_AXIS_IARG_1_DEPTH(S_AXIS_IARG_1_DEPTH),
        .S_AXIS_IARG_2_DEPTH(S_AXIS_IARG_2_DEPTH),
        .S_AXIS_IARG_3_DEPTH(S_AXIS_IARG_3_DEPTH),
        .S_AXIS_IARG_4_DEPTH(S_AXIS_IARG_4_DEPTH),
        .S_AXIS_IARG_5_DEPTH(S_AXIS_IARG_5_DEPTH),
        .S_AXIS_IARG_6_DEPTH(S_AXIS_IARG_6_DEPTH),
        .S_AXIS_IARG_7_DEPTH(S_AXIS_IARG_7_DEPTH),
        .S_AXIS_IARG_8_DEPTH(S_AXIS_IARG_8_DEPTH),
        .S_AXIS_IARG_9_DEPTH(S_AXIS_IARG_9_DEPTH),
        .S_AXIS_IARG_10_DEPTH(S_AXIS_IARG_10_DEPTH),
        .S_AXIS_IARG_11_DEPTH(S_AXIS_IARG_11_DEPTH),
        .S_AXIS_IARG_12_DEPTH(S_AXIS_IARG_12_DEPTH),
        .S_AXIS_IARG_13_DEPTH(S_AXIS_IARG_13_DEPTH),
        .S_AXIS_IARG_14_DEPTH(S_AXIS_IARG_14_DEPTH),
        .S_AXIS_IARG_15_DEPTH(S_AXIS_IARG_15_DEPTH),
        .S_AXIS_IARG_16_DEPTH(S_AXIS_IARG_16_DEPTH),
        .S_AXIS_IARG_17_DEPTH(S_AXIS_IARG_17_DEPTH),
        .S_AXIS_IARG_18_DEPTH(S_AXIS_IARG_18_DEPTH),
        .S_AXIS_IARG_19_DEPTH(S_AXIS_IARG_19_DEPTH),
        .S_AXIS_IARG_20_DEPTH(S_AXIS_IARG_20_DEPTH),
        .S_AXIS_IARG_21_DEPTH(S_AXIS_IARG_21_DEPTH),
        .S_AXIS_IARG_22_DEPTH(S_AXIS_IARG_22_DEPTH),
        .S_AXIS_IARG_23_DEPTH(S_AXIS_IARG_23_DEPTH),
        .S_AXIS_IARG_24_DEPTH(S_AXIS_IARG_24_DEPTH),
        .S_AXIS_IARG_25_DEPTH(S_AXIS_IARG_25_DEPTH),
        .S_AXIS_IARG_26_DEPTH(S_AXIS_IARG_26_DEPTH),
        .S_AXIS_IARG_27_DEPTH(S_AXIS_IARG_27_DEPTH),
        .S_AXIS_IARG_28_DEPTH(S_AXIS_IARG_28_DEPTH),
        .S_AXIS_IARG_29_DEPTH(S_AXIS_IARG_29_DEPTH),
        .S_AXIS_IARG_30_DEPTH(S_AXIS_IARG_30_DEPTH),
        .S_AXIS_IARG_31_DEPTH(S_AXIS_IARG_31_DEPTH),
        .S_AXIS_IARG_32_DEPTH(S_AXIS_IARG_32_DEPTH),
        .S_AXIS_IARG_33_DEPTH(S_AXIS_IARG_33_DEPTH),
        .S_AXIS_IARG_34_DEPTH(S_AXIS_IARG_34_DEPTH),
        .S_AXIS_IARG_35_DEPTH(S_AXIS_IARG_35_DEPTH),
        .S_AXIS_IARG_36_DEPTH(S_AXIS_IARG_36_DEPTH),
        .S_AXIS_IARG_37_DEPTH(S_AXIS_IARG_37_DEPTH),
        .S_AXIS_IARG_38_DEPTH(S_AXIS_IARG_38_DEPTH),
        .S_AXIS_IARG_39_DEPTH(S_AXIS_IARG_39_DEPTH),
        .S_AXIS_IARG_40_DEPTH(S_AXIS_IARG_40_DEPTH),
        .S_AXIS_IARG_41_DEPTH(S_AXIS_IARG_41_DEPTH),
        .S_AXIS_IARG_42_DEPTH(S_AXIS_IARG_42_DEPTH),
        .S_AXIS_IARG_43_DEPTH(S_AXIS_IARG_43_DEPTH),
        .S_AXIS_IARG_44_DEPTH(S_AXIS_IARG_44_DEPTH),
        .S_AXIS_IARG_45_DEPTH(S_AXIS_IARG_45_DEPTH),
        .S_AXIS_IARG_46_DEPTH(S_AXIS_IARG_46_DEPTH),
        .S_AXIS_IARG_47_DEPTH(S_AXIS_IARG_47_DEPTH),
        .S_AXIS_IARG_48_DEPTH(S_AXIS_IARG_48_DEPTH),
        .S_AXIS_IARG_49_DEPTH(S_AXIS_IARG_49_DEPTH),
        .S_AXIS_IARG_50_DEPTH(S_AXIS_IARG_50_DEPTH),
        .S_AXIS_IARG_51_DEPTH(S_AXIS_IARG_51_DEPTH),
        .S_AXIS_IARG_52_DEPTH(S_AXIS_IARG_52_DEPTH),
        .S_AXIS_IARG_53_DEPTH(S_AXIS_IARG_53_DEPTH),
        .S_AXIS_IARG_54_DEPTH(S_AXIS_IARG_54_DEPTH),
        .S_AXIS_IARG_55_DEPTH(S_AXIS_IARG_55_DEPTH),
        .S_AXIS_IARG_56_DEPTH(S_AXIS_IARG_56_DEPTH),
        .S_AXIS_IARG_57_DEPTH(S_AXIS_IARG_57_DEPTH),
        .S_AXIS_IARG_58_DEPTH(S_AXIS_IARG_58_DEPTH),
        .S_AXIS_IARG_59_DEPTH(S_AXIS_IARG_59_DEPTH),
        .S_AXIS_IARG_60_DEPTH(S_AXIS_IARG_60_DEPTH),
        .S_AXIS_IARG_61_DEPTH(S_AXIS_IARG_61_DEPTH),
        .S_AXIS_IARG_62_DEPTH(S_AXIS_IARG_62_DEPTH),
        .S_AXIS_IARG_63_DEPTH(S_AXIS_IARG_63_DEPTH),
        .S_AXIS_IARG_64_DEPTH(S_AXIS_IARG_64_DEPTH),
        .S_AXIS_IARG_65_DEPTH(S_AXIS_IARG_65_DEPTH),
        .S_AXIS_IARG_66_DEPTH(S_AXIS_IARG_66_DEPTH),
        .S_AXIS_IARG_67_DEPTH(S_AXIS_IARG_67_DEPTH),
        .S_AXIS_IARG_68_DEPTH(S_AXIS_IARG_68_DEPTH),
        .S_AXIS_IARG_69_DEPTH(S_AXIS_IARG_69_DEPTH),
        .S_AXIS_IARG_70_DEPTH(S_AXIS_IARG_70_DEPTH),
        .S_AXIS_IARG_71_DEPTH(S_AXIS_IARG_71_DEPTH),
        .S_AXIS_IARG_72_DEPTH(S_AXIS_IARG_72_DEPTH),
        .S_AXIS_IARG_73_DEPTH(S_AXIS_IARG_73_DEPTH),
        .S_AXIS_IARG_74_DEPTH(S_AXIS_IARG_74_DEPTH),
        .S_AXIS_IARG_75_DEPTH(S_AXIS_IARG_75_DEPTH),
        .S_AXIS_IARG_76_DEPTH(S_AXIS_IARG_76_DEPTH),
        .S_AXIS_IARG_77_DEPTH(S_AXIS_IARG_77_DEPTH),
        .S_AXIS_IARG_78_DEPTH(S_AXIS_IARG_78_DEPTH),
        .S_AXIS_IARG_79_DEPTH(S_AXIS_IARG_79_DEPTH),
        .S_AXIS_IARG_80_DEPTH(S_AXIS_IARG_80_DEPTH),
        .S_AXIS_IARG_81_DEPTH(S_AXIS_IARG_81_DEPTH),
        .S_AXIS_IARG_82_DEPTH(S_AXIS_IARG_82_DEPTH),
        .S_AXIS_IARG_83_DEPTH(S_AXIS_IARG_83_DEPTH),
        .S_AXIS_IARG_84_DEPTH(S_AXIS_IARG_84_DEPTH),
        .S_AXIS_IARG_85_DEPTH(S_AXIS_IARG_85_DEPTH),
        .S_AXIS_IARG_86_DEPTH(S_AXIS_IARG_86_DEPTH),
        .S_AXIS_IARG_87_DEPTH(S_AXIS_IARG_87_DEPTH),
        .S_AXIS_IARG_88_DEPTH(S_AXIS_IARG_88_DEPTH),
        .S_AXIS_IARG_89_DEPTH(S_AXIS_IARG_89_DEPTH),
        .S_AXIS_IARG_90_DEPTH(S_AXIS_IARG_90_DEPTH),
        .S_AXIS_IARG_91_DEPTH(S_AXIS_IARG_91_DEPTH),
        .S_AXIS_IARG_92_DEPTH(S_AXIS_IARG_92_DEPTH),
        .S_AXIS_IARG_93_DEPTH(S_AXIS_IARG_93_DEPTH),
        .S_AXIS_IARG_94_DEPTH(S_AXIS_IARG_94_DEPTH),
        .S_AXIS_IARG_95_DEPTH(S_AXIS_IARG_95_DEPTH),
        .S_AXIS_IARG_96_DEPTH(S_AXIS_IARG_96_DEPTH),
        .S_AXIS_IARG_97_DEPTH(S_AXIS_IARG_97_DEPTH),
        .S_AXIS_IARG_98_DEPTH(S_AXIS_IARG_98_DEPTH),
        .S_AXIS_IARG_99_DEPTH(S_AXIS_IARG_99_DEPTH),
        .S_AXIS_IARG_100_DEPTH(S_AXIS_IARG_100_DEPTH),
        .S_AXIS_IARG_101_DEPTH(S_AXIS_IARG_101_DEPTH),
        .S_AXIS_IARG_102_DEPTH(S_AXIS_IARG_102_DEPTH),
        .S_AXIS_IARG_103_DEPTH(S_AXIS_IARG_103_DEPTH),
        .S_AXIS_IARG_104_DEPTH(S_AXIS_IARG_104_DEPTH),
        .S_AXIS_IARG_105_DEPTH(S_AXIS_IARG_105_DEPTH),
        .S_AXIS_IARG_106_DEPTH(S_AXIS_IARG_106_DEPTH),
        .S_AXIS_IARG_107_DEPTH(S_AXIS_IARG_107_DEPTH),
        .S_AXIS_IARG_108_DEPTH(S_AXIS_IARG_108_DEPTH),
        .S_AXIS_IARG_109_DEPTH(S_AXIS_IARG_109_DEPTH),
        .S_AXIS_IARG_110_DEPTH(S_AXIS_IARG_110_DEPTH),
        .S_AXIS_IARG_111_DEPTH(S_AXIS_IARG_111_DEPTH),
        .S_AXIS_IARG_112_DEPTH(S_AXIS_IARG_112_DEPTH),
        .S_AXIS_IARG_113_DEPTH(S_AXIS_IARG_113_DEPTH),
        .S_AXIS_IARG_114_DEPTH(S_AXIS_IARG_114_DEPTH),
        .S_AXIS_IARG_115_DEPTH(S_AXIS_IARG_115_DEPTH),
        .S_AXIS_IARG_116_DEPTH(S_AXIS_IARG_116_DEPTH),
        .S_AXIS_IARG_117_DEPTH(S_AXIS_IARG_117_DEPTH),
        .S_AXIS_IARG_118_DEPTH(S_AXIS_IARG_118_DEPTH),
        .S_AXIS_IARG_119_DEPTH(S_AXIS_IARG_119_DEPTH),
        .S_AXIS_IARG_120_DEPTH(S_AXIS_IARG_120_DEPTH),
        .S_AXIS_IARG_121_DEPTH(S_AXIS_IARG_121_DEPTH),
        .S_AXIS_IARG_122_DEPTH(S_AXIS_IARG_122_DEPTH),
        .S_AXIS_IARG_123_DEPTH(S_AXIS_IARG_123_DEPTH),
        .S_AXIS_IARG_124_DEPTH(S_AXIS_IARG_124_DEPTH),
        .S_AXIS_IARG_125_DEPTH(S_AXIS_IARG_125_DEPTH),
        .S_AXIS_IARG_126_DEPTH(S_AXIS_IARG_126_DEPTH),
        .S_AXIS_IARG_127_DEPTH(S_AXIS_IARG_127_DEPTH),
        .S_AXIS_IARG_0_IS_ASYNC(S_AXIS_IARG_0_IS_ASYNC),
        .S_AXIS_IARG_1_IS_ASYNC(S_AXIS_IARG_1_IS_ASYNC),
        .S_AXIS_IARG_2_IS_ASYNC(S_AXIS_IARG_2_IS_ASYNC),
        .S_AXIS_IARG_3_IS_ASYNC(S_AXIS_IARG_3_IS_ASYNC),
        .S_AXIS_IARG_4_IS_ASYNC(S_AXIS_IARG_4_IS_ASYNC),
        .S_AXIS_IARG_5_IS_ASYNC(S_AXIS_IARG_5_IS_ASYNC),
        .S_AXIS_IARG_6_IS_ASYNC(S_AXIS_IARG_6_IS_ASYNC),
        .S_AXIS_IARG_7_IS_ASYNC(S_AXIS_IARG_7_IS_ASYNC),
        .S_AXIS_IARG_8_IS_ASYNC(S_AXIS_IARG_8_IS_ASYNC),
        .S_AXIS_IARG_9_IS_ASYNC(S_AXIS_IARG_9_IS_ASYNC),
        .S_AXIS_IARG_10_IS_ASYNC(S_AXIS_IARG_10_IS_ASYNC),
        .S_AXIS_IARG_11_IS_ASYNC(S_AXIS_IARG_11_IS_ASYNC),
        .S_AXIS_IARG_12_IS_ASYNC(S_AXIS_IARG_12_IS_ASYNC),
        .S_AXIS_IARG_13_IS_ASYNC(S_AXIS_IARG_13_IS_ASYNC),
        .S_AXIS_IARG_14_IS_ASYNC(S_AXIS_IARG_14_IS_ASYNC),
        .S_AXIS_IARG_15_IS_ASYNC(S_AXIS_IARG_15_IS_ASYNC),
        .S_AXIS_IARG_16_IS_ASYNC(S_AXIS_IARG_16_IS_ASYNC),
        .S_AXIS_IARG_17_IS_ASYNC(S_AXIS_IARG_17_IS_ASYNC),
        .S_AXIS_IARG_18_IS_ASYNC(S_AXIS_IARG_18_IS_ASYNC),
        .S_AXIS_IARG_19_IS_ASYNC(S_AXIS_IARG_19_IS_ASYNC),
        .S_AXIS_IARG_20_IS_ASYNC(S_AXIS_IARG_20_IS_ASYNC),
        .S_AXIS_IARG_21_IS_ASYNC(S_AXIS_IARG_21_IS_ASYNC),
        .S_AXIS_IARG_22_IS_ASYNC(S_AXIS_IARG_22_IS_ASYNC),
        .S_AXIS_IARG_23_IS_ASYNC(S_AXIS_IARG_23_IS_ASYNC),
        .S_AXIS_IARG_24_IS_ASYNC(S_AXIS_IARG_24_IS_ASYNC),
        .S_AXIS_IARG_25_IS_ASYNC(S_AXIS_IARG_25_IS_ASYNC),
        .S_AXIS_IARG_26_IS_ASYNC(S_AXIS_IARG_26_IS_ASYNC),
        .S_AXIS_IARG_27_IS_ASYNC(S_AXIS_IARG_27_IS_ASYNC),
        .S_AXIS_IARG_28_IS_ASYNC(S_AXIS_IARG_28_IS_ASYNC),
        .S_AXIS_IARG_29_IS_ASYNC(S_AXIS_IARG_29_IS_ASYNC),
        .S_AXIS_IARG_30_IS_ASYNC(S_AXIS_IARG_30_IS_ASYNC),
        .S_AXIS_IARG_31_IS_ASYNC(S_AXIS_IARG_31_IS_ASYNC),
        .S_AXIS_IARG_32_IS_ASYNC(S_AXIS_IARG_32_IS_ASYNC),
        .S_AXIS_IARG_33_IS_ASYNC(S_AXIS_IARG_33_IS_ASYNC),
        .S_AXIS_IARG_34_IS_ASYNC(S_AXIS_IARG_34_IS_ASYNC),
        .S_AXIS_IARG_35_IS_ASYNC(S_AXIS_IARG_35_IS_ASYNC),
        .S_AXIS_IARG_36_IS_ASYNC(S_AXIS_IARG_36_IS_ASYNC),
        .S_AXIS_IARG_37_IS_ASYNC(S_AXIS_IARG_37_IS_ASYNC),
        .S_AXIS_IARG_38_IS_ASYNC(S_AXIS_IARG_38_IS_ASYNC),
        .S_AXIS_IARG_39_IS_ASYNC(S_AXIS_IARG_39_IS_ASYNC),
        .S_AXIS_IARG_40_IS_ASYNC(S_AXIS_IARG_40_IS_ASYNC),
        .S_AXIS_IARG_41_IS_ASYNC(S_AXIS_IARG_41_IS_ASYNC),
        .S_AXIS_IARG_42_IS_ASYNC(S_AXIS_IARG_42_IS_ASYNC),
        .S_AXIS_IARG_43_IS_ASYNC(S_AXIS_IARG_43_IS_ASYNC),
        .S_AXIS_IARG_44_IS_ASYNC(S_AXIS_IARG_44_IS_ASYNC),
        .S_AXIS_IARG_45_IS_ASYNC(S_AXIS_IARG_45_IS_ASYNC),
        .S_AXIS_IARG_46_IS_ASYNC(S_AXIS_IARG_46_IS_ASYNC),
        .S_AXIS_IARG_47_IS_ASYNC(S_AXIS_IARG_47_IS_ASYNC),
        .S_AXIS_IARG_48_IS_ASYNC(S_AXIS_IARG_48_IS_ASYNC),
        .S_AXIS_IARG_49_IS_ASYNC(S_AXIS_IARG_49_IS_ASYNC),
        .S_AXIS_IARG_50_IS_ASYNC(S_AXIS_IARG_50_IS_ASYNC),
        .S_AXIS_IARG_51_IS_ASYNC(S_AXIS_IARG_51_IS_ASYNC),
        .S_AXIS_IARG_52_IS_ASYNC(S_AXIS_IARG_52_IS_ASYNC),
        .S_AXIS_IARG_53_IS_ASYNC(S_AXIS_IARG_53_IS_ASYNC),
        .S_AXIS_IARG_54_IS_ASYNC(S_AXIS_IARG_54_IS_ASYNC),
        .S_AXIS_IARG_55_IS_ASYNC(S_AXIS_IARG_55_IS_ASYNC),
        .S_AXIS_IARG_56_IS_ASYNC(S_AXIS_IARG_56_IS_ASYNC),
        .S_AXIS_IARG_57_IS_ASYNC(S_AXIS_IARG_57_IS_ASYNC),
        .S_AXIS_IARG_58_IS_ASYNC(S_AXIS_IARG_58_IS_ASYNC),
        .S_AXIS_IARG_59_IS_ASYNC(S_AXIS_IARG_59_IS_ASYNC),
        .S_AXIS_IARG_60_IS_ASYNC(S_AXIS_IARG_60_IS_ASYNC),
        .S_AXIS_IARG_61_IS_ASYNC(S_AXIS_IARG_61_IS_ASYNC),
        .S_AXIS_IARG_62_IS_ASYNC(S_AXIS_IARG_62_IS_ASYNC),
        .S_AXIS_IARG_63_IS_ASYNC(S_AXIS_IARG_63_IS_ASYNC),
        .S_AXIS_IARG_64_IS_ASYNC(S_AXIS_IARG_64_IS_ASYNC),
        .S_AXIS_IARG_65_IS_ASYNC(S_AXIS_IARG_65_IS_ASYNC),
        .S_AXIS_IARG_66_IS_ASYNC(S_AXIS_IARG_66_IS_ASYNC),
        .S_AXIS_IARG_67_IS_ASYNC(S_AXIS_IARG_67_IS_ASYNC),
        .S_AXIS_IARG_68_IS_ASYNC(S_AXIS_IARG_68_IS_ASYNC),
        .S_AXIS_IARG_69_IS_ASYNC(S_AXIS_IARG_69_IS_ASYNC),
        .S_AXIS_IARG_70_IS_ASYNC(S_AXIS_IARG_70_IS_ASYNC),
        .S_AXIS_IARG_71_IS_ASYNC(S_AXIS_IARG_71_IS_ASYNC),
        .S_AXIS_IARG_72_IS_ASYNC(S_AXIS_IARG_72_IS_ASYNC),
        .S_AXIS_IARG_73_IS_ASYNC(S_AXIS_IARG_73_IS_ASYNC),
        .S_AXIS_IARG_74_IS_ASYNC(S_AXIS_IARG_74_IS_ASYNC),
        .S_AXIS_IARG_75_IS_ASYNC(S_AXIS_IARG_75_IS_ASYNC),
        .S_AXIS_IARG_76_IS_ASYNC(S_AXIS_IARG_76_IS_ASYNC),
        .S_AXIS_IARG_77_IS_ASYNC(S_AXIS_IARG_77_IS_ASYNC),
        .S_AXIS_IARG_78_IS_ASYNC(S_AXIS_IARG_78_IS_ASYNC),
        .S_AXIS_IARG_79_IS_ASYNC(S_AXIS_IARG_79_IS_ASYNC),
        .S_AXIS_IARG_80_IS_ASYNC(S_AXIS_IARG_80_IS_ASYNC),
        .S_AXIS_IARG_81_IS_ASYNC(S_AXIS_IARG_81_IS_ASYNC),
        .S_AXIS_IARG_82_IS_ASYNC(S_AXIS_IARG_82_IS_ASYNC),
        .S_AXIS_IARG_83_IS_ASYNC(S_AXIS_IARG_83_IS_ASYNC),
        .S_AXIS_IARG_84_IS_ASYNC(S_AXIS_IARG_84_IS_ASYNC),
        .S_AXIS_IARG_85_IS_ASYNC(S_AXIS_IARG_85_IS_ASYNC),
        .S_AXIS_IARG_86_IS_ASYNC(S_AXIS_IARG_86_IS_ASYNC),
        .S_AXIS_IARG_87_IS_ASYNC(S_AXIS_IARG_87_IS_ASYNC),
        .S_AXIS_IARG_88_IS_ASYNC(S_AXIS_IARG_88_IS_ASYNC),
        .S_AXIS_IARG_89_IS_ASYNC(S_AXIS_IARG_89_IS_ASYNC),
        .S_AXIS_IARG_90_IS_ASYNC(S_AXIS_IARG_90_IS_ASYNC),
        .S_AXIS_IARG_91_IS_ASYNC(S_AXIS_IARG_91_IS_ASYNC),
        .S_AXIS_IARG_92_IS_ASYNC(S_AXIS_IARG_92_IS_ASYNC),
        .S_AXIS_IARG_93_IS_ASYNC(S_AXIS_IARG_93_IS_ASYNC),
        .S_AXIS_IARG_94_IS_ASYNC(S_AXIS_IARG_94_IS_ASYNC),
        .S_AXIS_IARG_95_IS_ASYNC(S_AXIS_IARG_95_IS_ASYNC),
        .S_AXIS_IARG_96_IS_ASYNC(S_AXIS_IARG_96_IS_ASYNC),
        .S_AXIS_IARG_97_IS_ASYNC(S_AXIS_IARG_97_IS_ASYNC),
        .S_AXIS_IARG_98_IS_ASYNC(S_AXIS_IARG_98_IS_ASYNC),
        .S_AXIS_IARG_99_IS_ASYNC(S_AXIS_IARG_99_IS_ASYNC),
        .S_AXIS_IARG_100_IS_ASYNC(S_AXIS_IARG_100_IS_ASYNC),
        .S_AXIS_IARG_101_IS_ASYNC(S_AXIS_IARG_101_IS_ASYNC),
        .S_AXIS_IARG_102_IS_ASYNC(S_AXIS_IARG_102_IS_ASYNC),
        .S_AXIS_IARG_103_IS_ASYNC(S_AXIS_IARG_103_IS_ASYNC),
        .S_AXIS_IARG_104_IS_ASYNC(S_AXIS_IARG_104_IS_ASYNC),
        .S_AXIS_IARG_105_IS_ASYNC(S_AXIS_IARG_105_IS_ASYNC),
        .S_AXIS_IARG_106_IS_ASYNC(S_AXIS_IARG_106_IS_ASYNC),
        .S_AXIS_IARG_107_IS_ASYNC(S_AXIS_IARG_107_IS_ASYNC),
        .S_AXIS_IARG_108_IS_ASYNC(S_AXIS_IARG_108_IS_ASYNC),
        .S_AXIS_IARG_109_IS_ASYNC(S_AXIS_IARG_109_IS_ASYNC),
        .S_AXIS_IARG_110_IS_ASYNC(S_AXIS_IARG_110_IS_ASYNC),
        .S_AXIS_IARG_111_IS_ASYNC(S_AXIS_IARG_111_IS_ASYNC),
        .S_AXIS_IARG_112_IS_ASYNC(S_AXIS_IARG_112_IS_ASYNC),
        .S_AXIS_IARG_113_IS_ASYNC(S_AXIS_IARG_113_IS_ASYNC),
        .S_AXIS_IARG_114_IS_ASYNC(S_AXIS_IARG_114_IS_ASYNC),
        .S_AXIS_IARG_115_IS_ASYNC(S_AXIS_IARG_115_IS_ASYNC),
        .S_AXIS_IARG_116_IS_ASYNC(S_AXIS_IARG_116_IS_ASYNC),
        .S_AXIS_IARG_117_IS_ASYNC(S_AXIS_IARG_117_IS_ASYNC),
        .S_AXIS_IARG_118_IS_ASYNC(S_AXIS_IARG_118_IS_ASYNC),
        .S_AXIS_IARG_119_IS_ASYNC(S_AXIS_IARG_119_IS_ASYNC),
        .S_AXIS_IARG_120_IS_ASYNC(S_AXIS_IARG_120_IS_ASYNC),
        .S_AXIS_IARG_121_IS_ASYNC(S_AXIS_IARG_121_IS_ASYNC),
        .S_AXIS_IARG_122_IS_ASYNC(S_AXIS_IARG_122_IS_ASYNC),
        .S_AXIS_IARG_123_IS_ASYNC(S_AXIS_IARG_123_IS_ASYNC),
        .S_AXIS_IARG_124_IS_ASYNC(S_AXIS_IARG_124_IS_ASYNC),
        .S_AXIS_IARG_125_IS_ASYNC(S_AXIS_IARG_125_IS_ASYNC),
        .S_AXIS_IARG_126_IS_ASYNC(S_AXIS_IARG_126_IS_ASYNC),
        .S_AXIS_IARG_127_IS_ASYNC(S_AXIS_IARG_127_IS_ASYNC),
        .S_AXIS_IARG_0_DMWIDTH(S_AXIS_IARG_0_DMWIDTH),
        .S_AXIS_IARG_1_DMWIDTH(S_AXIS_IARG_1_DMWIDTH),
        .S_AXIS_IARG_2_DMWIDTH(S_AXIS_IARG_2_DMWIDTH),
        .S_AXIS_IARG_3_DMWIDTH(S_AXIS_IARG_3_DMWIDTH),
        .S_AXIS_IARG_4_DMWIDTH(S_AXIS_IARG_4_DMWIDTH),
        .S_AXIS_IARG_5_DMWIDTH(S_AXIS_IARG_5_DMWIDTH),
        .S_AXIS_IARG_6_DMWIDTH(S_AXIS_IARG_6_DMWIDTH),
        .S_AXIS_IARG_7_DMWIDTH(S_AXIS_IARG_7_DMWIDTH),
        .S_AXIS_IARG_8_DMWIDTH(S_AXIS_IARG_8_DMWIDTH),
        .S_AXIS_IARG_9_DMWIDTH(S_AXIS_IARG_9_DMWIDTH),
        .S_AXIS_IARG_10_DMWIDTH(S_AXIS_IARG_10_DMWIDTH),
        .S_AXIS_IARG_11_DMWIDTH(S_AXIS_IARG_11_DMWIDTH),
        .S_AXIS_IARG_12_DMWIDTH(S_AXIS_IARG_12_DMWIDTH),
        .S_AXIS_IARG_13_DMWIDTH(S_AXIS_IARG_13_DMWIDTH),
        .S_AXIS_IARG_14_DMWIDTH(S_AXIS_IARG_14_DMWIDTH),
        .S_AXIS_IARG_15_DMWIDTH(S_AXIS_IARG_15_DMWIDTH),
        .S_AXIS_IARG_16_DMWIDTH(S_AXIS_IARG_16_DMWIDTH),
        .S_AXIS_IARG_17_DMWIDTH(S_AXIS_IARG_17_DMWIDTH),
        .S_AXIS_IARG_18_DMWIDTH(S_AXIS_IARG_18_DMWIDTH),
        .S_AXIS_IARG_19_DMWIDTH(S_AXIS_IARG_19_DMWIDTH),
        .S_AXIS_IARG_20_DMWIDTH(S_AXIS_IARG_20_DMWIDTH),
        .S_AXIS_IARG_21_DMWIDTH(S_AXIS_IARG_21_DMWIDTH),
        .S_AXIS_IARG_22_DMWIDTH(S_AXIS_IARG_22_DMWIDTH),
        .S_AXIS_IARG_23_DMWIDTH(S_AXIS_IARG_23_DMWIDTH),
        .S_AXIS_IARG_24_DMWIDTH(S_AXIS_IARG_24_DMWIDTH),
        .S_AXIS_IARG_25_DMWIDTH(S_AXIS_IARG_25_DMWIDTH),
        .S_AXIS_IARG_26_DMWIDTH(S_AXIS_IARG_26_DMWIDTH),
        .S_AXIS_IARG_27_DMWIDTH(S_AXIS_IARG_27_DMWIDTH),
        .S_AXIS_IARG_28_DMWIDTH(S_AXIS_IARG_28_DMWIDTH),
        .S_AXIS_IARG_29_DMWIDTH(S_AXIS_IARG_29_DMWIDTH),
        .S_AXIS_IARG_30_DMWIDTH(S_AXIS_IARG_30_DMWIDTH),
        .S_AXIS_IARG_31_DMWIDTH(S_AXIS_IARG_31_DMWIDTH),
        .S_AXIS_IARG_32_DMWIDTH(S_AXIS_IARG_32_DMWIDTH),
        .S_AXIS_IARG_33_DMWIDTH(S_AXIS_IARG_33_DMWIDTH),
        .S_AXIS_IARG_34_DMWIDTH(S_AXIS_IARG_34_DMWIDTH),
        .S_AXIS_IARG_35_DMWIDTH(S_AXIS_IARG_35_DMWIDTH),
        .S_AXIS_IARG_36_DMWIDTH(S_AXIS_IARG_36_DMWIDTH),
        .S_AXIS_IARG_37_DMWIDTH(S_AXIS_IARG_37_DMWIDTH),
        .S_AXIS_IARG_38_DMWIDTH(S_AXIS_IARG_38_DMWIDTH),
        .S_AXIS_IARG_39_DMWIDTH(S_AXIS_IARG_39_DMWIDTH),
        .S_AXIS_IARG_40_DMWIDTH(S_AXIS_IARG_40_DMWIDTH),
        .S_AXIS_IARG_41_DMWIDTH(S_AXIS_IARG_41_DMWIDTH),
        .S_AXIS_IARG_42_DMWIDTH(S_AXIS_IARG_42_DMWIDTH),
        .S_AXIS_IARG_43_DMWIDTH(S_AXIS_IARG_43_DMWIDTH),
        .S_AXIS_IARG_44_DMWIDTH(S_AXIS_IARG_44_DMWIDTH),
        .S_AXIS_IARG_45_DMWIDTH(S_AXIS_IARG_45_DMWIDTH),
        .S_AXIS_IARG_46_DMWIDTH(S_AXIS_IARG_46_DMWIDTH),
        .S_AXIS_IARG_47_DMWIDTH(S_AXIS_IARG_47_DMWIDTH),
        .S_AXIS_IARG_48_DMWIDTH(S_AXIS_IARG_48_DMWIDTH),
        .S_AXIS_IARG_49_DMWIDTH(S_AXIS_IARG_49_DMWIDTH),
        .S_AXIS_IARG_50_DMWIDTH(S_AXIS_IARG_50_DMWIDTH),
        .S_AXIS_IARG_51_DMWIDTH(S_AXIS_IARG_51_DMWIDTH),
        .S_AXIS_IARG_52_DMWIDTH(S_AXIS_IARG_52_DMWIDTH),
        .S_AXIS_IARG_53_DMWIDTH(S_AXIS_IARG_53_DMWIDTH),
        .S_AXIS_IARG_54_DMWIDTH(S_AXIS_IARG_54_DMWIDTH),
        .S_AXIS_IARG_55_DMWIDTH(S_AXIS_IARG_55_DMWIDTH),
        .S_AXIS_IARG_56_DMWIDTH(S_AXIS_IARG_56_DMWIDTH),
        .S_AXIS_IARG_57_DMWIDTH(S_AXIS_IARG_57_DMWIDTH),
        .S_AXIS_IARG_58_DMWIDTH(S_AXIS_IARG_58_DMWIDTH),
        .S_AXIS_IARG_59_DMWIDTH(S_AXIS_IARG_59_DMWIDTH),
        .S_AXIS_IARG_60_DMWIDTH(S_AXIS_IARG_60_DMWIDTH),
        .S_AXIS_IARG_61_DMWIDTH(S_AXIS_IARG_61_DMWIDTH),
        .S_AXIS_IARG_62_DMWIDTH(S_AXIS_IARG_62_DMWIDTH),
        .S_AXIS_IARG_63_DMWIDTH(S_AXIS_IARG_63_DMWIDTH),
        .S_AXIS_IARG_64_DMWIDTH(S_AXIS_IARG_64_DMWIDTH),
        .S_AXIS_IARG_65_DMWIDTH(S_AXIS_IARG_65_DMWIDTH),
        .S_AXIS_IARG_66_DMWIDTH(S_AXIS_IARG_66_DMWIDTH),
        .S_AXIS_IARG_67_DMWIDTH(S_AXIS_IARG_67_DMWIDTH),
        .S_AXIS_IARG_68_DMWIDTH(S_AXIS_IARG_68_DMWIDTH),
        .S_AXIS_IARG_69_DMWIDTH(S_AXIS_IARG_69_DMWIDTH),
        .S_AXIS_IARG_70_DMWIDTH(S_AXIS_IARG_70_DMWIDTH),
        .S_AXIS_IARG_71_DMWIDTH(S_AXIS_IARG_71_DMWIDTH),
        .S_AXIS_IARG_72_DMWIDTH(S_AXIS_IARG_72_DMWIDTH),
        .S_AXIS_IARG_73_DMWIDTH(S_AXIS_IARG_73_DMWIDTH),
        .S_AXIS_IARG_74_DMWIDTH(S_AXIS_IARG_74_DMWIDTH),
        .S_AXIS_IARG_75_DMWIDTH(S_AXIS_IARG_75_DMWIDTH),
        .S_AXIS_IARG_76_DMWIDTH(S_AXIS_IARG_76_DMWIDTH),
        .S_AXIS_IARG_77_DMWIDTH(S_AXIS_IARG_77_DMWIDTH),
        .S_AXIS_IARG_78_DMWIDTH(S_AXIS_IARG_78_DMWIDTH),
        .S_AXIS_IARG_79_DMWIDTH(S_AXIS_IARG_79_DMWIDTH),
        .S_AXIS_IARG_80_DMWIDTH(S_AXIS_IARG_80_DMWIDTH),
        .S_AXIS_IARG_81_DMWIDTH(S_AXIS_IARG_81_DMWIDTH),
        .S_AXIS_IARG_82_DMWIDTH(S_AXIS_IARG_82_DMWIDTH),
        .S_AXIS_IARG_83_DMWIDTH(S_AXIS_IARG_83_DMWIDTH),
        .S_AXIS_IARG_84_DMWIDTH(S_AXIS_IARG_84_DMWIDTH),
        .S_AXIS_IARG_85_DMWIDTH(S_AXIS_IARG_85_DMWIDTH),
        .S_AXIS_IARG_86_DMWIDTH(S_AXIS_IARG_86_DMWIDTH),
        .S_AXIS_IARG_87_DMWIDTH(S_AXIS_IARG_87_DMWIDTH),
        .S_AXIS_IARG_88_DMWIDTH(S_AXIS_IARG_88_DMWIDTH),
        .S_AXIS_IARG_89_DMWIDTH(S_AXIS_IARG_89_DMWIDTH),
        .S_AXIS_IARG_90_DMWIDTH(S_AXIS_IARG_90_DMWIDTH),
        .S_AXIS_IARG_91_DMWIDTH(S_AXIS_IARG_91_DMWIDTH),
        .S_AXIS_IARG_92_DMWIDTH(S_AXIS_IARG_92_DMWIDTH),
        .S_AXIS_IARG_93_DMWIDTH(S_AXIS_IARG_93_DMWIDTH),
        .S_AXIS_IARG_94_DMWIDTH(S_AXIS_IARG_94_DMWIDTH),
        .S_AXIS_IARG_95_DMWIDTH(S_AXIS_IARG_95_DMWIDTH),
        .S_AXIS_IARG_96_DMWIDTH(S_AXIS_IARG_96_DMWIDTH),
        .S_AXIS_IARG_97_DMWIDTH(S_AXIS_IARG_97_DMWIDTH),
        .S_AXIS_IARG_98_DMWIDTH(S_AXIS_IARG_98_DMWIDTH),
        .S_AXIS_IARG_99_DMWIDTH(S_AXIS_IARG_99_DMWIDTH),
        .S_AXIS_IARG_100_DMWIDTH(S_AXIS_IARG_100_DMWIDTH),
        .S_AXIS_IARG_101_DMWIDTH(S_AXIS_IARG_101_DMWIDTH),
        .S_AXIS_IARG_102_DMWIDTH(S_AXIS_IARG_102_DMWIDTH),
        .S_AXIS_IARG_103_DMWIDTH(S_AXIS_IARG_103_DMWIDTH),
        .S_AXIS_IARG_104_DMWIDTH(S_AXIS_IARG_104_DMWIDTH),
        .S_AXIS_IARG_105_DMWIDTH(S_AXIS_IARG_105_DMWIDTH),
        .S_AXIS_IARG_106_DMWIDTH(S_AXIS_IARG_106_DMWIDTH),
        .S_AXIS_IARG_107_DMWIDTH(S_AXIS_IARG_107_DMWIDTH),
        .S_AXIS_IARG_108_DMWIDTH(S_AXIS_IARG_108_DMWIDTH),
        .S_AXIS_IARG_109_DMWIDTH(S_AXIS_IARG_109_DMWIDTH),
        .S_AXIS_IARG_110_DMWIDTH(S_AXIS_IARG_110_DMWIDTH),
        .S_AXIS_IARG_111_DMWIDTH(S_AXIS_IARG_111_DMWIDTH),
        .S_AXIS_IARG_112_DMWIDTH(S_AXIS_IARG_112_DMWIDTH),
        .S_AXIS_IARG_113_DMWIDTH(S_AXIS_IARG_113_DMWIDTH),
        .S_AXIS_IARG_114_DMWIDTH(S_AXIS_IARG_114_DMWIDTH),
        .S_AXIS_IARG_115_DMWIDTH(S_AXIS_IARG_115_DMWIDTH),
        .S_AXIS_IARG_116_DMWIDTH(S_AXIS_IARG_116_DMWIDTH),
        .S_AXIS_IARG_117_DMWIDTH(S_AXIS_IARG_117_DMWIDTH),
        .S_AXIS_IARG_118_DMWIDTH(S_AXIS_IARG_118_DMWIDTH),
        .S_AXIS_IARG_119_DMWIDTH(S_AXIS_IARG_119_DMWIDTH),
        .S_AXIS_IARG_120_DMWIDTH(S_AXIS_IARG_120_DMWIDTH),
        .S_AXIS_IARG_121_DMWIDTH(S_AXIS_IARG_121_DMWIDTH),
        .S_AXIS_IARG_122_DMWIDTH(S_AXIS_IARG_122_DMWIDTH),
        .S_AXIS_IARG_123_DMWIDTH(S_AXIS_IARG_123_DMWIDTH),
        .S_AXIS_IARG_124_DMWIDTH(S_AXIS_IARG_124_DMWIDTH),
        .S_AXIS_IARG_125_DMWIDTH(S_AXIS_IARG_125_DMWIDTH),
        .S_AXIS_IARG_126_DMWIDTH(S_AXIS_IARG_126_DMWIDTH),
        .S_AXIS_IARG_127_DMWIDTH(S_AXIS_IARG_127_DMWIDTH)
    ) in_axis_args_i (
        .acc_clk(acc_aclk),
        .acc_aresetn(acc_aresetn),
        .in_axis_allow(inaxis_ctrl_allow),
        .s_axis_iarg_0_aclk(s_axis_iarg_0_aclk),
        .s_axis_iarg_0_aresetn(s_axis_iarg_0_aresetn),
        .s_axis_iarg_0_tlast(s_axis_iarg_0_tlast),
        .s_axis_iarg_0_tvalid(s_axis_iarg_0_tvalid),
        .s_axis_iarg_0_tkeep(s_axis_iarg_0_tkeep),
        .s_axis_iarg_0_tstrb(s_axis_iarg_0_tstrb),
        .s_axis_iarg_0_tdata(s_axis_iarg_0_tdata),
        .s_axis_iarg_0_tready(s_axis_iarg_0_tready),
        .ap_axis_iarg_0_tlast(ap_axis_iarg_0_tlast),
        .ap_axis_iarg_0_tvalid(ap_axis_iarg_0_tvalid),
        .ap_axis_iarg_0_tkeep(ap_axis_iarg_0_tkeep),
        .ap_axis_iarg_0_tstrb(ap_axis_iarg_0_tstrb),
        .ap_axis_iarg_0_tdata(ap_axis_iarg_0_tdata),
        .ap_axis_iarg_0_tready(ap_axis_iarg_0_tready),
        .s_axis_iarg_1_aclk(s_axis_iarg_1_aclk),
        .s_axis_iarg_1_aresetn(s_axis_iarg_1_aresetn),
        .s_axis_iarg_1_tlast(s_axis_iarg_1_tlast),
        .s_axis_iarg_1_tvalid(s_axis_iarg_1_tvalid),
        .s_axis_iarg_1_tkeep(s_axis_iarg_1_tkeep),
        .s_axis_iarg_1_tstrb(s_axis_iarg_1_tstrb),
        .s_axis_iarg_1_tdata(s_axis_iarg_1_tdata),
        .s_axis_iarg_1_tready(s_axis_iarg_1_tready),
        .ap_axis_iarg_1_tlast(ap_axis_iarg_1_tlast),
        .ap_axis_iarg_1_tvalid(ap_axis_iarg_1_tvalid),
        .ap_axis_iarg_1_tkeep(ap_axis_iarg_1_tkeep),
        .ap_axis_iarg_1_tstrb(ap_axis_iarg_1_tstrb),
        .ap_axis_iarg_1_tdata(ap_axis_iarg_1_tdata),
        .ap_axis_iarg_1_tready(ap_axis_iarg_1_tready),
        .s_axis_iarg_2_aclk(s_axis_iarg_2_aclk),
        .s_axis_iarg_2_aresetn(s_axis_iarg_2_aresetn),
        .s_axis_iarg_2_tlast(s_axis_iarg_2_tlast),
        .s_axis_iarg_2_tvalid(s_axis_iarg_2_tvalid),
        .s_axis_iarg_2_tkeep(s_axis_iarg_2_tkeep),
        .s_axis_iarg_2_tstrb(s_axis_iarg_2_tstrb),
        .s_axis_iarg_2_tdata(s_axis_iarg_2_tdata),
        .s_axis_iarg_2_tready(s_axis_iarg_2_tready),
        .ap_axis_iarg_2_tlast(ap_axis_iarg_2_tlast),
        .ap_axis_iarg_2_tvalid(ap_axis_iarg_2_tvalid),
        .ap_axis_iarg_2_tkeep(ap_axis_iarg_2_tkeep),
        .ap_axis_iarg_2_tstrb(ap_axis_iarg_2_tstrb),
        .ap_axis_iarg_2_tdata(ap_axis_iarg_2_tdata),
        .ap_axis_iarg_2_tready(ap_axis_iarg_2_tready),
        .s_axis_iarg_3_aclk(s_axis_iarg_3_aclk),
        .s_axis_iarg_3_aresetn(s_axis_iarg_3_aresetn),
        .s_axis_iarg_3_tlast(s_axis_iarg_3_tlast),
        .s_axis_iarg_3_tvalid(s_axis_iarg_3_tvalid),
        .s_axis_iarg_3_tkeep(s_axis_iarg_3_tkeep),
        .s_axis_iarg_3_tstrb(s_axis_iarg_3_tstrb),
        .s_axis_iarg_3_tdata(s_axis_iarg_3_tdata),
        .s_axis_iarg_3_tready(s_axis_iarg_3_tready),
        .ap_axis_iarg_3_tlast(ap_axis_iarg_3_tlast),
        .ap_axis_iarg_3_tvalid(ap_axis_iarg_3_tvalid),
        .ap_axis_iarg_3_tkeep(ap_axis_iarg_3_tkeep),
        .ap_axis_iarg_3_tstrb(ap_axis_iarg_3_tstrb),
        .ap_axis_iarg_3_tdata(ap_axis_iarg_3_tdata),
        .ap_axis_iarg_3_tready(ap_axis_iarg_3_tready),
        .s_axis_iarg_4_aclk(s_axis_iarg_4_aclk),
        .s_axis_iarg_4_aresetn(s_axis_iarg_4_aresetn),
        .s_axis_iarg_4_tlast(s_axis_iarg_4_tlast),
        .s_axis_iarg_4_tvalid(s_axis_iarg_4_tvalid),
        .s_axis_iarg_4_tkeep(s_axis_iarg_4_tkeep),
        .s_axis_iarg_4_tstrb(s_axis_iarg_4_tstrb),
        .s_axis_iarg_4_tdata(s_axis_iarg_4_tdata),
        .s_axis_iarg_4_tready(s_axis_iarg_4_tready),
        .ap_axis_iarg_4_tlast(ap_axis_iarg_4_tlast),
        .ap_axis_iarg_4_tvalid(ap_axis_iarg_4_tvalid),
        .ap_axis_iarg_4_tkeep(ap_axis_iarg_4_tkeep),
        .ap_axis_iarg_4_tstrb(ap_axis_iarg_4_tstrb),
        .ap_axis_iarg_4_tdata(ap_axis_iarg_4_tdata),
        .ap_axis_iarg_4_tready(ap_axis_iarg_4_tready),
        .s_axis_iarg_5_aclk(s_axis_iarg_5_aclk),
        .s_axis_iarg_5_aresetn(s_axis_iarg_5_aresetn),
        .s_axis_iarg_5_tlast(s_axis_iarg_5_tlast),
        .s_axis_iarg_5_tvalid(s_axis_iarg_5_tvalid),
        .s_axis_iarg_5_tkeep(s_axis_iarg_5_tkeep),
        .s_axis_iarg_5_tstrb(s_axis_iarg_5_tstrb),
        .s_axis_iarg_5_tdata(s_axis_iarg_5_tdata),
        .s_axis_iarg_5_tready(s_axis_iarg_5_tready),
        .ap_axis_iarg_5_tlast(ap_axis_iarg_5_tlast),
        .ap_axis_iarg_5_tvalid(ap_axis_iarg_5_tvalid),
        .ap_axis_iarg_5_tkeep(ap_axis_iarg_5_tkeep),
        .ap_axis_iarg_5_tstrb(ap_axis_iarg_5_tstrb),
        .ap_axis_iarg_5_tdata(ap_axis_iarg_5_tdata),
        .ap_axis_iarg_5_tready(ap_axis_iarg_5_tready),
        .s_axis_iarg_6_aclk(s_axis_iarg_6_aclk),
        .s_axis_iarg_6_aresetn(s_axis_iarg_6_aresetn),
        .s_axis_iarg_6_tlast(s_axis_iarg_6_tlast),
        .s_axis_iarg_6_tvalid(s_axis_iarg_6_tvalid),
        .s_axis_iarg_6_tkeep(s_axis_iarg_6_tkeep),
        .s_axis_iarg_6_tstrb(s_axis_iarg_6_tstrb),
        .s_axis_iarg_6_tdata(s_axis_iarg_6_tdata),
        .s_axis_iarg_6_tready(s_axis_iarg_6_tready),
        .ap_axis_iarg_6_tlast(ap_axis_iarg_6_tlast),
        .ap_axis_iarg_6_tvalid(ap_axis_iarg_6_tvalid),
        .ap_axis_iarg_6_tkeep(ap_axis_iarg_6_tkeep),
        .ap_axis_iarg_6_tstrb(ap_axis_iarg_6_tstrb),
        .ap_axis_iarg_6_tdata(ap_axis_iarg_6_tdata),
        .ap_axis_iarg_6_tready(ap_axis_iarg_6_tready),
        .s_axis_iarg_7_aclk(s_axis_iarg_7_aclk),
        .s_axis_iarg_7_aresetn(s_axis_iarg_7_aresetn),
        .s_axis_iarg_7_tlast(s_axis_iarg_7_tlast),
        .s_axis_iarg_7_tvalid(s_axis_iarg_7_tvalid),
        .s_axis_iarg_7_tkeep(s_axis_iarg_7_tkeep),
        .s_axis_iarg_7_tstrb(s_axis_iarg_7_tstrb),
        .s_axis_iarg_7_tdata(s_axis_iarg_7_tdata),
        .s_axis_iarg_7_tready(s_axis_iarg_7_tready),
        .ap_axis_iarg_7_tlast(ap_axis_iarg_7_tlast),
        .ap_axis_iarg_7_tvalid(ap_axis_iarg_7_tvalid),
        .ap_axis_iarg_7_tkeep(ap_axis_iarg_7_tkeep),
        .ap_axis_iarg_7_tstrb(ap_axis_iarg_7_tstrb),
        .ap_axis_iarg_7_tdata(ap_axis_iarg_7_tdata),
        .ap_axis_iarg_7_tready(ap_axis_iarg_7_tready),
        .s_axis_iarg_8_aclk(s_axis_iarg_8_aclk),
        .s_axis_iarg_8_aresetn(s_axis_iarg_8_aresetn),
        .s_axis_iarg_8_tlast(s_axis_iarg_8_tlast),
        .s_axis_iarg_8_tvalid(s_axis_iarg_8_tvalid),
        .s_axis_iarg_8_tkeep(s_axis_iarg_8_tkeep),
        .s_axis_iarg_8_tstrb(s_axis_iarg_8_tstrb),
        .s_axis_iarg_8_tdata(s_axis_iarg_8_tdata),
        .s_axis_iarg_8_tready(s_axis_iarg_8_tready),
        .ap_axis_iarg_8_tlast(ap_axis_iarg_8_tlast),
        .ap_axis_iarg_8_tvalid(ap_axis_iarg_8_tvalid),
        .ap_axis_iarg_8_tkeep(ap_axis_iarg_8_tkeep),
        .ap_axis_iarg_8_tstrb(ap_axis_iarg_8_tstrb),
        .ap_axis_iarg_8_tdata(ap_axis_iarg_8_tdata),
        .ap_axis_iarg_8_tready(ap_axis_iarg_8_tready),
        .s_axis_iarg_9_aclk(s_axis_iarg_9_aclk),
        .s_axis_iarg_9_aresetn(s_axis_iarg_9_aresetn),
        .s_axis_iarg_9_tlast(s_axis_iarg_9_tlast),
        .s_axis_iarg_9_tvalid(s_axis_iarg_9_tvalid),
        .s_axis_iarg_9_tkeep(s_axis_iarg_9_tkeep),
        .s_axis_iarg_9_tstrb(s_axis_iarg_9_tstrb),
        .s_axis_iarg_9_tdata(s_axis_iarg_9_tdata),
        .s_axis_iarg_9_tready(s_axis_iarg_9_tready),
        .ap_axis_iarg_9_tlast(ap_axis_iarg_9_tlast),
        .ap_axis_iarg_9_tvalid(ap_axis_iarg_9_tvalid),
        .ap_axis_iarg_9_tkeep(ap_axis_iarg_9_tkeep),
        .ap_axis_iarg_9_tstrb(ap_axis_iarg_9_tstrb),
        .ap_axis_iarg_9_tdata(ap_axis_iarg_9_tdata),
        .ap_axis_iarg_9_tready(ap_axis_iarg_9_tready),
        .s_axis_iarg_10_aclk(s_axis_iarg_10_aclk),
        .s_axis_iarg_10_aresetn(s_axis_iarg_10_aresetn),
        .s_axis_iarg_10_tlast(s_axis_iarg_10_tlast),
        .s_axis_iarg_10_tvalid(s_axis_iarg_10_tvalid),
        .s_axis_iarg_10_tkeep(s_axis_iarg_10_tkeep),
        .s_axis_iarg_10_tstrb(s_axis_iarg_10_tstrb),
        .s_axis_iarg_10_tdata(s_axis_iarg_10_tdata),
        .s_axis_iarg_10_tready(s_axis_iarg_10_tready),
        .ap_axis_iarg_10_tlast(ap_axis_iarg_10_tlast),
        .ap_axis_iarg_10_tvalid(ap_axis_iarg_10_tvalid),
        .ap_axis_iarg_10_tkeep(ap_axis_iarg_10_tkeep),
        .ap_axis_iarg_10_tstrb(ap_axis_iarg_10_tstrb),
        .ap_axis_iarg_10_tdata(ap_axis_iarg_10_tdata),
        .ap_axis_iarg_10_tready(ap_axis_iarg_10_tready),
        .s_axis_iarg_11_aclk(s_axis_iarg_11_aclk),
        .s_axis_iarg_11_aresetn(s_axis_iarg_11_aresetn),
        .s_axis_iarg_11_tlast(s_axis_iarg_11_tlast),
        .s_axis_iarg_11_tvalid(s_axis_iarg_11_tvalid),
        .s_axis_iarg_11_tkeep(s_axis_iarg_11_tkeep),
        .s_axis_iarg_11_tstrb(s_axis_iarg_11_tstrb),
        .s_axis_iarg_11_tdata(s_axis_iarg_11_tdata),
        .s_axis_iarg_11_tready(s_axis_iarg_11_tready),
        .ap_axis_iarg_11_tlast(ap_axis_iarg_11_tlast),
        .ap_axis_iarg_11_tvalid(ap_axis_iarg_11_tvalid),
        .ap_axis_iarg_11_tkeep(ap_axis_iarg_11_tkeep),
        .ap_axis_iarg_11_tstrb(ap_axis_iarg_11_tstrb),
        .ap_axis_iarg_11_tdata(ap_axis_iarg_11_tdata),
        .ap_axis_iarg_11_tready(ap_axis_iarg_11_tready),
        .s_axis_iarg_12_aclk(s_axis_iarg_12_aclk),
        .s_axis_iarg_12_aresetn(s_axis_iarg_12_aresetn),
        .s_axis_iarg_12_tlast(s_axis_iarg_12_tlast),
        .s_axis_iarg_12_tvalid(s_axis_iarg_12_tvalid),
        .s_axis_iarg_12_tkeep(s_axis_iarg_12_tkeep),
        .s_axis_iarg_12_tstrb(s_axis_iarg_12_tstrb),
        .s_axis_iarg_12_tdata(s_axis_iarg_12_tdata),
        .s_axis_iarg_12_tready(s_axis_iarg_12_tready),
        .ap_axis_iarg_12_tlast(ap_axis_iarg_12_tlast),
        .ap_axis_iarg_12_tvalid(ap_axis_iarg_12_tvalid),
        .ap_axis_iarg_12_tkeep(ap_axis_iarg_12_tkeep),
        .ap_axis_iarg_12_tstrb(ap_axis_iarg_12_tstrb),
        .ap_axis_iarg_12_tdata(ap_axis_iarg_12_tdata),
        .ap_axis_iarg_12_tready(ap_axis_iarg_12_tready),
        .s_axis_iarg_13_aclk(s_axis_iarg_13_aclk),
        .s_axis_iarg_13_aresetn(s_axis_iarg_13_aresetn),
        .s_axis_iarg_13_tlast(s_axis_iarg_13_tlast),
        .s_axis_iarg_13_tvalid(s_axis_iarg_13_tvalid),
        .s_axis_iarg_13_tkeep(s_axis_iarg_13_tkeep),
        .s_axis_iarg_13_tstrb(s_axis_iarg_13_tstrb),
        .s_axis_iarg_13_tdata(s_axis_iarg_13_tdata),
        .s_axis_iarg_13_tready(s_axis_iarg_13_tready),
        .ap_axis_iarg_13_tlast(ap_axis_iarg_13_tlast),
        .ap_axis_iarg_13_tvalid(ap_axis_iarg_13_tvalid),
        .ap_axis_iarg_13_tkeep(ap_axis_iarg_13_tkeep),
        .ap_axis_iarg_13_tstrb(ap_axis_iarg_13_tstrb),
        .ap_axis_iarg_13_tdata(ap_axis_iarg_13_tdata),
        .ap_axis_iarg_13_tready(ap_axis_iarg_13_tready),
        .s_axis_iarg_14_aclk(s_axis_iarg_14_aclk),
        .s_axis_iarg_14_aresetn(s_axis_iarg_14_aresetn),
        .s_axis_iarg_14_tlast(s_axis_iarg_14_tlast),
        .s_axis_iarg_14_tvalid(s_axis_iarg_14_tvalid),
        .s_axis_iarg_14_tkeep(s_axis_iarg_14_tkeep),
        .s_axis_iarg_14_tstrb(s_axis_iarg_14_tstrb),
        .s_axis_iarg_14_tdata(s_axis_iarg_14_tdata),
        .s_axis_iarg_14_tready(s_axis_iarg_14_tready),
        .ap_axis_iarg_14_tlast(ap_axis_iarg_14_tlast),
        .ap_axis_iarg_14_tvalid(ap_axis_iarg_14_tvalid),
        .ap_axis_iarg_14_tkeep(ap_axis_iarg_14_tkeep),
        .ap_axis_iarg_14_tstrb(ap_axis_iarg_14_tstrb),
        .ap_axis_iarg_14_tdata(ap_axis_iarg_14_tdata),
        .ap_axis_iarg_14_tready(ap_axis_iarg_14_tready),
        .s_axis_iarg_15_aclk(s_axis_iarg_15_aclk),
        .s_axis_iarg_15_aresetn(s_axis_iarg_15_aresetn),
        .s_axis_iarg_15_tlast(s_axis_iarg_15_tlast),
        .s_axis_iarg_15_tvalid(s_axis_iarg_15_tvalid),
        .s_axis_iarg_15_tkeep(s_axis_iarg_15_tkeep),
        .s_axis_iarg_15_tstrb(s_axis_iarg_15_tstrb),
        .s_axis_iarg_15_tdata(s_axis_iarg_15_tdata),
        .s_axis_iarg_15_tready(s_axis_iarg_15_tready),
        .ap_axis_iarg_15_tlast(ap_axis_iarg_15_tlast),
        .ap_axis_iarg_15_tvalid(ap_axis_iarg_15_tvalid),
        .ap_axis_iarg_15_tkeep(ap_axis_iarg_15_tkeep),
        .ap_axis_iarg_15_tstrb(ap_axis_iarg_15_tstrb),
        .ap_axis_iarg_15_tdata(ap_axis_iarg_15_tdata),
        .ap_axis_iarg_15_tready(ap_axis_iarg_15_tready),
        .s_axis_iarg_16_aclk(s_axis_iarg_16_aclk),
        .s_axis_iarg_16_aresetn(s_axis_iarg_16_aresetn),
        .s_axis_iarg_16_tlast(s_axis_iarg_16_tlast),
        .s_axis_iarg_16_tvalid(s_axis_iarg_16_tvalid),
        .s_axis_iarg_16_tkeep(s_axis_iarg_16_tkeep),
        .s_axis_iarg_16_tstrb(s_axis_iarg_16_tstrb),
        .s_axis_iarg_16_tdata(s_axis_iarg_16_tdata),
        .s_axis_iarg_16_tready(s_axis_iarg_16_tready),
        .ap_axis_iarg_16_tlast(ap_axis_iarg_16_tlast),
        .ap_axis_iarg_16_tvalid(ap_axis_iarg_16_tvalid),
        .ap_axis_iarg_16_tkeep(ap_axis_iarg_16_tkeep),
        .ap_axis_iarg_16_tstrb(ap_axis_iarg_16_tstrb),
        .ap_axis_iarg_16_tdata(ap_axis_iarg_16_tdata),
        .ap_axis_iarg_16_tready(ap_axis_iarg_16_tready),
        .s_axis_iarg_17_aclk(s_axis_iarg_17_aclk),
        .s_axis_iarg_17_aresetn(s_axis_iarg_17_aresetn),
        .s_axis_iarg_17_tlast(s_axis_iarg_17_tlast),
        .s_axis_iarg_17_tvalid(s_axis_iarg_17_tvalid),
        .s_axis_iarg_17_tkeep(s_axis_iarg_17_tkeep),
        .s_axis_iarg_17_tstrb(s_axis_iarg_17_tstrb),
        .s_axis_iarg_17_tdata(s_axis_iarg_17_tdata),
        .s_axis_iarg_17_tready(s_axis_iarg_17_tready),
        .ap_axis_iarg_17_tlast(ap_axis_iarg_17_tlast),
        .ap_axis_iarg_17_tvalid(ap_axis_iarg_17_tvalid),
        .ap_axis_iarg_17_tkeep(ap_axis_iarg_17_tkeep),
        .ap_axis_iarg_17_tstrb(ap_axis_iarg_17_tstrb),
        .ap_axis_iarg_17_tdata(ap_axis_iarg_17_tdata),
        .ap_axis_iarg_17_tready(ap_axis_iarg_17_tready),
        .s_axis_iarg_18_aclk(s_axis_iarg_18_aclk),
        .s_axis_iarg_18_aresetn(s_axis_iarg_18_aresetn),
        .s_axis_iarg_18_tlast(s_axis_iarg_18_tlast),
        .s_axis_iarg_18_tvalid(s_axis_iarg_18_tvalid),
        .s_axis_iarg_18_tkeep(s_axis_iarg_18_tkeep),
        .s_axis_iarg_18_tstrb(s_axis_iarg_18_tstrb),
        .s_axis_iarg_18_tdata(s_axis_iarg_18_tdata),
        .s_axis_iarg_18_tready(s_axis_iarg_18_tready),
        .ap_axis_iarg_18_tlast(ap_axis_iarg_18_tlast),
        .ap_axis_iarg_18_tvalid(ap_axis_iarg_18_tvalid),
        .ap_axis_iarg_18_tkeep(ap_axis_iarg_18_tkeep),
        .ap_axis_iarg_18_tstrb(ap_axis_iarg_18_tstrb),
        .ap_axis_iarg_18_tdata(ap_axis_iarg_18_tdata),
        .ap_axis_iarg_18_tready(ap_axis_iarg_18_tready),
        .s_axis_iarg_19_aclk(s_axis_iarg_19_aclk),
        .s_axis_iarg_19_aresetn(s_axis_iarg_19_aresetn),
        .s_axis_iarg_19_tlast(s_axis_iarg_19_tlast),
        .s_axis_iarg_19_tvalid(s_axis_iarg_19_tvalid),
        .s_axis_iarg_19_tkeep(s_axis_iarg_19_tkeep),
        .s_axis_iarg_19_tstrb(s_axis_iarg_19_tstrb),
        .s_axis_iarg_19_tdata(s_axis_iarg_19_tdata),
        .s_axis_iarg_19_tready(s_axis_iarg_19_tready),
        .ap_axis_iarg_19_tlast(ap_axis_iarg_19_tlast),
        .ap_axis_iarg_19_tvalid(ap_axis_iarg_19_tvalid),
        .ap_axis_iarg_19_tkeep(ap_axis_iarg_19_tkeep),
        .ap_axis_iarg_19_tstrb(ap_axis_iarg_19_tstrb),
        .ap_axis_iarg_19_tdata(ap_axis_iarg_19_tdata),
        .ap_axis_iarg_19_tready(ap_axis_iarg_19_tready),
        .s_axis_iarg_20_aclk(s_axis_iarg_20_aclk),
        .s_axis_iarg_20_aresetn(s_axis_iarg_20_aresetn),
        .s_axis_iarg_20_tlast(s_axis_iarg_20_tlast),
        .s_axis_iarg_20_tvalid(s_axis_iarg_20_tvalid),
        .s_axis_iarg_20_tkeep(s_axis_iarg_20_tkeep),
        .s_axis_iarg_20_tstrb(s_axis_iarg_20_tstrb),
        .s_axis_iarg_20_tdata(s_axis_iarg_20_tdata),
        .s_axis_iarg_20_tready(s_axis_iarg_20_tready),
        .ap_axis_iarg_20_tlast(ap_axis_iarg_20_tlast),
        .ap_axis_iarg_20_tvalid(ap_axis_iarg_20_tvalid),
        .ap_axis_iarg_20_tkeep(ap_axis_iarg_20_tkeep),
        .ap_axis_iarg_20_tstrb(ap_axis_iarg_20_tstrb),
        .ap_axis_iarg_20_tdata(ap_axis_iarg_20_tdata),
        .ap_axis_iarg_20_tready(ap_axis_iarg_20_tready),
        .s_axis_iarg_21_aclk(s_axis_iarg_21_aclk),
        .s_axis_iarg_21_aresetn(s_axis_iarg_21_aresetn),
        .s_axis_iarg_21_tlast(s_axis_iarg_21_tlast),
        .s_axis_iarg_21_tvalid(s_axis_iarg_21_tvalid),
        .s_axis_iarg_21_tkeep(s_axis_iarg_21_tkeep),
        .s_axis_iarg_21_tstrb(s_axis_iarg_21_tstrb),
        .s_axis_iarg_21_tdata(s_axis_iarg_21_tdata),
        .s_axis_iarg_21_tready(s_axis_iarg_21_tready),
        .ap_axis_iarg_21_tlast(ap_axis_iarg_21_tlast),
        .ap_axis_iarg_21_tvalid(ap_axis_iarg_21_tvalid),
        .ap_axis_iarg_21_tkeep(ap_axis_iarg_21_tkeep),
        .ap_axis_iarg_21_tstrb(ap_axis_iarg_21_tstrb),
        .ap_axis_iarg_21_tdata(ap_axis_iarg_21_tdata),
        .ap_axis_iarg_21_tready(ap_axis_iarg_21_tready),
        .s_axis_iarg_22_aclk(s_axis_iarg_22_aclk),
        .s_axis_iarg_22_aresetn(s_axis_iarg_22_aresetn),
        .s_axis_iarg_22_tlast(s_axis_iarg_22_tlast),
        .s_axis_iarg_22_tvalid(s_axis_iarg_22_tvalid),
        .s_axis_iarg_22_tkeep(s_axis_iarg_22_tkeep),
        .s_axis_iarg_22_tstrb(s_axis_iarg_22_tstrb),
        .s_axis_iarg_22_tdata(s_axis_iarg_22_tdata),
        .s_axis_iarg_22_tready(s_axis_iarg_22_tready),
        .ap_axis_iarg_22_tlast(ap_axis_iarg_22_tlast),
        .ap_axis_iarg_22_tvalid(ap_axis_iarg_22_tvalid),
        .ap_axis_iarg_22_tkeep(ap_axis_iarg_22_tkeep),
        .ap_axis_iarg_22_tstrb(ap_axis_iarg_22_tstrb),
        .ap_axis_iarg_22_tdata(ap_axis_iarg_22_tdata),
        .ap_axis_iarg_22_tready(ap_axis_iarg_22_tready),
        .s_axis_iarg_23_aclk(s_axis_iarg_23_aclk),
        .s_axis_iarg_23_aresetn(s_axis_iarg_23_aresetn),
        .s_axis_iarg_23_tlast(s_axis_iarg_23_tlast),
        .s_axis_iarg_23_tvalid(s_axis_iarg_23_tvalid),
        .s_axis_iarg_23_tkeep(s_axis_iarg_23_tkeep),
        .s_axis_iarg_23_tstrb(s_axis_iarg_23_tstrb),
        .s_axis_iarg_23_tdata(s_axis_iarg_23_tdata),
        .s_axis_iarg_23_tready(s_axis_iarg_23_tready),
        .ap_axis_iarg_23_tlast(ap_axis_iarg_23_tlast),
        .ap_axis_iarg_23_tvalid(ap_axis_iarg_23_tvalid),
        .ap_axis_iarg_23_tkeep(ap_axis_iarg_23_tkeep),
        .ap_axis_iarg_23_tstrb(ap_axis_iarg_23_tstrb),
        .ap_axis_iarg_23_tdata(ap_axis_iarg_23_tdata),
        .ap_axis_iarg_23_tready(ap_axis_iarg_23_tready),
        .s_axis_iarg_24_aclk(s_axis_iarg_24_aclk),
        .s_axis_iarg_24_aresetn(s_axis_iarg_24_aresetn),
        .s_axis_iarg_24_tlast(s_axis_iarg_24_tlast),
        .s_axis_iarg_24_tvalid(s_axis_iarg_24_tvalid),
        .s_axis_iarg_24_tkeep(s_axis_iarg_24_tkeep),
        .s_axis_iarg_24_tstrb(s_axis_iarg_24_tstrb),
        .s_axis_iarg_24_tdata(s_axis_iarg_24_tdata),
        .s_axis_iarg_24_tready(s_axis_iarg_24_tready),
        .ap_axis_iarg_24_tlast(ap_axis_iarg_24_tlast),
        .ap_axis_iarg_24_tvalid(ap_axis_iarg_24_tvalid),
        .ap_axis_iarg_24_tkeep(ap_axis_iarg_24_tkeep),
        .ap_axis_iarg_24_tstrb(ap_axis_iarg_24_tstrb),
        .ap_axis_iarg_24_tdata(ap_axis_iarg_24_tdata),
        .ap_axis_iarg_24_tready(ap_axis_iarg_24_tready),
        .s_axis_iarg_25_aclk(s_axis_iarg_25_aclk),
        .s_axis_iarg_25_aresetn(s_axis_iarg_25_aresetn),
        .s_axis_iarg_25_tlast(s_axis_iarg_25_tlast),
        .s_axis_iarg_25_tvalid(s_axis_iarg_25_tvalid),
        .s_axis_iarg_25_tkeep(s_axis_iarg_25_tkeep),
        .s_axis_iarg_25_tstrb(s_axis_iarg_25_tstrb),
        .s_axis_iarg_25_tdata(s_axis_iarg_25_tdata),
        .s_axis_iarg_25_tready(s_axis_iarg_25_tready),
        .ap_axis_iarg_25_tlast(ap_axis_iarg_25_tlast),
        .ap_axis_iarg_25_tvalid(ap_axis_iarg_25_tvalid),
        .ap_axis_iarg_25_tkeep(ap_axis_iarg_25_tkeep),
        .ap_axis_iarg_25_tstrb(ap_axis_iarg_25_tstrb),
        .ap_axis_iarg_25_tdata(ap_axis_iarg_25_tdata),
        .ap_axis_iarg_25_tready(ap_axis_iarg_25_tready),
        .s_axis_iarg_26_aclk(s_axis_iarg_26_aclk),
        .s_axis_iarg_26_aresetn(s_axis_iarg_26_aresetn),
        .s_axis_iarg_26_tlast(s_axis_iarg_26_tlast),
        .s_axis_iarg_26_tvalid(s_axis_iarg_26_tvalid),
        .s_axis_iarg_26_tkeep(s_axis_iarg_26_tkeep),
        .s_axis_iarg_26_tstrb(s_axis_iarg_26_tstrb),
        .s_axis_iarg_26_tdata(s_axis_iarg_26_tdata),
        .s_axis_iarg_26_tready(s_axis_iarg_26_tready),
        .ap_axis_iarg_26_tlast(ap_axis_iarg_26_tlast),
        .ap_axis_iarg_26_tvalid(ap_axis_iarg_26_tvalid),
        .ap_axis_iarg_26_tkeep(ap_axis_iarg_26_tkeep),
        .ap_axis_iarg_26_tstrb(ap_axis_iarg_26_tstrb),
        .ap_axis_iarg_26_tdata(ap_axis_iarg_26_tdata),
        .ap_axis_iarg_26_tready(ap_axis_iarg_26_tready),
        .s_axis_iarg_27_aclk(s_axis_iarg_27_aclk),
        .s_axis_iarg_27_aresetn(s_axis_iarg_27_aresetn),
        .s_axis_iarg_27_tlast(s_axis_iarg_27_tlast),
        .s_axis_iarg_27_tvalid(s_axis_iarg_27_tvalid),
        .s_axis_iarg_27_tkeep(s_axis_iarg_27_tkeep),
        .s_axis_iarg_27_tstrb(s_axis_iarg_27_tstrb),
        .s_axis_iarg_27_tdata(s_axis_iarg_27_tdata),
        .s_axis_iarg_27_tready(s_axis_iarg_27_tready),
        .ap_axis_iarg_27_tlast(ap_axis_iarg_27_tlast),
        .ap_axis_iarg_27_tvalid(ap_axis_iarg_27_tvalid),
        .ap_axis_iarg_27_tkeep(ap_axis_iarg_27_tkeep),
        .ap_axis_iarg_27_tstrb(ap_axis_iarg_27_tstrb),
        .ap_axis_iarg_27_tdata(ap_axis_iarg_27_tdata),
        .ap_axis_iarg_27_tready(ap_axis_iarg_27_tready),
        .s_axis_iarg_28_aclk(s_axis_iarg_28_aclk),
        .s_axis_iarg_28_aresetn(s_axis_iarg_28_aresetn),
        .s_axis_iarg_28_tlast(s_axis_iarg_28_tlast),
        .s_axis_iarg_28_tvalid(s_axis_iarg_28_tvalid),
        .s_axis_iarg_28_tkeep(s_axis_iarg_28_tkeep),
        .s_axis_iarg_28_tstrb(s_axis_iarg_28_tstrb),
        .s_axis_iarg_28_tdata(s_axis_iarg_28_tdata),
        .s_axis_iarg_28_tready(s_axis_iarg_28_tready),
        .ap_axis_iarg_28_tlast(ap_axis_iarg_28_tlast),
        .ap_axis_iarg_28_tvalid(ap_axis_iarg_28_tvalid),
        .ap_axis_iarg_28_tkeep(ap_axis_iarg_28_tkeep),
        .ap_axis_iarg_28_tstrb(ap_axis_iarg_28_tstrb),
        .ap_axis_iarg_28_tdata(ap_axis_iarg_28_tdata),
        .ap_axis_iarg_28_tready(ap_axis_iarg_28_tready),
        .s_axis_iarg_29_aclk(s_axis_iarg_29_aclk),
        .s_axis_iarg_29_aresetn(s_axis_iarg_29_aresetn),
        .s_axis_iarg_29_tlast(s_axis_iarg_29_tlast),
        .s_axis_iarg_29_tvalid(s_axis_iarg_29_tvalid),
        .s_axis_iarg_29_tkeep(s_axis_iarg_29_tkeep),
        .s_axis_iarg_29_tstrb(s_axis_iarg_29_tstrb),
        .s_axis_iarg_29_tdata(s_axis_iarg_29_tdata),
        .s_axis_iarg_29_tready(s_axis_iarg_29_tready),
        .ap_axis_iarg_29_tlast(ap_axis_iarg_29_tlast),
        .ap_axis_iarg_29_tvalid(ap_axis_iarg_29_tvalid),
        .ap_axis_iarg_29_tkeep(ap_axis_iarg_29_tkeep),
        .ap_axis_iarg_29_tstrb(ap_axis_iarg_29_tstrb),
        .ap_axis_iarg_29_tdata(ap_axis_iarg_29_tdata),
        .ap_axis_iarg_29_tready(ap_axis_iarg_29_tready),
        .s_axis_iarg_30_aclk(s_axis_iarg_30_aclk),
        .s_axis_iarg_30_aresetn(s_axis_iarg_30_aresetn),
        .s_axis_iarg_30_tlast(s_axis_iarg_30_tlast),
        .s_axis_iarg_30_tvalid(s_axis_iarg_30_tvalid),
        .s_axis_iarg_30_tkeep(s_axis_iarg_30_tkeep),
        .s_axis_iarg_30_tstrb(s_axis_iarg_30_tstrb),
        .s_axis_iarg_30_tdata(s_axis_iarg_30_tdata),
        .s_axis_iarg_30_tready(s_axis_iarg_30_tready),
        .ap_axis_iarg_30_tlast(ap_axis_iarg_30_tlast),
        .ap_axis_iarg_30_tvalid(ap_axis_iarg_30_tvalid),
        .ap_axis_iarg_30_tkeep(ap_axis_iarg_30_tkeep),
        .ap_axis_iarg_30_tstrb(ap_axis_iarg_30_tstrb),
        .ap_axis_iarg_30_tdata(ap_axis_iarg_30_tdata),
        .ap_axis_iarg_30_tready(ap_axis_iarg_30_tready),
        .s_axis_iarg_31_aclk(s_axis_iarg_31_aclk),
        .s_axis_iarg_31_aresetn(s_axis_iarg_31_aresetn),
        .s_axis_iarg_31_tlast(s_axis_iarg_31_tlast),
        .s_axis_iarg_31_tvalid(s_axis_iarg_31_tvalid),
        .s_axis_iarg_31_tkeep(s_axis_iarg_31_tkeep),
        .s_axis_iarg_31_tstrb(s_axis_iarg_31_tstrb),
        .s_axis_iarg_31_tdata(s_axis_iarg_31_tdata),
        .s_axis_iarg_31_tready(s_axis_iarg_31_tready),
        .ap_axis_iarg_31_tlast(ap_axis_iarg_31_tlast),
        .ap_axis_iarg_31_tvalid(ap_axis_iarg_31_tvalid),
        .ap_axis_iarg_31_tkeep(ap_axis_iarg_31_tkeep),
        .ap_axis_iarg_31_tstrb(ap_axis_iarg_31_tstrb),
        .ap_axis_iarg_31_tdata(ap_axis_iarg_31_tdata),
        .ap_axis_iarg_31_tready(ap_axis_iarg_31_tready),
        .s_axis_iarg_32_aclk(s_axis_iarg_32_aclk),
        .s_axis_iarg_32_aresetn(s_axis_iarg_32_aresetn),
        .s_axis_iarg_32_tlast(s_axis_iarg_32_tlast),
        .s_axis_iarg_32_tvalid(s_axis_iarg_32_tvalid),
        .s_axis_iarg_32_tkeep(s_axis_iarg_32_tkeep),
        .s_axis_iarg_32_tstrb(s_axis_iarg_32_tstrb),
        .s_axis_iarg_32_tdata(s_axis_iarg_32_tdata),
        .s_axis_iarg_32_tready(s_axis_iarg_32_tready),
        .ap_axis_iarg_32_tlast(ap_axis_iarg_32_tlast),
        .ap_axis_iarg_32_tvalid(ap_axis_iarg_32_tvalid),
        .ap_axis_iarg_32_tkeep(ap_axis_iarg_32_tkeep),
        .ap_axis_iarg_32_tstrb(ap_axis_iarg_32_tstrb),
        .ap_axis_iarg_32_tdata(ap_axis_iarg_32_tdata),
        .ap_axis_iarg_32_tready(ap_axis_iarg_32_tready),
        .s_axis_iarg_33_aclk(s_axis_iarg_33_aclk),
        .s_axis_iarg_33_aresetn(s_axis_iarg_33_aresetn),
        .s_axis_iarg_33_tlast(s_axis_iarg_33_tlast),
        .s_axis_iarg_33_tvalid(s_axis_iarg_33_tvalid),
        .s_axis_iarg_33_tkeep(s_axis_iarg_33_tkeep),
        .s_axis_iarg_33_tstrb(s_axis_iarg_33_tstrb),
        .s_axis_iarg_33_tdata(s_axis_iarg_33_tdata),
        .s_axis_iarg_33_tready(s_axis_iarg_33_tready),
        .ap_axis_iarg_33_tlast(ap_axis_iarg_33_tlast),
        .ap_axis_iarg_33_tvalid(ap_axis_iarg_33_tvalid),
        .ap_axis_iarg_33_tkeep(ap_axis_iarg_33_tkeep),
        .ap_axis_iarg_33_tstrb(ap_axis_iarg_33_tstrb),
        .ap_axis_iarg_33_tdata(ap_axis_iarg_33_tdata),
        .ap_axis_iarg_33_tready(ap_axis_iarg_33_tready),
        .s_axis_iarg_34_aclk(s_axis_iarg_34_aclk),
        .s_axis_iarg_34_aresetn(s_axis_iarg_34_aresetn),
        .s_axis_iarg_34_tlast(s_axis_iarg_34_tlast),
        .s_axis_iarg_34_tvalid(s_axis_iarg_34_tvalid),
        .s_axis_iarg_34_tkeep(s_axis_iarg_34_tkeep),
        .s_axis_iarg_34_tstrb(s_axis_iarg_34_tstrb),
        .s_axis_iarg_34_tdata(s_axis_iarg_34_tdata),
        .s_axis_iarg_34_tready(s_axis_iarg_34_tready),
        .ap_axis_iarg_34_tlast(ap_axis_iarg_34_tlast),
        .ap_axis_iarg_34_tvalid(ap_axis_iarg_34_tvalid),
        .ap_axis_iarg_34_tkeep(ap_axis_iarg_34_tkeep),
        .ap_axis_iarg_34_tstrb(ap_axis_iarg_34_tstrb),
        .ap_axis_iarg_34_tdata(ap_axis_iarg_34_tdata),
        .ap_axis_iarg_34_tready(ap_axis_iarg_34_tready),
        .s_axis_iarg_35_aclk(s_axis_iarg_35_aclk),
        .s_axis_iarg_35_aresetn(s_axis_iarg_35_aresetn),
        .s_axis_iarg_35_tlast(s_axis_iarg_35_tlast),
        .s_axis_iarg_35_tvalid(s_axis_iarg_35_tvalid),
        .s_axis_iarg_35_tkeep(s_axis_iarg_35_tkeep),
        .s_axis_iarg_35_tstrb(s_axis_iarg_35_tstrb),
        .s_axis_iarg_35_tdata(s_axis_iarg_35_tdata),
        .s_axis_iarg_35_tready(s_axis_iarg_35_tready),
        .ap_axis_iarg_35_tlast(ap_axis_iarg_35_tlast),
        .ap_axis_iarg_35_tvalid(ap_axis_iarg_35_tvalid),
        .ap_axis_iarg_35_tkeep(ap_axis_iarg_35_tkeep),
        .ap_axis_iarg_35_tstrb(ap_axis_iarg_35_tstrb),
        .ap_axis_iarg_35_tdata(ap_axis_iarg_35_tdata),
        .ap_axis_iarg_35_tready(ap_axis_iarg_35_tready),
        .s_axis_iarg_36_aclk(s_axis_iarg_36_aclk),
        .s_axis_iarg_36_aresetn(s_axis_iarg_36_aresetn),
        .s_axis_iarg_36_tlast(s_axis_iarg_36_tlast),
        .s_axis_iarg_36_tvalid(s_axis_iarg_36_tvalid),
        .s_axis_iarg_36_tkeep(s_axis_iarg_36_tkeep),
        .s_axis_iarg_36_tstrb(s_axis_iarg_36_tstrb),
        .s_axis_iarg_36_tdata(s_axis_iarg_36_tdata),
        .s_axis_iarg_36_tready(s_axis_iarg_36_tready),
        .ap_axis_iarg_36_tlast(ap_axis_iarg_36_tlast),
        .ap_axis_iarg_36_tvalid(ap_axis_iarg_36_tvalid),
        .ap_axis_iarg_36_tkeep(ap_axis_iarg_36_tkeep),
        .ap_axis_iarg_36_tstrb(ap_axis_iarg_36_tstrb),
        .ap_axis_iarg_36_tdata(ap_axis_iarg_36_tdata),
        .ap_axis_iarg_36_tready(ap_axis_iarg_36_tready),
        .s_axis_iarg_37_aclk(s_axis_iarg_37_aclk),
        .s_axis_iarg_37_aresetn(s_axis_iarg_37_aresetn),
        .s_axis_iarg_37_tlast(s_axis_iarg_37_tlast),
        .s_axis_iarg_37_tvalid(s_axis_iarg_37_tvalid),
        .s_axis_iarg_37_tkeep(s_axis_iarg_37_tkeep),
        .s_axis_iarg_37_tstrb(s_axis_iarg_37_tstrb),
        .s_axis_iarg_37_tdata(s_axis_iarg_37_tdata),
        .s_axis_iarg_37_tready(s_axis_iarg_37_tready),
        .ap_axis_iarg_37_tlast(ap_axis_iarg_37_tlast),
        .ap_axis_iarg_37_tvalid(ap_axis_iarg_37_tvalid),
        .ap_axis_iarg_37_tkeep(ap_axis_iarg_37_tkeep),
        .ap_axis_iarg_37_tstrb(ap_axis_iarg_37_tstrb),
        .ap_axis_iarg_37_tdata(ap_axis_iarg_37_tdata),
        .ap_axis_iarg_37_tready(ap_axis_iarg_37_tready),
        .s_axis_iarg_38_aclk(s_axis_iarg_38_aclk),
        .s_axis_iarg_38_aresetn(s_axis_iarg_38_aresetn),
        .s_axis_iarg_38_tlast(s_axis_iarg_38_tlast),
        .s_axis_iarg_38_tvalid(s_axis_iarg_38_tvalid),
        .s_axis_iarg_38_tkeep(s_axis_iarg_38_tkeep),
        .s_axis_iarg_38_tstrb(s_axis_iarg_38_tstrb),
        .s_axis_iarg_38_tdata(s_axis_iarg_38_tdata),
        .s_axis_iarg_38_tready(s_axis_iarg_38_tready),
        .ap_axis_iarg_38_tlast(ap_axis_iarg_38_tlast),
        .ap_axis_iarg_38_tvalid(ap_axis_iarg_38_tvalid),
        .ap_axis_iarg_38_tkeep(ap_axis_iarg_38_tkeep),
        .ap_axis_iarg_38_tstrb(ap_axis_iarg_38_tstrb),
        .ap_axis_iarg_38_tdata(ap_axis_iarg_38_tdata),
        .ap_axis_iarg_38_tready(ap_axis_iarg_38_tready),
        .s_axis_iarg_39_aclk(s_axis_iarg_39_aclk),
        .s_axis_iarg_39_aresetn(s_axis_iarg_39_aresetn),
        .s_axis_iarg_39_tlast(s_axis_iarg_39_tlast),
        .s_axis_iarg_39_tvalid(s_axis_iarg_39_tvalid),
        .s_axis_iarg_39_tkeep(s_axis_iarg_39_tkeep),
        .s_axis_iarg_39_tstrb(s_axis_iarg_39_tstrb),
        .s_axis_iarg_39_tdata(s_axis_iarg_39_tdata),
        .s_axis_iarg_39_tready(s_axis_iarg_39_tready),
        .ap_axis_iarg_39_tlast(ap_axis_iarg_39_tlast),
        .ap_axis_iarg_39_tvalid(ap_axis_iarg_39_tvalid),
        .ap_axis_iarg_39_tkeep(ap_axis_iarg_39_tkeep),
        .ap_axis_iarg_39_tstrb(ap_axis_iarg_39_tstrb),
        .ap_axis_iarg_39_tdata(ap_axis_iarg_39_tdata),
        .ap_axis_iarg_39_tready(ap_axis_iarg_39_tready),
        .s_axis_iarg_40_aclk(s_axis_iarg_40_aclk),
        .s_axis_iarg_40_aresetn(s_axis_iarg_40_aresetn),
        .s_axis_iarg_40_tlast(s_axis_iarg_40_tlast),
        .s_axis_iarg_40_tvalid(s_axis_iarg_40_tvalid),
        .s_axis_iarg_40_tkeep(s_axis_iarg_40_tkeep),
        .s_axis_iarg_40_tstrb(s_axis_iarg_40_tstrb),
        .s_axis_iarg_40_tdata(s_axis_iarg_40_tdata),
        .s_axis_iarg_40_tready(s_axis_iarg_40_tready),
        .ap_axis_iarg_40_tlast(ap_axis_iarg_40_tlast),
        .ap_axis_iarg_40_tvalid(ap_axis_iarg_40_tvalid),
        .ap_axis_iarg_40_tkeep(ap_axis_iarg_40_tkeep),
        .ap_axis_iarg_40_tstrb(ap_axis_iarg_40_tstrb),
        .ap_axis_iarg_40_tdata(ap_axis_iarg_40_tdata),
        .ap_axis_iarg_40_tready(ap_axis_iarg_40_tready),
        .s_axis_iarg_41_aclk(s_axis_iarg_41_aclk),
        .s_axis_iarg_41_aresetn(s_axis_iarg_41_aresetn),
        .s_axis_iarg_41_tlast(s_axis_iarg_41_tlast),
        .s_axis_iarg_41_tvalid(s_axis_iarg_41_tvalid),
        .s_axis_iarg_41_tkeep(s_axis_iarg_41_tkeep),
        .s_axis_iarg_41_tstrb(s_axis_iarg_41_tstrb),
        .s_axis_iarg_41_tdata(s_axis_iarg_41_tdata),
        .s_axis_iarg_41_tready(s_axis_iarg_41_tready),
        .ap_axis_iarg_41_tlast(ap_axis_iarg_41_tlast),
        .ap_axis_iarg_41_tvalid(ap_axis_iarg_41_tvalid),
        .ap_axis_iarg_41_tkeep(ap_axis_iarg_41_tkeep),
        .ap_axis_iarg_41_tstrb(ap_axis_iarg_41_tstrb),
        .ap_axis_iarg_41_tdata(ap_axis_iarg_41_tdata),
        .ap_axis_iarg_41_tready(ap_axis_iarg_41_tready),
        .s_axis_iarg_42_aclk(s_axis_iarg_42_aclk),
        .s_axis_iarg_42_aresetn(s_axis_iarg_42_aresetn),
        .s_axis_iarg_42_tlast(s_axis_iarg_42_tlast),
        .s_axis_iarg_42_tvalid(s_axis_iarg_42_tvalid),
        .s_axis_iarg_42_tkeep(s_axis_iarg_42_tkeep),
        .s_axis_iarg_42_tstrb(s_axis_iarg_42_tstrb),
        .s_axis_iarg_42_tdata(s_axis_iarg_42_tdata),
        .s_axis_iarg_42_tready(s_axis_iarg_42_tready),
        .ap_axis_iarg_42_tlast(ap_axis_iarg_42_tlast),
        .ap_axis_iarg_42_tvalid(ap_axis_iarg_42_tvalid),
        .ap_axis_iarg_42_tkeep(ap_axis_iarg_42_tkeep),
        .ap_axis_iarg_42_tstrb(ap_axis_iarg_42_tstrb),
        .ap_axis_iarg_42_tdata(ap_axis_iarg_42_tdata),
        .ap_axis_iarg_42_tready(ap_axis_iarg_42_tready),
        .s_axis_iarg_43_aclk(s_axis_iarg_43_aclk),
        .s_axis_iarg_43_aresetn(s_axis_iarg_43_aresetn),
        .s_axis_iarg_43_tlast(s_axis_iarg_43_tlast),
        .s_axis_iarg_43_tvalid(s_axis_iarg_43_tvalid),
        .s_axis_iarg_43_tkeep(s_axis_iarg_43_tkeep),
        .s_axis_iarg_43_tstrb(s_axis_iarg_43_tstrb),
        .s_axis_iarg_43_tdata(s_axis_iarg_43_tdata),
        .s_axis_iarg_43_tready(s_axis_iarg_43_tready),
        .ap_axis_iarg_43_tlast(ap_axis_iarg_43_tlast),
        .ap_axis_iarg_43_tvalid(ap_axis_iarg_43_tvalid),
        .ap_axis_iarg_43_tkeep(ap_axis_iarg_43_tkeep),
        .ap_axis_iarg_43_tstrb(ap_axis_iarg_43_tstrb),
        .ap_axis_iarg_43_tdata(ap_axis_iarg_43_tdata),
        .ap_axis_iarg_43_tready(ap_axis_iarg_43_tready),
        .s_axis_iarg_44_aclk(s_axis_iarg_44_aclk),
        .s_axis_iarg_44_aresetn(s_axis_iarg_44_aresetn),
        .s_axis_iarg_44_tlast(s_axis_iarg_44_tlast),
        .s_axis_iarg_44_tvalid(s_axis_iarg_44_tvalid),
        .s_axis_iarg_44_tkeep(s_axis_iarg_44_tkeep),
        .s_axis_iarg_44_tstrb(s_axis_iarg_44_tstrb),
        .s_axis_iarg_44_tdata(s_axis_iarg_44_tdata),
        .s_axis_iarg_44_tready(s_axis_iarg_44_tready),
        .ap_axis_iarg_44_tlast(ap_axis_iarg_44_tlast),
        .ap_axis_iarg_44_tvalid(ap_axis_iarg_44_tvalid),
        .ap_axis_iarg_44_tkeep(ap_axis_iarg_44_tkeep),
        .ap_axis_iarg_44_tstrb(ap_axis_iarg_44_tstrb),
        .ap_axis_iarg_44_tdata(ap_axis_iarg_44_tdata),
        .ap_axis_iarg_44_tready(ap_axis_iarg_44_tready),
        .s_axis_iarg_45_aclk(s_axis_iarg_45_aclk),
        .s_axis_iarg_45_aresetn(s_axis_iarg_45_aresetn),
        .s_axis_iarg_45_tlast(s_axis_iarg_45_tlast),
        .s_axis_iarg_45_tvalid(s_axis_iarg_45_tvalid),
        .s_axis_iarg_45_tkeep(s_axis_iarg_45_tkeep),
        .s_axis_iarg_45_tstrb(s_axis_iarg_45_tstrb),
        .s_axis_iarg_45_tdata(s_axis_iarg_45_tdata),
        .s_axis_iarg_45_tready(s_axis_iarg_45_tready),
        .ap_axis_iarg_45_tlast(ap_axis_iarg_45_tlast),
        .ap_axis_iarg_45_tvalid(ap_axis_iarg_45_tvalid),
        .ap_axis_iarg_45_tkeep(ap_axis_iarg_45_tkeep),
        .ap_axis_iarg_45_tstrb(ap_axis_iarg_45_tstrb),
        .ap_axis_iarg_45_tdata(ap_axis_iarg_45_tdata),
        .ap_axis_iarg_45_tready(ap_axis_iarg_45_tready),
        .s_axis_iarg_46_aclk(s_axis_iarg_46_aclk),
        .s_axis_iarg_46_aresetn(s_axis_iarg_46_aresetn),
        .s_axis_iarg_46_tlast(s_axis_iarg_46_tlast),
        .s_axis_iarg_46_tvalid(s_axis_iarg_46_tvalid),
        .s_axis_iarg_46_tkeep(s_axis_iarg_46_tkeep),
        .s_axis_iarg_46_tstrb(s_axis_iarg_46_tstrb),
        .s_axis_iarg_46_tdata(s_axis_iarg_46_tdata),
        .s_axis_iarg_46_tready(s_axis_iarg_46_tready),
        .ap_axis_iarg_46_tlast(ap_axis_iarg_46_tlast),
        .ap_axis_iarg_46_tvalid(ap_axis_iarg_46_tvalid),
        .ap_axis_iarg_46_tkeep(ap_axis_iarg_46_tkeep),
        .ap_axis_iarg_46_tstrb(ap_axis_iarg_46_tstrb),
        .ap_axis_iarg_46_tdata(ap_axis_iarg_46_tdata),
        .ap_axis_iarg_46_tready(ap_axis_iarg_46_tready),
        .s_axis_iarg_47_aclk(s_axis_iarg_47_aclk),
        .s_axis_iarg_47_aresetn(s_axis_iarg_47_aresetn),
        .s_axis_iarg_47_tlast(s_axis_iarg_47_tlast),
        .s_axis_iarg_47_tvalid(s_axis_iarg_47_tvalid),
        .s_axis_iarg_47_tkeep(s_axis_iarg_47_tkeep),
        .s_axis_iarg_47_tstrb(s_axis_iarg_47_tstrb),
        .s_axis_iarg_47_tdata(s_axis_iarg_47_tdata),
        .s_axis_iarg_47_tready(s_axis_iarg_47_tready),
        .ap_axis_iarg_47_tlast(ap_axis_iarg_47_tlast),
        .ap_axis_iarg_47_tvalid(ap_axis_iarg_47_tvalid),
        .ap_axis_iarg_47_tkeep(ap_axis_iarg_47_tkeep),
        .ap_axis_iarg_47_tstrb(ap_axis_iarg_47_tstrb),
        .ap_axis_iarg_47_tdata(ap_axis_iarg_47_tdata),
        .ap_axis_iarg_47_tready(ap_axis_iarg_47_tready),
        .s_axis_iarg_48_aclk(s_axis_iarg_48_aclk),
        .s_axis_iarg_48_aresetn(s_axis_iarg_48_aresetn),
        .s_axis_iarg_48_tlast(s_axis_iarg_48_tlast),
        .s_axis_iarg_48_tvalid(s_axis_iarg_48_tvalid),
        .s_axis_iarg_48_tkeep(s_axis_iarg_48_tkeep),
        .s_axis_iarg_48_tstrb(s_axis_iarg_48_tstrb),
        .s_axis_iarg_48_tdata(s_axis_iarg_48_tdata),
        .s_axis_iarg_48_tready(s_axis_iarg_48_tready),
        .ap_axis_iarg_48_tlast(ap_axis_iarg_48_tlast),
        .ap_axis_iarg_48_tvalid(ap_axis_iarg_48_tvalid),
        .ap_axis_iarg_48_tkeep(ap_axis_iarg_48_tkeep),
        .ap_axis_iarg_48_tstrb(ap_axis_iarg_48_tstrb),
        .ap_axis_iarg_48_tdata(ap_axis_iarg_48_tdata),
        .ap_axis_iarg_48_tready(ap_axis_iarg_48_tready),
        .s_axis_iarg_49_aclk(s_axis_iarg_49_aclk),
        .s_axis_iarg_49_aresetn(s_axis_iarg_49_aresetn),
        .s_axis_iarg_49_tlast(s_axis_iarg_49_tlast),
        .s_axis_iarg_49_tvalid(s_axis_iarg_49_tvalid),
        .s_axis_iarg_49_tkeep(s_axis_iarg_49_tkeep),
        .s_axis_iarg_49_tstrb(s_axis_iarg_49_tstrb),
        .s_axis_iarg_49_tdata(s_axis_iarg_49_tdata),
        .s_axis_iarg_49_tready(s_axis_iarg_49_tready),
        .ap_axis_iarg_49_tlast(ap_axis_iarg_49_tlast),
        .ap_axis_iarg_49_tvalid(ap_axis_iarg_49_tvalid),
        .ap_axis_iarg_49_tkeep(ap_axis_iarg_49_tkeep),
        .ap_axis_iarg_49_tstrb(ap_axis_iarg_49_tstrb),
        .ap_axis_iarg_49_tdata(ap_axis_iarg_49_tdata),
        .ap_axis_iarg_49_tready(ap_axis_iarg_49_tready),
        .s_axis_iarg_50_aclk(s_axis_iarg_50_aclk),
        .s_axis_iarg_50_aresetn(s_axis_iarg_50_aresetn),
        .s_axis_iarg_50_tlast(s_axis_iarg_50_tlast),
        .s_axis_iarg_50_tvalid(s_axis_iarg_50_tvalid),
        .s_axis_iarg_50_tkeep(s_axis_iarg_50_tkeep),
        .s_axis_iarg_50_tstrb(s_axis_iarg_50_tstrb),
        .s_axis_iarg_50_tdata(s_axis_iarg_50_tdata),
        .s_axis_iarg_50_tready(s_axis_iarg_50_tready),
        .ap_axis_iarg_50_tlast(ap_axis_iarg_50_tlast),
        .ap_axis_iarg_50_tvalid(ap_axis_iarg_50_tvalid),
        .ap_axis_iarg_50_tkeep(ap_axis_iarg_50_tkeep),
        .ap_axis_iarg_50_tstrb(ap_axis_iarg_50_tstrb),
        .ap_axis_iarg_50_tdata(ap_axis_iarg_50_tdata),
        .ap_axis_iarg_50_tready(ap_axis_iarg_50_tready),
        .s_axis_iarg_51_aclk(s_axis_iarg_51_aclk),
        .s_axis_iarg_51_aresetn(s_axis_iarg_51_aresetn),
        .s_axis_iarg_51_tlast(s_axis_iarg_51_tlast),
        .s_axis_iarg_51_tvalid(s_axis_iarg_51_tvalid),
        .s_axis_iarg_51_tkeep(s_axis_iarg_51_tkeep),
        .s_axis_iarg_51_tstrb(s_axis_iarg_51_tstrb),
        .s_axis_iarg_51_tdata(s_axis_iarg_51_tdata),
        .s_axis_iarg_51_tready(s_axis_iarg_51_tready),
        .ap_axis_iarg_51_tlast(ap_axis_iarg_51_tlast),
        .ap_axis_iarg_51_tvalid(ap_axis_iarg_51_tvalid),
        .ap_axis_iarg_51_tkeep(ap_axis_iarg_51_tkeep),
        .ap_axis_iarg_51_tstrb(ap_axis_iarg_51_tstrb),
        .ap_axis_iarg_51_tdata(ap_axis_iarg_51_tdata),
        .ap_axis_iarg_51_tready(ap_axis_iarg_51_tready),
        .s_axis_iarg_52_aclk(s_axis_iarg_52_aclk),
        .s_axis_iarg_52_aresetn(s_axis_iarg_52_aresetn),
        .s_axis_iarg_52_tlast(s_axis_iarg_52_tlast),
        .s_axis_iarg_52_tvalid(s_axis_iarg_52_tvalid),
        .s_axis_iarg_52_tkeep(s_axis_iarg_52_tkeep),
        .s_axis_iarg_52_tstrb(s_axis_iarg_52_tstrb),
        .s_axis_iarg_52_tdata(s_axis_iarg_52_tdata),
        .s_axis_iarg_52_tready(s_axis_iarg_52_tready),
        .ap_axis_iarg_52_tlast(ap_axis_iarg_52_tlast),
        .ap_axis_iarg_52_tvalid(ap_axis_iarg_52_tvalid),
        .ap_axis_iarg_52_tkeep(ap_axis_iarg_52_tkeep),
        .ap_axis_iarg_52_tstrb(ap_axis_iarg_52_tstrb),
        .ap_axis_iarg_52_tdata(ap_axis_iarg_52_tdata),
        .ap_axis_iarg_52_tready(ap_axis_iarg_52_tready),
        .s_axis_iarg_53_aclk(s_axis_iarg_53_aclk),
        .s_axis_iarg_53_aresetn(s_axis_iarg_53_aresetn),
        .s_axis_iarg_53_tlast(s_axis_iarg_53_tlast),
        .s_axis_iarg_53_tvalid(s_axis_iarg_53_tvalid),
        .s_axis_iarg_53_tkeep(s_axis_iarg_53_tkeep),
        .s_axis_iarg_53_tstrb(s_axis_iarg_53_tstrb),
        .s_axis_iarg_53_tdata(s_axis_iarg_53_tdata),
        .s_axis_iarg_53_tready(s_axis_iarg_53_tready),
        .ap_axis_iarg_53_tlast(ap_axis_iarg_53_tlast),
        .ap_axis_iarg_53_tvalid(ap_axis_iarg_53_tvalid),
        .ap_axis_iarg_53_tkeep(ap_axis_iarg_53_tkeep),
        .ap_axis_iarg_53_tstrb(ap_axis_iarg_53_tstrb),
        .ap_axis_iarg_53_tdata(ap_axis_iarg_53_tdata),
        .ap_axis_iarg_53_tready(ap_axis_iarg_53_tready),
        .s_axis_iarg_54_aclk(s_axis_iarg_54_aclk),
        .s_axis_iarg_54_aresetn(s_axis_iarg_54_aresetn),
        .s_axis_iarg_54_tlast(s_axis_iarg_54_tlast),
        .s_axis_iarg_54_tvalid(s_axis_iarg_54_tvalid),
        .s_axis_iarg_54_tkeep(s_axis_iarg_54_tkeep),
        .s_axis_iarg_54_tstrb(s_axis_iarg_54_tstrb),
        .s_axis_iarg_54_tdata(s_axis_iarg_54_tdata),
        .s_axis_iarg_54_tready(s_axis_iarg_54_tready),
        .ap_axis_iarg_54_tlast(ap_axis_iarg_54_tlast),
        .ap_axis_iarg_54_tvalid(ap_axis_iarg_54_tvalid),
        .ap_axis_iarg_54_tkeep(ap_axis_iarg_54_tkeep),
        .ap_axis_iarg_54_tstrb(ap_axis_iarg_54_tstrb),
        .ap_axis_iarg_54_tdata(ap_axis_iarg_54_tdata),
        .ap_axis_iarg_54_tready(ap_axis_iarg_54_tready),
        .s_axis_iarg_55_aclk(s_axis_iarg_55_aclk),
        .s_axis_iarg_55_aresetn(s_axis_iarg_55_aresetn),
        .s_axis_iarg_55_tlast(s_axis_iarg_55_tlast),
        .s_axis_iarg_55_tvalid(s_axis_iarg_55_tvalid),
        .s_axis_iarg_55_tkeep(s_axis_iarg_55_tkeep),
        .s_axis_iarg_55_tstrb(s_axis_iarg_55_tstrb),
        .s_axis_iarg_55_tdata(s_axis_iarg_55_tdata),
        .s_axis_iarg_55_tready(s_axis_iarg_55_tready),
        .ap_axis_iarg_55_tlast(ap_axis_iarg_55_tlast),
        .ap_axis_iarg_55_tvalid(ap_axis_iarg_55_tvalid),
        .ap_axis_iarg_55_tkeep(ap_axis_iarg_55_tkeep),
        .ap_axis_iarg_55_tstrb(ap_axis_iarg_55_tstrb),
        .ap_axis_iarg_55_tdata(ap_axis_iarg_55_tdata),
        .ap_axis_iarg_55_tready(ap_axis_iarg_55_tready),
        .s_axis_iarg_56_aclk(s_axis_iarg_56_aclk),
        .s_axis_iarg_56_aresetn(s_axis_iarg_56_aresetn),
        .s_axis_iarg_56_tlast(s_axis_iarg_56_tlast),
        .s_axis_iarg_56_tvalid(s_axis_iarg_56_tvalid),
        .s_axis_iarg_56_tkeep(s_axis_iarg_56_tkeep),
        .s_axis_iarg_56_tstrb(s_axis_iarg_56_tstrb),
        .s_axis_iarg_56_tdata(s_axis_iarg_56_tdata),
        .s_axis_iarg_56_tready(s_axis_iarg_56_tready),
        .ap_axis_iarg_56_tlast(ap_axis_iarg_56_tlast),
        .ap_axis_iarg_56_tvalid(ap_axis_iarg_56_tvalid),
        .ap_axis_iarg_56_tkeep(ap_axis_iarg_56_tkeep),
        .ap_axis_iarg_56_tstrb(ap_axis_iarg_56_tstrb),
        .ap_axis_iarg_56_tdata(ap_axis_iarg_56_tdata),
        .ap_axis_iarg_56_tready(ap_axis_iarg_56_tready),
        .s_axis_iarg_57_aclk(s_axis_iarg_57_aclk),
        .s_axis_iarg_57_aresetn(s_axis_iarg_57_aresetn),
        .s_axis_iarg_57_tlast(s_axis_iarg_57_tlast),
        .s_axis_iarg_57_tvalid(s_axis_iarg_57_tvalid),
        .s_axis_iarg_57_tkeep(s_axis_iarg_57_tkeep),
        .s_axis_iarg_57_tstrb(s_axis_iarg_57_tstrb),
        .s_axis_iarg_57_tdata(s_axis_iarg_57_tdata),
        .s_axis_iarg_57_tready(s_axis_iarg_57_tready),
        .ap_axis_iarg_57_tlast(ap_axis_iarg_57_tlast),
        .ap_axis_iarg_57_tvalid(ap_axis_iarg_57_tvalid),
        .ap_axis_iarg_57_tkeep(ap_axis_iarg_57_tkeep),
        .ap_axis_iarg_57_tstrb(ap_axis_iarg_57_tstrb),
        .ap_axis_iarg_57_tdata(ap_axis_iarg_57_tdata),
        .ap_axis_iarg_57_tready(ap_axis_iarg_57_tready),
        .s_axis_iarg_58_aclk(s_axis_iarg_58_aclk),
        .s_axis_iarg_58_aresetn(s_axis_iarg_58_aresetn),
        .s_axis_iarg_58_tlast(s_axis_iarg_58_tlast),
        .s_axis_iarg_58_tvalid(s_axis_iarg_58_tvalid),
        .s_axis_iarg_58_tkeep(s_axis_iarg_58_tkeep),
        .s_axis_iarg_58_tstrb(s_axis_iarg_58_tstrb),
        .s_axis_iarg_58_tdata(s_axis_iarg_58_tdata),
        .s_axis_iarg_58_tready(s_axis_iarg_58_tready),
        .ap_axis_iarg_58_tlast(ap_axis_iarg_58_tlast),
        .ap_axis_iarg_58_tvalid(ap_axis_iarg_58_tvalid),
        .ap_axis_iarg_58_tkeep(ap_axis_iarg_58_tkeep),
        .ap_axis_iarg_58_tstrb(ap_axis_iarg_58_tstrb),
        .ap_axis_iarg_58_tdata(ap_axis_iarg_58_tdata),
        .ap_axis_iarg_58_tready(ap_axis_iarg_58_tready),
        .s_axis_iarg_59_aclk(s_axis_iarg_59_aclk),
        .s_axis_iarg_59_aresetn(s_axis_iarg_59_aresetn),
        .s_axis_iarg_59_tlast(s_axis_iarg_59_tlast),
        .s_axis_iarg_59_tvalid(s_axis_iarg_59_tvalid),
        .s_axis_iarg_59_tkeep(s_axis_iarg_59_tkeep),
        .s_axis_iarg_59_tstrb(s_axis_iarg_59_tstrb),
        .s_axis_iarg_59_tdata(s_axis_iarg_59_tdata),
        .s_axis_iarg_59_tready(s_axis_iarg_59_tready),
        .ap_axis_iarg_59_tlast(ap_axis_iarg_59_tlast),
        .ap_axis_iarg_59_tvalid(ap_axis_iarg_59_tvalid),
        .ap_axis_iarg_59_tkeep(ap_axis_iarg_59_tkeep),
        .ap_axis_iarg_59_tstrb(ap_axis_iarg_59_tstrb),
        .ap_axis_iarg_59_tdata(ap_axis_iarg_59_tdata),
        .ap_axis_iarg_59_tready(ap_axis_iarg_59_tready),
        .s_axis_iarg_60_aclk(s_axis_iarg_60_aclk),
        .s_axis_iarg_60_aresetn(s_axis_iarg_60_aresetn),
        .s_axis_iarg_60_tlast(s_axis_iarg_60_tlast),
        .s_axis_iarg_60_tvalid(s_axis_iarg_60_tvalid),
        .s_axis_iarg_60_tkeep(s_axis_iarg_60_tkeep),
        .s_axis_iarg_60_tstrb(s_axis_iarg_60_tstrb),
        .s_axis_iarg_60_tdata(s_axis_iarg_60_tdata),
        .s_axis_iarg_60_tready(s_axis_iarg_60_tready),
        .ap_axis_iarg_60_tlast(ap_axis_iarg_60_tlast),
        .ap_axis_iarg_60_tvalid(ap_axis_iarg_60_tvalid),
        .ap_axis_iarg_60_tkeep(ap_axis_iarg_60_tkeep),
        .ap_axis_iarg_60_tstrb(ap_axis_iarg_60_tstrb),
        .ap_axis_iarg_60_tdata(ap_axis_iarg_60_tdata),
        .ap_axis_iarg_60_tready(ap_axis_iarg_60_tready),
        .s_axis_iarg_61_aclk(s_axis_iarg_61_aclk),
        .s_axis_iarg_61_aresetn(s_axis_iarg_61_aresetn),
        .s_axis_iarg_61_tlast(s_axis_iarg_61_tlast),
        .s_axis_iarg_61_tvalid(s_axis_iarg_61_tvalid),
        .s_axis_iarg_61_tkeep(s_axis_iarg_61_tkeep),
        .s_axis_iarg_61_tstrb(s_axis_iarg_61_tstrb),
        .s_axis_iarg_61_tdata(s_axis_iarg_61_tdata),
        .s_axis_iarg_61_tready(s_axis_iarg_61_tready),
        .ap_axis_iarg_61_tlast(ap_axis_iarg_61_tlast),
        .ap_axis_iarg_61_tvalid(ap_axis_iarg_61_tvalid),
        .ap_axis_iarg_61_tkeep(ap_axis_iarg_61_tkeep),
        .ap_axis_iarg_61_tstrb(ap_axis_iarg_61_tstrb),
        .ap_axis_iarg_61_tdata(ap_axis_iarg_61_tdata),
        .ap_axis_iarg_61_tready(ap_axis_iarg_61_tready),
        .s_axis_iarg_62_aclk(s_axis_iarg_62_aclk),
        .s_axis_iarg_62_aresetn(s_axis_iarg_62_aresetn),
        .s_axis_iarg_62_tlast(s_axis_iarg_62_tlast),
        .s_axis_iarg_62_tvalid(s_axis_iarg_62_tvalid),
        .s_axis_iarg_62_tkeep(s_axis_iarg_62_tkeep),
        .s_axis_iarg_62_tstrb(s_axis_iarg_62_tstrb),
        .s_axis_iarg_62_tdata(s_axis_iarg_62_tdata),
        .s_axis_iarg_62_tready(s_axis_iarg_62_tready),
        .ap_axis_iarg_62_tlast(ap_axis_iarg_62_tlast),
        .ap_axis_iarg_62_tvalid(ap_axis_iarg_62_tvalid),
        .ap_axis_iarg_62_tkeep(ap_axis_iarg_62_tkeep),
        .ap_axis_iarg_62_tstrb(ap_axis_iarg_62_tstrb),
        .ap_axis_iarg_62_tdata(ap_axis_iarg_62_tdata),
        .ap_axis_iarg_62_tready(ap_axis_iarg_62_tready),
        .s_axis_iarg_63_aclk(s_axis_iarg_63_aclk),
        .s_axis_iarg_63_aresetn(s_axis_iarg_63_aresetn),
        .s_axis_iarg_63_tlast(s_axis_iarg_63_tlast),
        .s_axis_iarg_63_tvalid(s_axis_iarg_63_tvalid),
        .s_axis_iarg_63_tkeep(s_axis_iarg_63_tkeep),
        .s_axis_iarg_63_tstrb(s_axis_iarg_63_tstrb),
        .s_axis_iarg_63_tdata(s_axis_iarg_63_tdata),
        .s_axis_iarg_63_tready(s_axis_iarg_63_tready),
        .ap_axis_iarg_63_tlast(ap_axis_iarg_63_tlast),
        .ap_axis_iarg_63_tvalid(ap_axis_iarg_63_tvalid),
        .ap_axis_iarg_63_tkeep(ap_axis_iarg_63_tkeep),
        .ap_axis_iarg_63_tstrb(ap_axis_iarg_63_tstrb),
        .ap_axis_iarg_63_tdata(ap_axis_iarg_63_tdata),
        .ap_axis_iarg_63_tready(ap_axis_iarg_63_tready),
        .s_axis_iarg_64_aclk(s_axis_iarg_64_aclk),
        .s_axis_iarg_64_aresetn(s_axis_iarg_64_aresetn),
        .s_axis_iarg_64_tlast(s_axis_iarg_64_tlast),
        .s_axis_iarg_64_tvalid(s_axis_iarg_64_tvalid),
        .s_axis_iarg_64_tkeep(s_axis_iarg_64_tkeep),
        .s_axis_iarg_64_tstrb(s_axis_iarg_64_tstrb),
        .s_axis_iarg_64_tdata(s_axis_iarg_64_tdata),
        .s_axis_iarg_64_tready(s_axis_iarg_64_tready),
        .ap_axis_iarg_64_tlast(ap_axis_iarg_64_tlast),
        .ap_axis_iarg_64_tvalid(ap_axis_iarg_64_tvalid),
        .ap_axis_iarg_64_tkeep(ap_axis_iarg_64_tkeep),
        .ap_axis_iarg_64_tstrb(ap_axis_iarg_64_tstrb),
        .ap_axis_iarg_64_tdata(ap_axis_iarg_64_tdata),
        .ap_axis_iarg_64_tready(ap_axis_iarg_64_tready),
        .s_axis_iarg_65_aclk(s_axis_iarg_65_aclk),
        .s_axis_iarg_65_aresetn(s_axis_iarg_65_aresetn),
        .s_axis_iarg_65_tlast(s_axis_iarg_65_tlast),
        .s_axis_iarg_65_tvalid(s_axis_iarg_65_tvalid),
        .s_axis_iarg_65_tkeep(s_axis_iarg_65_tkeep),
        .s_axis_iarg_65_tstrb(s_axis_iarg_65_tstrb),
        .s_axis_iarg_65_tdata(s_axis_iarg_65_tdata),
        .s_axis_iarg_65_tready(s_axis_iarg_65_tready),
        .ap_axis_iarg_65_tlast(ap_axis_iarg_65_tlast),
        .ap_axis_iarg_65_tvalid(ap_axis_iarg_65_tvalid),
        .ap_axis_iarg_65_tkeep(ap_axis_iarg_65_tkeep),
        .ap_axis_iarg_65_tstrb(ap_axis_iarg_65_tstrb),
        .ap_axis_iarg_65_tdata(ap_axis_iarg_65_tdata),
        .ap_axis_iarg_65_tready(ap_axis_iarg_65_tready),
        .s_axis_iarg_66_aclk(s_axis_iarg_66_aclk),
        .s_axis_iarg_66_aresetn(s_axis_iarg_66_aresetn),
        .s_axis_iarg_66_tlast(s_axis_iarg_66_tlast),
        .s_axis_iarg_66_tvalid(s_axis_iarg_66_tvalid),
        .s_axis_iarg_66_tkeep(s_axis_iarg_66_tkeep),
        .s_axis_iarg_66_tstrb(s_axis_iarg_66_tstrb),
        .s_axis_iarg_66_tdata(s_axis_iarg_66_tdata),
        .s_axis_iarg_66_tready(s_axis_iarg_66_tready),
        .ap_axis_iarg_66_tlast(ap_axis_iarg_66_tlast),
        .ap_axis_iarg_66_tvalid(ap_axis_iarg_66_tvalid),
        .ap_axis_iarg_66_tkeep(ap_axis_iarg_66_tkeep),
        .ap_axis_iarg_66_tstrb(ap_axis_iarg_66_tstrb),
        .ap_axis_iarg_66_tdata(ap_axis_iarg_66_tdata),
        .ap_axis_iarg_66_tready(ap_axis_iarg_66_tready),
        .s_axis_iarg_67_aclk(s_axis_iarg_67_aclk),
        .s_axis_iarg_67_aresetn(s_axis_iarg_67_aresetn),
        .s_axis_iarg_67_tlast(s_axis_iarg_67_tlast),
        .s_axis_iarg_67_tvalid(s_axis_iarg_67_tvalid),
        .s_axis_iarg_67_tkeep(s_axis_iarg_67_tkeep),
        .s_axis_iarg_67_tstrb(s_axis_iarg_67_tstrb),
        .s_axis_iarg_67_tdata(s_axis_iarg_67_tdata),
        .s_axis_iarg_67_tready(s_axis_iarg_67_tready),
        .ap_axis_iarg_67_tlast(ap_axis_iarg_67_tlast),
        .ap_axis_iarg_67_tvalid(ap_axis_iarg_67_tvalid),
        .ap_axis_iarg_67_tkeep(ap_axis_iarg_67_tkeep),
        .ap_axis_iarg_67_tstrb(ap_axis_iarg_67_tstrb),
        .ap_axis_iarg_67_tdata(ap_axis_iarg_67_tdata),
        .ap_axis_iarg_67_tready(ap_axis_iarg_67_tready),
        .s_axis_iarg_68_aclk(s_axis_iarg_68_aclk),
        .s_axis_iarg_68_aresetn(s_axis_iarg_68_aresetn),
        .s_axis_iarg_68_tlast(s_axis_iarg_68_tlast),
        .s_axis_iarg_68_tvalid(s_axis_iarg_68_tvalid),
        .s_axis_iarg_68_tkeep(s_axis_iarg_68_tkeep),
        .s_axis_iarg_68_tstrb(s_axis_iarg_68_tstrb),
        .s_axis_iarg_68_tdata(s_axis_iarg_68_tdata),
        .s_axis_iarg_68_tready(s_axis_iarg_68_tready),
        .ap_axis_iarg_68_tlast(ap_axis_iarg_68_tlast),
        .ap_axis_iarg_68_tvalid(ap_axis_iarg_68_tvalid),
        .ap_axis_iarg_68_tkeep(ap_axis_iarg_68_tkeep),
        .ap_axis_iarg_68_tstrb(ap_axis_iarg_68_tstrb),
        .ap_axis_iarg_68_tdata(ap_axis_iarg_68_tdata),
        .ap_axis_iarg_68_tready(ap_axis_iarg_68_tready),
        .s_axis_iarg_69_aclk(s_axis_iarg_69_aclk),
        .s_axis_iarg_69_aresetn(s_axis_iarg_69_aresetn),
        .s_axis_iarg_69_tlast(s_axis_iarg_69_tlast),
        .s_axis_iarg_69_tvalid(s_axis_iarg_69_tvalid),
        .s_axis_iarg_69_tkeep(s_axis_iarg_69_tkeep),
        .s_axis_iarg_69_tstrb(s_axis_iarg_69_tstrb),
        .s_axis_iarg_69_tdata(s_axis_iarg_69_tdata),
        .s_axis_iarg_69_tready(s_axis_iarg_69_tready),
        .ap_axis_iarg_69_tlast(ap_axis_iarg_69_tlast),
        .ap_axis_iarg_69_tvalid(ap_axis_iarg_69_tvalid),
        .ap_axis_iarg_69_tkeep(ap_axis_iarg_69_tkeep),
        .ap_axis_iarg_69_tstrb(ap_axis_iarg_69_tstrb),
        .ap_axis_iarg_69_tdata(ap_axis_iarg_69_tdata),
        .ap_axis_iarg_69_tready(ap_axis_iarg_69_tready),
        .s_axis_iarg_70_aclk(s_axis_iarg_70_aclk),
        .s_axis_iarg_70_aresetn(s_axis_iarg_70_aresetn),
        .s_axis_iarg_70_tlast(s_axis_iarg_70_tlast),
        .s_axis_iarg_70_tvalid(s_axis_iarg_70_tvalid),
        .s_axis_iarg_70_tkeep(s_axis_iarg_70_tkeep),
        .s_axis_iarg_70_tstrb(s_axis_iarg_70_tstrb),
        .s_axis_iarg_70_tdata(s_axis_iarg_70_tdata),
        .s_axis_iarg_70_tready(s_axis_iarg_70_tready),
        .ap_axis_iarg_70_tlast(ap_axis_iarg_70_tlast),
        .ap_axis_iarg_70_tvalid(ap_axis_iarg_70_tvalid),
        .ap_axis_iarg_70_tkeep(ap_axis_iarg_70_tkeep),
        .ap_axis_iarg_70_tstrb(ap_axis_iarg_70_tstrb),
        .ap_axis_iarg_70_tdata(ap_axis_iarg_70_tdata),
        .ap_axis_iarg_70_tready(ap_axis_iarg_70_tready),
        .s_axis_iarg_71_aclk(s_axis_iarg_71_aclk),
        .s_axis_iarg_71_aresetn(s_axis_iarg_71_aresetn),
        .s_axis_iarg_71_tlast(s_axis_iarg_71_tlast),
        .s_axis_iarg_71_tvalid(s_axis_iarg_71_tvalid),
        .s_axis_iarg_71_tkeep(s_axis_iarg_71_tkeep),
        .s_axis_iarg_71_tstrb(s_axis_iarg_71_tstrb),
        .s_axis_iarg_71_tdata(s_axis_iarg_71_tdata),
        .s_axis_iarg_71_tready(s_axis_iarg_71_tready),
        .ap_axis_iarg_71_tlast(ap_axis_iarg_71_tlast),
        .ap_axis_iarg_71_tvalid(ap_axis_iarg_71_tvalid),
        .ap_axis_iarg_71_tkeep(ap_axis_iarg_71_tkeep),
        .ap_axis_iarg_71_tstrb(ap_axis_iarg_71_tstrb),
        .ap_axis_iarg_71_tdata(ap_axis_iarg_71_tdata),
        .ap_axis_iarg_71_tready(ap_axis_iarg_71_tready),
        .s_axis_iarg_72_aclk(s_axis_iarg_72_aclk),
        .s_axis_iarg_72_aresetn(s_axis_iarg_72_aresetn),
        .s_axis_iarg_72_tlast(s_axis_iarg_72_tlast),
        .s_axis_iarg_72_tvalid(s_axis_iarg_72_tvalid),
        .s_axis_iarg_72_tkeep(s_axis_iarg_72_tkeep),
        .s_axis_iarg_72_tstrb(s_axis_iarg_72_tstrb),
        .s_axis_iarg_72_tdata(s_axis_iarg_72_tdata),
        .s_axis_iarg_72_tready(s_axis_iarg_72_tready),
        .ap_axis_iarg_72_tlast(ap_axis_iarg_72_tlast),
        .ap_axis_iarg_72_tvalid(ap_axis_iarg_72_tvalid),
        .ap_axis_iarg_72_tkeep(ap_axis_iarg_72_tkeep),
        .ap_axis_iarg_72_tstrb(ap_axis_iarg_72_tstrb),
        .ap_axis_iarg_72_tdata(ap_axis_iarg_72_tdata),
        .ap_axis_iarg_72_tready(ap_axis_iarg_72_tready),
        .s_axis_iarg_73_aclk(s_axis_iarg_73_aclk),
        .s_axis_iarg_73_aresetn(s_axis_iarg_73_aresetn),
        .s_axis_iarg_73_tlast(s_axis_iarg_73_tlast),
        .s_axis_iarg_73_tvalid(s_axis_iarg_73_tvalid),
        .s_axis_iarg_73_tkeep(s_axis_iarg_73_tkeep),
        .s_axis_iarg_73_tstrb(s_axis_iarg_73_tstrb),
        .s_axis_iarg_73_tdata(s_axis_iarg_73_tdata),
        .s_axis_iarg_73_tready(s_axis_iarg_73_tready),
        .ap_axis_iarg_73_tlast(ap_axis_iarg_73_tlast),
        .ap_axis_iarg_73_tvalid(ap_axis_iarg_73_tvalid),
        .ap_axis_iarg_73_tkeep(ap_axis_iarg_73_tkeep),
        .ap_axis_iarg_73_tstrb(ap_axis_iarg_73_tstrb),
        .ap_axis_iarg_73_tdata(ap_axis_iarg_73_tdata),
        .ap_axis_iarg_73_tready(ap_axis_iarg_73_tready),
        .s_axis_iarg_74_aclk(s_axis_iarg_74_aclk),
        .s_axis_iarg_74_aresetn(s_axis_iarg_74_aresetn),
        .s_axis_iarg_74_tlast(s_axis_iarg_74_tlast),
        .s_axis_iarg_74_tvalid(s_axis_iarg_74_tvalid),
        .s_axis_iarg_74_tkeep(s_axis_iarg_74_tkeep),
        .s_axis_iarg_74_tstrb(s_axis_iarg_74_tstrb),
        .s_axis_iarg_74_tdata(s_axis_iarg_74_tdata),
        .s_axis_iarg_74_tready(s_axis_iarg_74_tready),
        .ap_axis_iarg_74_tlast(ap_axis_iarg_74_tlast),
        .ap_axis_iarg_74_tvalid(ap_axis_iarg_74_tvalid),
        .ap_axis_iarg_74_tkeep(ap_axis_iarg_74_tkeep),
        .ap_axis_iarg_74_tstrb(ap_axis_iarg_74_tstrb),
        .ap_axis_iarg_74_tdata(ap_axis_iarg_74_tdata),
        .ap_axis_iarg_74_tready(ap_axis_iarg_74_tready),
        .s_axis_iarg_75_aclk(s_axis_iarg_75_aclk),
        .s_axis_iarg_75_aresetn(s_axis_iarg_75_aresetn),
        .s_axis_iarg_75_tlast(s_axis_iarg_75_tlast),
        .s_axis_iarg_75_tvalid(s_axis_iarg_75_tvalid),
        .s_axis_iarg_75_tkeep(s_axis_iarg_75_tkeep),
        .s_axis_iarg_75_tstrb(s_axis_iarg_75_tstrb),
        .s_axis_iarg_75_tdata(s_axis_iarg_75_tdata),
        .s_axis_iarg_75_tready(s_axis_iarg_75_tready),
        .ap_axis_iarg_75_tlast(ap_axis_iarg_75_tlast),
        .ap_axis_iarg_75_tvalid(ap_axis_iarg_75_tvalid),
        .ap_axis_iarg_75_tkeep(ap_axis_iarg_75_tkeep),
        .ap_axis_iarg_75_tstrb(ap_axis_iarg_75_tstrb),
        .ap_axis_iarg_75_tdata(ap_axis_iarg_75_tdata),
        .ap_axis_iarg_75_tready(ap_axis_iarg_75_tready),
        .s_axis_iarg_76_aclk(s_axis_iarg_76_aclk),
        .s_axis_iarg_76_aresetn(s_axis_iarg_76_aresetn),
        .s_axis_iarg_76_tlast(s_axis_iarg_76_tlast),
        .s_axis_iarg_76_tvalid(s_axis_iarg_76_tvalid),
        .s_axis_iarg_76_tkeep(s_axis_iarg_76_tkeep),
        .s_axis_iarg_76_tstrb(s_axis_iarg_76_tstrb),
        .s_axis_iarg_76_tdata(s_axis_iarg_76_tdata),
        .s_axis_iarg_76_tready(s_axis_iarg_76_tready),
        .ap_axis_iarg_76_tlast(ap_axis_iarg_76_tlast),
        .ap_axis_iarg_76_tvalid(ap_axis_iarg_76_tvalid),
        .ap_axis_iarg_76_tkeep(ap_axis_iarg_76_tkeep),
        .ap_axis_iarg_76_tstrb(ap_axis_iarg_76_tstrb),
        .ap_axis_iarg_76_tdata(ap_axis_iarg_76_tdata),
        .ap_axis_iarg_76_tready(ap_axis_iarg_76_tready),
        .s_axis_iarg_77_aclk(s_axis_iarg_77_aclk),
        .s_axis_iarg_77_aresetn(s_axis_iarg_77_aresetn),
        .s_axis_iarg_77_tlast(s_axis_iarg_77_tlast),
        .s_axis_iarg_77_tvalid(s_axis_iarg_77_tvalid),
        .s_axis_iarg_77_tkeep(s_axis_iarg_77_tkeep),
        .s_axis_iarg_77_tstrb(s_axis_iarg_77_tstrb),
        .s_axis_iarg_77_tdata(s_axis_iarg_77_tdata),
        .s_axis_iarg_77_tready(s_axis_iarg_77_tready),
        .ap_axis_iarg_77_tlast(ap_axis_iarg_77_tlast),
        .ap_axis_iarg_77_tvalid(ap_axis_iarg_77_tvalid),
        .ap_axis_iarg_77_tkeep(ap_axis_iarg_77_tkeep),
        .ap_axis_iarg_77_tstrb(ap_axis_iarg_77_tstrb),
        .ap_axis_iarg_77_tdata(ap_axis_iarg_77_tdata),
        .ap_axis_iarg_77_tready(ap_axis_iarg_77_tready),
        .s_axis_iarg_78_aclk(s_axis_iarg_78_aclk),
        .s_axis_iarg_78_aresetn(s_axis_iarg_78_aresetn),
        .s_axis_iarg_78_tlast(s_axis_iarg_78_tlast),
        .s_axis_iarg_78_tvalid(s_axis_iarg_78_tvalid),
        .s_axis_iarg_78_tkeep(s_axis_iarg_78_tkeep),
        .s_axis_iarg_78_tstrb(s_axis_iarg_78_tstrb),
        .s_axis_iarg_78_tdata(s_axis_iarg_78_tdata),
        .s_axis_iarg_78_tready(s_axis_iarg_78_tready),
        .ap_axis_iarg_78_tlast(ap_axis_iarg_78_tlast),
        .ap_axis_iarg_78_tvalid(ap_axis_iarg_78_tvalid),
        .ap_axis_iarg_78_tkeep(ap_axis_iarg_78_tkeep),
        .ap_axis_iarg_78_tstrb(ap_axis_iarg_78_tstrb),
        .ap_axis_iarg_78_tdata(ap_axis_iarg_78_tdata),
        .ap_axis_iarg_78_tready(ap_axis_iarg_78_tready),
        .s_axis_iarg_79_aclk(s_axis_iarg_79_aclk),
        .s_axis_iarg_79_aresetn(s_axis_iarg_79_aresetn),
        .s_axis_iarg_79_tlast(s_axis_iarg_79_tlast),
        .s_axis_iarg_79_tvalid(s_axis_iarg_79_tvalid),
        .s_axis_iarg_79_tkeep(s_axis_iarg_79_tkeep),
        .s_axis_iarg_79_tstrb(s_axis_iarg_79_tstrb),
        .s_axis_iarg_79_tdata(s_axis_iarg_79_tdata),
        .s_axis_iarg_79_tready(s_axis_iarg_79_tready),
        .ap_axis_iarg_79_tlast(ap_axis_iarg_79_tlast),
        .ap_axis_iarg_79_tvalid(ap_axis_iarg_79_tvalid),
        .ap_axis_iarg_79_tkeep(ap_axis_iarg_79_tkeep),
        .ap_axis_iarg_79_tstrb(ap_axis_iarg_79_tstrb),
        .ap_axis_iarg_79_tdata(ap_axis_iarg_79_tdata),
        .ap_axis_iarg_79_tready(ap_axis_iarg_79_tready),
        .s_axis_iarg_80_aclk(s_axis_iarg_80_aclk),
        .s_axis_iarg_80_aresetn(s_axis_iarg_80_aresetn),
        .s_axis_iarg_80_tlast(s_axis_iarg_80_tlast),
        .s_axis_iarg_80_tvalid(s_axis_iarg_80_tvalid),
        .s_axis_iarg_80_tkeep(s_axis_iarg_80_tkeep),
        .s_axis_iarg_80_tstrb(s_axis_iarg_80_tstrb),
        .s_axis_iarg_80_tdata(s_axis_iarg_80_tdata),
        .s_axis_iarg_80_tready(s_axis_iarg_80_tready),
        .ap_axis_iarg_80_tlast(ap_axis_iarg_80_tlast),
        .ap_axis_iarg_80_tvalid(ap_axis_iarg_80_tvalid),
        .ap_axis_iarg_80_tkeep(ap_axis_iarg_80_tkeep),
        .ap_axis_iarg_80_tstrb(ap_axis_iarg_80_tstrb),
        .ap_axis_iarg_80_tdata(ap_axis_iarg_80_tdata),
        .ap_axis_iarg_80_tready(ap_axis_iarg_80_tready),
        .s_axis_iarg_81_aclk(s_axis_iarg_81_aclk),
        .s_axis_iarg_81_aresetn(s_axis_iarg_81_aresetn),
        .s_axis_iarg_81_tlast(s_axis_iarg_81_tlast),
        .s_axis_iarg_81_tvalid(s_axis_iarg_81_tvalid),
        .s_axis_iarg_81_tkeep(s_axis_iarg_81_tkeep),
        .s_axis_iarg_81_tstrb(s_axis_iarg_81_tstrb),
        .s_axis_iarg_81_tdata(s_axis_iarg_81_tdata),
        .s_axis_iarg_81_tready(s_axis_iarg_81_tready),
        .ap_axis_iarg_81_tlast(ap_axis_iarg_81_tlast),
        .ap_axis_iarg_81_tvalid(ap_axis_iarg_81_tvalid),
        .ap_axis_iarg_81_tkeep(ap_axis_iarg_81_tkeep),
        .ap_axis_iarg_81_tstrb(ap_axis_iarg_81_tstrb),
        .ap_axis_iarg_81_tdata(ap_axis_iarg_81_tdata),
        .ap_axis_iarg_81_tready(ap_axis_iarg_81_tready),
        .s_axis_iarg_82_aclk(s_axis_iarg_82_aclk),
        .s_axis_iarg_82_aresetn(s_axis_iarg_82_aresetn),
        .s_axis_iarg_82_tlast(s_axis_iarg_82_tlast),
        .s_axis_iarg_82_tvalid(s_axis_iarg_82_tvalid),
        .s_axis_iarg_82_tkeep(s_axis_iarg_82_tkeep),
        .s_axis_iarg_82_tstrb(s_axis_iarg_82_tstrb),
        .s_axis_iarg_82_tdata(s_axis_iarg_82_tdata),
        .s_axis_iarg_82_tready(s_axis_iarg_82_tready),
        .ap_axis_iarg_82_tlast(ap_axis_iarg_82_tlast),
        .ap_axis_iarg_82_tvalid(ap_axis_iarg_82_tvalid),
        .ap_axis_iarg_82_tkeep(ap_axis_iarg_82_tkeep),
        .ap_axis_iarg_82_tstrb(ap_axis_iarg_82_tstrb),
        .ap_axis_iarg_82_tdata(ap_axis_iarg_82_tdata),
        .ap_axis_iarg_82_tready(ap_axis_iarg_82_tready),
        .s_axis_iarg_83_aclk(s_axis_iarg_83_aclk),
        .s_axis_iarg_83_aresetn(s_axis_iarg_83_aresetn),
        .s_axis_iarg_83_tlast(s_axis_iarg_83_tlast),
        .s_axis_iarg_83_tvalid(s_axis_iarg_83_tvalid),
        .s_axis_iarg_83_tkeep(s_axis_iarg_83_tkeep),
        .s_axis_iarg_83_tstrb(s_axis_iarg_83_tstrb),
        .s_axis_iarg_83_tdata(s_axis_iarg_83_tdata),
        .s_axis_iarg_83_tready(s_axis_iarg_83_tready),
        .ap_axis_iarg_83_tlast(ap_axis_iarg_83_tlast),
        .ap_axis_iarg_83_tvalid(ap_axis_iarg_83_tvalid),
        .ap_axis_iarg_83_tkeep(ap_axis_iarg_83_tkeep),
        .ap_axis_iarg_83_tstrb(ap_axis_iarg_83_tstrb),
        .ap_axis_iarg_83_tdata(ap_axis_iarg_83_tdata),
        .ap_axis_iarg_83_tready(ap_axis_iarg_83_tready),
        .s_axis_iarg_84_aclk(s_axis_iarg_84_aclk),
        .s_axis_iarg_84_aresetn(s_axis_iarg_84_aresetn),
        .s_axis_iarg_84_tlast(s_axis_iarg_84_tlast),
        .s_axis_iarg_84_tvalid(s_axis_iarg_84_tvalid),
        .s_axis_iarg_84_tkeep(s_axis_iarg_84_tkeep),
        .s_axis_iarg_84_tstrb(s_axis_iarg_84_tstrb),
        .s_axis_iarg_84_tdata(s_axis_iarg_84_tdata),
        .s_axis_iarg_84_tready(s_axis_iarg_84_tready),
        .ap_axis_iarg_84_tlast(ap_axis_iarg_84_tlast),
        .ap_axis_iarg_84_tvalid(ap_axis_iarg_84_tvalid),
        .ap_axis_iarg_84_tkeep(ap_axis_iarg_84_tkeep),
        .ap_axis_iarg_84_tstrb(ap_axis_iarg_84_tstrb),
        .ap_axis_iarg_84_tdata(ap_axis_iarg_84_tdata),
        .ap_axis_iarg_84_tready(ap_axis_iarg_84_tready),
        .s_axis_iarg_85_aclk(s_axis_iarg_85_aclk),
        .s_axis_iarg_85_aresetn(s_axis_iarg_85_aresetn),
        .s_axis_iarg_85_tlast(s_axis_iarg_85_tlast),
        .s_axis_iarg_85_tvalid(s_axis_iarg_85_tvalid),
        .s_axis_iarg_85_tkeep(s_axis_iarg_85_tkeep),
        .s_axis_iarg_85_tstrb(s_axis_iarg_85_tstrb),
        .s_axis_iarg_85_tdata(s_axis_iarg_85_tdata),
        .s_axis_iarg_85_tready(s_axis_iarg_85_tready),
        .ap_axis_iarg_85_tlast(ap_axis_iarg_85_tlast),
        .ap_axis_iarg_85_tvalid(ap_axis_iarg_85_tvalid),
        .ap_axis_iarg_85_tkeep(ap_axis_iarg_85_tkeep),
        .ap_axis_iarg_85_tstrb(ap_axis_iarg_85_tstrb),
        .ap_axis_iarg_85_tdata(ap_axis_iarg_85_tdata),
        .ap_axis_iarg_85_tready(ap_axis_iarg_85_tready),
        .s_axis_iarg_86_aclk(s_axis_iarg_86_aclk),
        .s_axis_iarg_86_aresetn(s_axis_iarg_86_aresetn),
        .s_axis_iarg_86_tlast(s_axis_iarg_86_tlast),
        .s_axis_iarg_86_tvalid(s_axis_iarg_86_tvalid),
        .s_axis_iarg_86_tkeep(s_axis_iarg_86_tkeep),
        .s_axis_iarg_86_tstrb(s_axis_iarg_86_tstrb),
        .s_axis_iarg_86_tdata(s_axis_iarg_86_tdata),
        .s_axis_iarg_86_tready(s_axis_iarg_86_tready),
        .ap_axis_iarg_86_tlast(ap_axis_iarg_86_tlast),
        .ap_axis_iarg_86_tvalid(ap_axis_iarg_86_tvalid),
        .ap_axis_iarg_86_tkeep(ap_axis_iarg_86_tkeep),
        .ap_axis_iarg_86_tstrb(ap_axis_iarg_86_tstrb),
        .ap_axis_iarg_86_tdata(ap_axis_iarg_86_tdata),
        .ap_axis_iarg_86_tready(ap_axis_iarg_86_tready),
        .s_axis_iarg_87_aclk(s_axis_iarg_87_aclk),
        .s_axis_iarg_87_aresetn(s_axis_iarg_87_aresetn),
        .s_axis_iarg_87_tlast(s_axis_iarg_87_tlast),
        .s_axis_iarg_87_tvalid(s_axis_iarg_87_tvalid),
        .s_axis_iarg_87_tkeep(s_axis_iarg_87_tkeep),
        .s_axis_iarg_87_tstrb(s_axis_iarg_87_tstrb),
        .s_axis_iarg_87_tdata(s_axis_iarg_87_tdata),
        .s_axis_iarg_87_tready(s_axis_iarg_87_tready),
        .ap_axis_iarg_87_tlast(ap_axis_iarg_87_tlast),
        .ap_axis_iarg_87_tvalid(ap_axis_iarg_87_tvalid),
        .ap_axis_iarg_87_tkeep(ap_axis_iarg_87_tkeep),
        .ap_axis_iarg_87_tstrb(ap_axis_iarg_87_tstrb),
        .ap_axis_iarg_87_tdata(ap_axis_iarg_87_tdata),
        .ap_axis_iarg_87_tready(ap_axis_iarg_87_tready),
        .s_axis_iarg_88_aclk(s_axis_iarg_88_aclk),
        .s_axis_iarg_88_aresetn(s_axis_iarg_88_aresetn),
        .s_axis_iarg_88_tlast(s_axis_iarg_88_tlast),
        .s_axis_iarg_88_tvalid(s_axis_iarg_88_tvalid),
        .s_axis_iarg_88_tkeep(s_axis_iarg_88_tkeep),
        .s_axis_iarg_88_tstrb(s_axis_iarg_88_tstrb),
        .s_axis_iarg_88_tdata(s_axis_iarg_88_tdata),
        .s_axis_iarg_88_tready(s_axis_iarg_88_tready),
        .ap_axis_iarg_88_tlast(ap_axis_iarg_88_tlast),
        .ap_axis_iarg_88_tvalid(ap_axis_iarg_88_tvalid),
        .ap_axis_iarg_88_tkeep(ap_axis_iarg_88_tkeep),
        .ap_axis_iarg_88_tstrb(ap_axis_iarg_88_tstrb),
        .ap_axis_iarg_88_tdata(ap_axis_iarg_88_tdata),
        .ap_axis_iarg_88_tready(ap_axis_iarg_88_tready),
        .s_axis_iarg_89_aclk(s_axis_iarg_89_aclk),
        .s_axis_iarg_89_aresetn(s_axis_iarg_89_aresetn),
        .s_axis_iarg_89_tlast(s_axis_iarg_89_tlast),
        .s_axis_iarg_89_tvalid(s_axis_iarg_89_tvalid),
        .s_axis_iarg_89_tkeep(s_axis_iarg_89_tkeep),
        .s_axis_iarg_89_tstrb(s_axis_iarg_89_tstrb),
        .s_axis_iarg_89_tdata(s_axis_iarg_89_tdata),
        .s_axis_iarg_89_tready(s_axis_iarg_89_tready),
        .ap_axis_iarg_89_tlast(ap_axis_iarg_89_tlast),
        .ap_axis_iarg_89_tvalid(ap_axis_iarg_89_tvalid),
        .ap_axis_iarg_89_tkeep(ap_axis_iarg_89_tkeep),
        .ap_axis_iarg_89_tstrb(ap_axis_iarg_89_tstrb),
        .ap_axis_iarg_89_tdata(ap_axis_iarg_89_tdata),
        .ap_axis_iarg_89_tready(ap_axis_iarg_89_tready),
        .s_axis_iarg_90_aclk(s_axis_iarg_90_aclk),
        .s_axis_iarg_90_aresetn(s_axis_iarg_90_aresetn),
        .s_axis_iarg_90_tlast(s_axis_iarg_90_tlast),
        .s_axis_iarg_90_tvalid(s_axis_iarg_90_tvalid),
        .s_axis_iarg_90_tkeep(s_axis_iarg_90_tkeep),
        .s_axis_iarg_90_tstrb(s_axis_iarg_90_tstrb),
        .s_axis_iarg_90_tdata(s_axis_iarg_90_tdata),
        .s_axis_iarg_90_tready(s_axis_iarg_90_tready),
        .ap_axis_iarg_90_tlast(ap_axis_iarg_90_tlast),
        .ap_axis_iarg_90_tvalid(ap_axis_iarg_90_tvalid),
        .ap_axis_iarg_90_tkeep(ap_axis_iarg_90_tkeep),
        .ap_axis_iarg_90_tstrb(ap_axis_iarg_90_tstrb),
        .ap_axis_iarg_90_tdata(ap_axis_iarg_90_tdata),
        .ap_axis_iarg_90_tready(ap_axis_iarg_90_tready),
        .s_axis_iarg_91_aclk(s_axis_iarg_91_aclk),
        .s_axis_iarg_91_aresetn(s_axis_iarg_91_aresetn),
        .s_axis_iarg_91_tlast(s_axis_iarg_91_tlast),
        .s_axis_iarg_91_tvalid(s_axis_iarg_91_tvalid),
        .s_axis_iarg_91_tkeep(s_axis_iarg_91_tkeep),
        .s_axis_iarg_91_tstrb(s_axis_iarg_91_tstrb),
        .s_axis_iarg_91_tdata(s_axis_iarg_91_tdata),
        .s_axis_iarg_91_tready(s_axis_iarg_91_tready),
        .ap_axis_iarg_91_tlast(ap_axis_iarg_91_tlast),
        .ap_axis_iarg_91_tvalid(ap_axis_iarg_91_tvalid),
        .ap_axis_iarg_91_tkeep(ap_axis_iarg_91_tkeep),
        .ap_axis_iarg_91_tstrb(ap_axis_iarg_91_tstrb),
        .ap_axis_iarg_91_tdata(ap_axis_iarg_91_tdata),
        .ap_axis_iarg_91_tready(ap_axis_iarg_91_tready),
        .s_axis_iarg_92_aclk(s_axis_iarg_92_aclk),
        .s_axis_iarg_92_aresetn(s_axis_iarg_92_aresetn),
        .s_axis_iarg_92_tlast(s_axis_iarg_92_tlast),
        .s_axis_iarg_92_tvalid(s_axis_iarg_92_tvalid),
        .s_axis_iarg_92_tkeep(s_axis_iarg_92_tkeep),
        .s_axis_iarg_92_tstrb(s_axis_iarg_92_tstrb),
        .s_axis_iarg_92_tdata(s_axis_iarg_92_tdata),
        .s_axis_iarg_92_tready(s_axis_iarg_92_tready),
        .ap_axis_iarg_92_tlast(ap_axis_iarg_92_tlast),
        .ap_axis_iarg_92_tvalid(ap_axis_iarg_92_tvalid),
        .ap_axis_iarg_92_tkeep(ap_axis_iarg_92_tkeep),
        .ap_axis_iarg_92_tstrb(ap_axis_iarg_92_tstrb),
        .ap_axis_iarg_92_tdata(ap_axis_iarg_92_tdata),
        .ap_axis_iarg_92_tready(ap_axis_iarg_92_tready),
        .s_axis_iarg_93_aclk(s_axis_iarg_93_aclk),
        .s_axis_iarg_93_aresetn(s_axis_iarg_93_aresetn),
        .s_axis_iarg_93_tlast(s_axis_iarg_93_tlast),
        .s_axis_iarg_93_tvalid(s_axis_iarg_93_tvalid),
        .s_axis_iarg_93_tkeep(s_axis_iarg_93_tkeep),
        .s_axis_iarg_93_tstrb(s_axis_iarg_93_tstrb),
        .s_axis_iarg_93_tdata(s_axis_iarg_93_tdata),
        .s_axis_iarg_93_tready(s_axis_iarg_93_tready),
        .ap_axis_iarg_93_tlast(ap_axis_iarg_93_tlast),
        .ap_axis_iarg_93_tvalid(ap_axis_iarg_93_tvalid),
        .ap_axis_iarg_93_tkeep(ap_axis_iarg_93_tkeep),
        .ap_axis_iarg_93_tstrb(ap_axis_iarg_93_tstrb),
        .ap_axis_iarg_93_tdata(ap_axis_iarg_93_tdata),
        .ap_axis_iarg_93_tready(ap_axis_iarg_93_tready),
        .s_axis_iarg_94_aclk(s_axis_iarg_94_aclk),
        .s_axis_iarg_94_aresetn(s_axis_iarg_94_aresetn),
        .s_axis_iarg_94_tlast(s_axis_iarg_94_tlast),
        .s_axis_iarg_94_tvalid(s_axis_iarg_94_tvalid),
        .s_axis_iarg_94_tkeep(s_axis_iarg_94_tkeep),
        .s_axis_iarg_94_tstrb(s_axis_iarg_94_tstrb),
        .s_axis_iarg_94_tdata(s_axis_iarg_94_tdata),
        .s_axis_iarg_94_tready(s_axis_iarg_94_tready),
        .ap_axis_iarg_94_tlast(ap_axis_iarg_94_tlast),
        .ap_axis_iarg_94_tvalid(ap_axis_iarg_94_tvalid),
        .ap_axis_iarg_94_tkeep(ap_axis_iarg_94_tkeep),
        .ap_axis_iarg_94_tstrb(ap_axis_iarg_94_tstrb),
        .ap_axis_iarg_94_tdata(ap_axis_iarg_94_tdata),
        .ap_axis_iarg_94_tready(ap_axis_iarg_94_tready),
        .s_axis_iarg_95_aclk(s_axis_iarg_95_aclk),
        .s_axis_iarg_95_aresetn(s_axis_iarg_95_aresetn),
        .s_axis_iarg_95_tlast(s_axis_iarg_95_tlast),
        .s_axis_iarg_95_tvalid(s_axis_iarg_95_tvalid),
        .s_axis_iarg_95_tkeep(s_axis_iarg_95_tkeep),
        .s_axis_iarg_95_tstrb(s_axis_iarg_95_tstrb),
        .s_axis_iarg_95_tdata(s_axis_iarg_95_tdata),
        .s_axis_iarg_95_tready(s_axis_iarg_95_tready),
        .ap_axis_iarg_95_tlast(ap_axis_iarg_95_tlast),
        .ap_axis_iarg_95_tvalid(ap_axis_iarg_95_tvalid),
        .ap_axis_iarg_95_tkeep(ap_axis_iarg_95_tkeep),
        .ap_axis_iarg_95_tstrb(ap_axis_iarg_95_tstrb),
        .ap_axis_iarg_95_tdata(ap_axis_iarg_95_tdata),
        .ap_axis_iarg_95_tready(ap_axis_iarg_95_tready),
        .s_axis_iarg_96_aclk(s_axis_iarg_96_aclk),
        .s_axis_iarg_96_aresetn(s_axis_iarg_96_aresetn),
        .s_axis_iarg_96_tlast(s_axis_iarg_96_tlast),
        .s_axis_iarg_96_tvalid(s_axis_iarg_96_tvalid),
        .s_axis_iarg_96_tkeep(s_axis_iarg_96_tkeep),
        .s_axis_iarg_96_tstrb(s_axis_iarg_96_tstrb),
        .s_axis_iarg_96_tdata(s_axis_iarg_96_tdata),
        .s_axis_iarg_96_tready(s_axis_iarg_96_tready),
        .ap_axis_iarg_96_tlast(ap_axis_iarg_96_tlast),
        .ap_axis_iarg_96_tvalid(ap_axis_iarg_96_tvalid),
        .ap_axis_iarg_96_tkeep(ap_axis_iarg_96_tkeep),
        .ap_axis_iarg_96_tstrb(ap_axis_iarg_96_tstrb),
        .ap_axis_iarg_96_tdata(ap_axis_iarg_96_tdata),
        .ap_axis_iarg_96_tready(ap_axis_iarg_96_tready),
        .s_axis_iarg_97_aclk(s_axis_iarg_97_aclk),
        .s_axis_iarg_97_aresetn(s_axis_iarg_97_aresetn),
        .s_axis_iarg_97_tlast(s_axis_iarg_97_tlast),
        .s_axis_iarg_97_tvalid(s_axis_iarg_97_tvalid),
        .s_axis_iarg_97_tkeep(s_axis_iarg_97_tkeep),
        .s_axis_iarg_97_tstrb(s_axis_iarg_97_tstrb),
        .s_axis_iarg_97_tdata(s_axis_iarg_97_tdata),
        .s_axis_iarg_97_tready(s_axis_iarg_97_tready),
        .ap_axis_iarg_97_tlast(ap_axis_iarg_97_tlast),
        .ap_axis_iarg_97_tvalid(ap_axis_iarg_97_tvalid),
        .ap_axis_iarg_97_tkeep(ap_axis_iarg_97_tkeep),
        .ap_axis_iarg_97_tstrb(ap_axis_iarg_97_tstrb),
        .ap_axis_iarg_97_tdata(ap_axis_iarg_97_tdata),
        .ap_axis_iarg_97_tready(ap_axis_iarg_97_tready),
        .s_axis_iarg_98_aclk(s_axis_iarg_98_aclk),
        .s_axis_iarg_98_aresetn(s_axis_iarg_98_aresetn),
        .s_axis_iarg_98_tlast(s_axis_iarg_98_tlast),
        .s_axis_iarg_98_tvalid(s_axis_iarg_98_tvalid),
        .s_axis_iarg_98_tkeep(s_axis_iarg_98_tkeep),
        .s_axis_iarg_98_tstrb(s_axis_iarg_98_tstrb),
        .s_axis_iarg_98_tdata(s_axis_iarg_98_tdata),
        .s_axis_iarg_98_tready(s_axis_iarg_98_tready),
        .ap_axis_iarg_98_tlast(ap_axis_iarg_98_tlast),
        .ap_axis_iarg_98_tvalid(ap_axis_iarg_98_tvalid),
        .ap_axis_iarg_98_tkeep(ap_axis_iarg_98_tkeep),
        .ap_axis_iarg_98_tstrb(ap_axis_iarg_98_tstrb),
        .ap_axis_iarg_98_tdata(ap_axis_iarg_98_tdata),
        .ap_axis_iarg_98_tready(ap_axis_iarg_98_tready),
        .s_axis_iarg_99_aclk(s_axis_iarg_99_aclk),
        .s_axis_iarg_99_aresetn(s_axis_iarg_99_aresetn),
        .s_axis_iarg_99_tlast(s_axis_iarg_99_tlast),
        .s_axis_iarg_99_tvalid(s_axis_iarg_99_tvalid),
        .s_axis_iarg_99_tkeep(s_axis_iarg_99_tkeep),
        .s_axis_iarg_99_tstrb(s_axis_iarg_99_tstrb),
        .s_axis_iarg_99_tdata(s_axis_iarg_99_tdata),
        .s_axis_iarg_99_tready(s_axis_iarg_99_tready),
        .ap_axis_iarg_99_tlast(ap_axis_iarg_99_tlast),
        .ap_axis_iarg_99_tvalid(ap_axis_iarg_99_tvalid),
        .ap_axis_iarg_99_tkeep(ap_axis_iarg_99_tkeep),
        .ap_axis_iarg_99_tstrb(ap_axis_iarg_99_tstrb),
        .ap_axis_iarg_99_tdata(ap_axis_iarg_99_tdata),
        .ap_axis_iarg_99_tready(ap_axis_iarg_99_tready),
        .s_axis_iarg_100_aclk(s_axis_iarg_100_aclk),
        .s_axis_iarg_100_aresetn(s_axis_iarg_100_aresetn),
        .s_axis_iarg_100_tlast(s_axis_iarg_100_tlast),
        .s_axis_iarg_100_tvalid(s_axis_iarg_100_tvalid),
        .s_axis_iarg_100_tkeep(s_axis_iarg_100_tkeep),
        .s_axis_iarg_100_tstrb(s_axis_iarg_100_tstrb),
        .s_axis_iarg_100_tdata(s_axis_iarg_100_tdata),
        .s_axis_iarg_100_tready(s_axis_iarg_100_tready),
        .ap_axis_iarg_100_tlast(ap_axis_iarg_100_tlast),
        .ap_axis_iarg_100_tvalid(ap_axis_iarg_100_tvalid),
        .ap_axis_iarg_100_tkeep(ap_axis_iarg_100_tkeep),
        .ap_axis_iarg_100_tstrb(ap_axis_iarg_100_tstrb),
        .ap_axis_iarg_100_tdata(ap_axis_iarg_100_tdata),
        .ap_axis_iarg_100_tready(ap_axis_iarg_100_tready),
        .s_axis_iarg_101_aclk(s_axis_iarg_101_aclk),
        .s_axis_iarg_101_aresetn(s_axis_iarg_101_aresetn),
        .s_axis_iarg_101_tlast(s_axis_iarg_101_tlast),
        .s_axis_iarg_101_tvalid(s_axis_iarg_101_tvalid),
        .s_axis_iarg_101_tkeep(s_axis_iarg_101_tkeep),
        .s_axis_iarg_101_tstrb(s_axis_iarg_101_tstrb),
        .s_axis_iarg_101_tdata(s_axis_iarg_101_tdata),
        .s_axis_iarg_101_tready(s_axis_iarg_101_tready),
        .ap_axis_iarg_101_tlast(ap_axis_iarg_101_tlast),
        .ap_axis_iarg_101_tvalid(ap_axis_iarg_101_tvalid),
        .ap_axis_iarg_101_tkeep(ap_axis_iarg_101_tkeep),
        .ap_axis_iarg_101_tstrb(ap_axis_iarg_101_tstrb),
        .ap_axis_iarg_101_tdata(ap_axis_iarg_101_tdata),
        .ap_axis_iarg_101_tready(ap_axis_iarg_101_tready),
        .s_axis_iarg_102_aclk(s_axis_iarg_102_aclk),
        .s_axis_iarg_102_aresetn(s_axis_iarg_102_aresetn),
        .s_axis_iarg_102_tlast(s_axis_iarg_102_tlast),
        .s_axis_iarg_102_tvalid(s_axis_iarg_102_tvalid),
        .s_axis_iarg_102_tkeep(s_axis_iarg_102_tkeep),
        .s_axis_iarg_102_tstrb(s_axis_iarg_102_tstrb),
        .s_axis_iarg_102_tdata(s_axis_iarg_102_tdata),
        .s_axis_iarg_102_tready(s_axis_iarg_102_tready),
        .ap_axis_iarg_102_tlast(ap_axis_iarg_102_tlast),
        .ap_axis_iarg_102_tvalid(ap_axis_iarg_102_tvalid),
        .ap_axis_iarg_102_tkeep(ap_axis_iarg_102_tkeep),
        .ap_axis_iarg_102_tstrb(ap_axis_iarg_102_tstrb),
        .ap_axis_iarg_102_tdata(ap_axis_iarg_102_tdata),
        .ap_axis_iarg_102_tready(ap_axis_iarg_102_tready),
        .s_axis_iarg_103_aclk(s_axis_iarg_103_aclk),
        .s_axis_iarg_103_aresetn(s_axis_iarg_103_aresetn),
        .s_axis_iarg_103_tlast(s_axis_iarg_103_tlast),
        .s_axis_iarg_103_tvalid(s_axis_iarg_103_tvalid),
        .s_axis_iarg_103_tkeep(s_axis_iarg_103_tkeep),
        .s_axis_iarg_103_tstrb(s_axis_iarg_103_tstrb),
        .s_axis_iarg_103_tdata(s_axis_iarg_103_tdata),
        .s_axis_iarg_103_tready(s_axis_iarg_103_tready),
        .ap_axis_iarg_103_tlast(ap_axis_iarg_103_tlast),
        .ap_axis_iarg_103_tvalid(ap_axis_iarg_103_tvalid),
        .ap_axis_iarg_103_tkeep(ap_axis_iarg_103_tkeep),
        .ap_axis_iarg_103_tstrb(ap_axis_iarg_103_tstrb),
        .ap_axis_iarg_103_tdata(ap_axis_iarg_103_tdata),
        .ap_axis_iarg_103_tready(ap_axis_iarg_103_tready),
        .s_axis_iarg_104_aclk(s_axis_iarg_104_aclk),
        .s_axis_iarg_104_aresetn(s_axis_iarg_104_aresetn),
        .s_axis_iarg_104_tlast(s_axis_iarg_104_tlast),
        .s_axis_iarg_104_tvalid(s_axis_iarg_104_tvalid),
        .s_axis_iarg_104_tkeep(s_axis_iarg_104_tkeep),
        .s_axis_iarg_104_tstrb(s_axis_iarg_104_tstrb),
        .s_axis_iarg_104_tdata(s_axis_iarg_104_tdata),
        .s_axis_iarg_104_tready(s_axis_iarg_104_tready),
        .ap_axis_iarg_104_tlast(ap_axis_iarg_104_tlast),
        .ap_axis_iarg_104_tvalid(ap_axis_iarg_104_tvalid),
        .ap_axis_iarg_104_tkeep(ap_axis_iarg_104_tkeep),
        .ap_axis_iarg_104_tstrb(ap_axis_iarg_104_tstrb),
        .ap_axis_iarg_104_tdata(ap_axis_iarg_104_tdata),
        .ap_axis_iarg_104_tready(ap_axis_iarg_104_tready),
        .s_axis_iarg_105_aclk(s_axis_iarg_105_aclk),
        .s_axis_iarg_105_aresetn(s_axis_iarg_105_aresetn),
        .s_axis_iarg_105_tlast(s_axis_iarg_105_tlast),
        .s_axis_iarg_105_tvalid(s_axis_iarg_105_tvalid),
        .s_axis_iarg_105_tkeep(s_axis_iarg_105_tkeep),
        .s_axis_iarg_105_tstrb(s_axis_iarg_105_tstrb),
        .s_axis_iarg_105_tdata(s_axis_iarg_105_tdata),
        .s_axis_iarg_105_tready(s_axis_iarg_105_tready),
        .ap_axis_iarg_105_tlast(ap_axis_iarg_105_tlast),
        .ap_axis_iarg_105_tvalid(ap_axis_iarg_105_tvalid),
        .ap_axis_iarg_105_tkeep(ap_axis_iarg_105_tkeep),
        .ap_axis_iarg_105_tstrb(ap_axis_iarg_105_tstrb),
        .ap_axis_iarg_105_tdata(ap_axis_iarg_105_tdata),
        .ap_axis_iarg_105_tready(ap_axis_iarg_105_tready),
        .s_axis_iarg_106_aclk(s_axis_iarg_106_aclk),
        .s_axis_iarg_106_aresetn(s_axis_iarg_106_aresetn),
        .s_axis_iarg_106_tlast(s_axis_iarg_106_tlast),
        .s_axis_iarg_106_tvalid(s_axis_iarg_106_tvalid),
        .s_axis_iarg_106_tkeep(s_axis_iarg_106_tkeep),
        .s_axis_iarg_106_tstrb(s_axis_iarg_106_tstrb),
        .s_axis_iarg_106_tdata(s_axis_iarg_106_tdata),
        .s_axis_iarg_106_tready(s_axis_iarg_106_tready),
        .ap_axis_iarg_106_tlast(ap_axis_iarg_106_tlast),
        .ap_axis_iarg_106_tvalid(ap_axis_iarg_106_tvalid),
        .ap_axis_iarg_106_tkeep(ap_axis_iarg_106_tkeep),
        .ap_axis_iarg_106_tstrb(ap_axis_iarg_106_tstrb),
        .ap_axis_iarg_106_tdata(ap_axis_iarg_106_tdata),
        .ap_axis_iarg_106_tready(ap_axis_iarg_106_tready),
        .s_axis_iarg_107_aclk(s_axis_iarg_107_aclk),
        .s_axis_iarg_107_aresetn(s_axis_iarg_107_aresetn),
        .s_axis_iarg_107_tlast(s_axis_iarg_107_tlast),
        .s_axis_iarg_107_tvalid(s_axis_iarg_107_tvalid),
        .s_axis_iarg_107_tkeep(s_axis_iarg_107_tkeep),
        .s_axis_iarg_107_tstrb(s_axis_iarg_107_tstrb),
        .s_axis_iarg_107_tdata(s_axis_iarg_107_tdata),
        .s_axis_iarg_107_tready(s_axis_iarg_107_tready),
        .ap_axis_iarg_107_tlast(ap_axis_iarg_107_tlast),
        .ap_axis_iarg_107_tvalid(ap_axis_iarg_107_tvalid),
        .ap_axis_iarg_107_tkeep(ap_axis_iarg_107_tkeep),
        .ap_axis_iarg_107_tstrb(ap_axis_iarg_107_tstrb),
        .ap_axis_iarg_107_tdata(ap_axis_iarg_107_tdata),
        .ap_axis_iarg_107_tready(ap_axis_iarg_107_tready),
        .s_axis_iarg_108_aclk(s_axis_iarg_108_aclk),
        .s_axis_iarg_108_aresetn(s_axis_iarg_108_aresetn),
        .s_axis_iarg_108_tlast(s_axis_iarg_108_tlast),
        .s_axis_iarg_108_tvalid(s_axis_iarg_108_tvalid),
        .s_axis_iarg_108_tkeep(s_axis_iarg_108_tkeep),
        .s_axis_iarg_108_tstrb(s_axis_iarg_108_tstrb),
        .s_axis_iarg_108_tdata(s_axis_iarg_108_tdata),
        .s_axis_iarg_108_tready(s_axis_iarg_108_tready),
        .ap_axis_iarg_108_tlast(ap_axis_iarg_108_tlast),
        .ap_axis_iarg_108_tvalid(ap_axis_iarg_108_tvalid),
        .ap_axis_iarg_108_tkeep(ap_axis_iarg_108_tkeep),
        .ap_axis_iarg_108_tstrb(ap_axis_iarg_108_tstrb),
        .ap_axis_iarg_108_tdata(ap_axis_iarg_108_tdata),
        .ap_axis_iarg_108_tready(ap_axis_iarg_108_tready),
        .s_axis_iarg_109_aclk(s_axis_iarg_109_aclk),
        .s_axis_iarg_109_aresetn(s_axis_iarg_109_aresetn),
        .s_axis_iarg_109_tlast(s_axis_iarg_109_tlast),
        .s_axis_iarg_109_tvalid(s_axis_iarg_109_tvalid),
        .s_axis_iarg_109_tkeep(s_axis_iarg_109_tkeep),
        .s_axis_iarg_109_tstrb(s_axis_iarg_109_tstrb),
        .s_axis_iarg_109_tdata(s_axis_iarg_109_tdata),
        .s_axis_iarg_109_tready(s_axis_iarg_109_tready),
        .ap_axis_iarg_109_tlast(ap_axis_iarg_109_tlast),
        .ap_axis_iarg_109_tvalid(ap_axis_iarg_109_tvalid),
        .ap_axis_iarg_109_tkeep(ap_axis_iarg_109_tkeep),
        .ap_axis_iarg_109_tstrb(ap_axis_iarg_109_tstrb),
        .ap_axis_iarg_109_tdata(ap_axis_iarg_109_tdata),
        .ap_axis_iarg_109_tready(ap_axis_iarg_109_tready),
        .s_axis_iarg_110_aclk(s_axis_iarg_110_aclk),
        .s_axis_iarg_110_aresetn(s_axis_iarg_110_aresetn),
        .s_axis_iarg_110_tlast(s_axis_iarg_110_tlast),
        .s_axis_iarg_110_tvalid(s_axis_iarg_110_tvalid),
        .s_axis_iarg_110_tkeep(s_axis_iarg_110_tkeep),
        .s_axis_iarg_110_tstrb(s_axis_iarg_110_tstrb),
        .s_axis_iarg_110_tdata(s_axis_iarg_110_tdata),
        .s_axis_iarg_110_tready(s_axis_iarg_110_tready),
        .ap_axis_iarg_110_tlast(ap_axis_iarg_110_tlast),
        .ap_axis_iarg_110_tvalid(ap_axis_iarg_110_tvalid),
        .ap_axis_iarg_110_tkeep(ap_axis_iarg_110_tkeep),
        .ap_axis_iarg_110_tstrb(ap_axis_iarg_110_tstrb),
        .ap_axis_iarg_110_tdata(ap_axis_iarg_110_tdata),
        .ap_axis_iarg_110_tready(ap_axis_iarg_110_tready),
        .s_axis_iarg_111_aclk(s_axis_iarg_111_aclk),
        .s_axis_iarg_111_aresetn(s_axis_iarg_111_aresetn),
        .s_axis_iarg_111_tlast(s_axis_iarg_111_tlast),
        .s_axis_iarg_111_tvalid(s_axis_iarg_111_tvalid),
        .s_axis_iarg_111_tkeep(s_axis_iarg_111_tkeep),
        .s_axis_iarg_111_tstrb(s_axis_iarg_111_tstrb),
        .s_axis_iarg_111_tdata(s_axis_iarg_111_tdata),
        .s_axis_iarg_111_tready(s_axis_iarg_111_tready),
        .ap_axis_iarg_111_tlast(ap_axis_iarg_111_tlast),
        .ap_axis_iarg_111_tvalid(ap_axis_iarg_111_tvalid),
        .ap_axis_iarg_111_tkeep(ap_axis_iarg_111_tkeep),
        .ap_axis_iarg_111_tstrb(ap_axis_iarg_111_tstrb),
        .ap_axis_iarg_111_tdata(ap_axis_iarg_111_tdata),
        .ap_axis_iarg_111_tready(ap_axis_iarg_111_tready),
        .s_axis_iarg_112_aclk(s_axis_iarg_112_aclk),
        .s_axis_iarg_112_aresetn(s_axis_iarg_112_aresetn),
        .s_axis_iarg_112_tlast(s_axis_iarg_112_tlast),
        .s_axis_iarg_112_tvalid(s_axis_iarg_112_tvalid),
        .s_axis_iarg_112_tkeep(s_axis_iarg_112_tkeep),
        .s_axis_iarg_112_tstrb(s_axis_iarg_112_tstrb),
        .s_axis_iarg_112_tdata(s_axis_iarg_112_tdata),
        .s_axis_iarg_112_tready(s_axis_iarg_112_tready),
        .ap_axis_iarg_112_tlast(ap_axis_iarg_112_tlast),
        .ap_axis_iarg_112_tvalid(ap_axis_iarg_112_tvalid),
        .ap_axis_iarg_112_tkeep(ap_axis_iarg_112_tkeep),
        .ap_axis_iarg_112_tstrb(ap_axis_iarg_112_tstrb),
        .ap_axis_iarg_112_tdata(ap_axis_iarg_112_tdata),
        .ap_axis_iarg_112_tready(ap_axis_iarg_112_tready),
        .s_axis_iarg_113_aclk(s_axis_iarg_113_aclk),
        .s_axis_iarg_113_aresetn(s_axis_iarg_113_aresetn),
        .s_axis_iarg_113_tlast(s_axis_iarg_113_tlast),
        .s_axis_iarg_113_tvalid(s_axis_iarg_113_tvalid),
        .s_axis_iarg_113_tkeep(s_axis_iarg_113_tkeep),
        .s_axis_iarg_113_tstrb(s_axis_iarg_113_tstrb),
        .s_axis_iarg_113_tdata(s_axis_iarg_113_tdata),
        .s_axis_iarg_113_tready(s_axis_iarg_113_tready),
        .ap_axis_iarg_113_tlast(ap_axis_iarg_113_tlast),
        .ap_axis_iarg_113_tvalid(ap_axis_iarg_113_tvalid),
        .ap_axis_iarg_113_tkeep(ap_axis_iarg_113_tkeep),
        .ap_axis_iarg_113_tstrb(ap_axis_iarg_113_tstrb),
        .ap_axis_iarg_113_tdata(ap_axis_iarg_113_tdata),
        .ap_axis_iarg_113_tready(ap_axis_iarg_113_tready),
        .s_axis_iarg_114_aclk(s_axis_iarg_114_aclk),
        .s_axis_iarg_114_aresetn(s_axis_iarg_114_aresetn),
        .s_axis_iarg_114_tlast(s_axis_iarg_114_tlast),
        .s_axis_iarg_114_tvalid(s_axis_iarg_114_tvalid),
        .s_axis_iarg_114_tkeep(s_axis_iarg_114_tkeep),
        .s_axis_iarg_114_tstrb(s_axis_iarg_114_tstrb),
        .s_axis_iarg_114_tdata(s_axis_iarg_114_tdata),
        .s_axis_iarg_114_tready(s_axis_iarg_114_tready),
        .ap_axis_iarg_114_tlast(ap_axis_iarg_114_tlast),
        .ap_axis_iarg_114_tvalid(ap_axis_iarg_114_tvalid),
        .ap_axis_iarg_114_tkeep(ap_axis_iarg_114_tkeep),
        .ap_axis_iarg_114_tstrb(ap_axis_iarg_114_tstrb),
        .ap_axis_iarg_114_tdata(ap_axis_iarg_114_tdata),
        .ap_axis_iarg_114_tready(ap_axis_iarg_114_tready),
        .s_axis_iarg_115_aclk(s_axis_iarg_115_aclk),
        .s_axis_iarg_115_aresetn(s_axis_iarg_115_aresetn),
        .s_axis_iarg_115_tlast(s_axis_iarg_115_tlast),
        .s_axis_iarg_115_tvalid(s_axis_iarg_115_tvalid),
        .s_axis_iarg_115_tkeep(s_axis_iarg_115_tkeep),
        .s_axis_iarg_115_tstrb(s_axis_iarg_115_tstrb),
        .s_axis_iarg_115_tdata(s_axis_iarg_115_tdata),
        .s_axis_iarg_115_tready(s_axis_iarg_115_tready),
        .ap_axis_iarg_115_tlast(ap_axis_iarg_115_tlast),
        .ap_axis_iarg_115_tvalid(ap_axis_iarg_115_tvalid),
        .ap_axis_iarg_115_tkeep(ap_axis_iarg_115_tkeep),
        .ap_axis_iarg_115_tstrb(ap_axis_iarg_115_tstrb),
        .ap_axis_iarg_115_tdata(ap_axis_iarg_115_tdata),
        .ap_axis_iarg_115_tready(ap_axis_iarg_115_tready),
        .s_axis_iarg_116_aclk(s_axis_iarg_116_aclk),
        .s_axis_iarg_116_aresetn(s_axis_iarg_116_aresetn),
        .s_axis_iarg_116_tlast(s_axis_iarg_116_tlast),
        .s_axis_iarg_116_tvalid(s_axis_iarg_116_tvalid),
        .s_axis_iarg_116_tkeep(s_axis_iarg_116_tkeep),
        .s_axis_iarg_116_tstrb(s_axis_iarg_116_tstrb),
        .s_axis_iarg_116_tdata(s_axis_iarg_116_tdata),
        .s_axis_iarg_116_tready(s_axis_iarg_116_tready),
        .ap_axis_iarg_116_tlast(ap_axis_iarg_116_tlast),
        .ap_axis_iarg_116_tvalid(ap_axis_iarg_116_tvalid),
        .ap_axis_iarg_116_tkeep(ap_axis_iarg_116_tkeep),
        .ap_axis_iarg_116_tstrb(ap_axis_iarg_116_tstrb),
        .ap_axis_iarg_116_tdata(ap_axis_iarg_116_tdata),
        .ap_axis_iarg_116_tready(ap_axis_iarg_116_tready),
        .s_axis_iarg_117_aclk(s_axis_iarg_117_aclk),
        .s_axis_iarg_117_aresetn(s_axis_iarg_117_aresetn),
        .s_axis_iarg_117_tlast(s_axis_iarg_117_tlast),
        .s_axis_iarg_117_tvalid(s_axis_iarg_117_tvalid),
        .s_axis_iarg_117_tkeep(s_axis_iarg_117_tkeep),
        .s_axis_iarg_117_tstrb(s_axis_iarg_117_tstrb),
        .s_axis_iarg_117_tdata(s_axis_iarg_117_tdata),
        .s_axis_iarg_117_tready(s_axis_iarg_117_tready),
        .ap_axis_iarg_117_tlast(ap_axis_iarg_117_tlast),
        .ap_axis_iarg_117_tvalid(ap_axis_iarg_117_tvalid),
        .ap_axis_iarg_117_tkeep(ap_axis_iarg_117_tkeep),
        .ap_axis_iarg_117_tstrb(ap_axis_iarg_117_tstrb),
        .ap_axis_iarg_117_tdata(ap_axis_iarg_117_tdata),
        .ap_axis_iarg_117_tready(ap_axis_iarg_117_tready),
        .s_axis_iarg_118_aclk(s_axis_iarg_118_aclk),
        .s_axis_iarg_118_aresetn(s_axis_iarg_118_aresetn),
        .s_axis_iarg_118_tlast(s_axis_iarg_118_tlast),
        .s_axis_iarg_118_tvalid(s_axis_iarg_118_tvalid),
        .s_axis_iarg_118_tkeep(s_axis_iarg_118_tkeep),
        .s_axis_iarg_118_tstrb(s_axis_iarg_118_tstrb),
        .s_axis_iarg_118_tdata(s_axis_iarg_118_tdata),
        .s_axis_iarg_118_tready(s_axis_iarg_118_tready),
        .ap_axis_iarg_118_tlast(ap_axis_iarg_118_tlast),
        .ap_axis_iarg_118_tvalid(ap_axis_iarg_118_tvalid),
        .ap_axis_iarg_118_tkeep(ap_axis_iarg_118_tkeep),
        .ap_axis_iarg_118_tstrb(ap_axis_iarg_118_tstrb),
        .ap_axis_iarg_118_tdata(ap_axis_iarg_118_tdata),
        .ap_axis_iarg_118_tready(ap_axis_iarg_118_tready),
        .s_axis_iarg_119_aclk(s_axis_iarg_119_aclk),
        .s_axis_iarg_119_aresetn(s_axis_iarg_119_aresetn),
        .s_axis_iarg_119_tlast(s_axis_iarg_119_tlast),
        .s_axis_iarg_119_tvalid(s_axis_iarg_119_tvalid),
        .s_axis_iarg_119_tkeep(s_axis_iarg_119_tkeep),
        .s_axis_iarg_119_tstrb(s_axis_iarg_119_tstrb),
        .s_axis_iarg_119_tdata(s_axis_iarg_119_tdata),
        .s_axis_iarg_119_tready(s_axis_iarg_119_tready),
        .ap_axis_iarg_119_tlast(ap_axis_iarg_119_tlast),
        .ap_axis_iarg_119_tvalid(ap_axis_iarg_119_tvalid),
        .ap_axis_iarg_119_tkeep(ap_axis_iarg_119_tkeep),
        .ap_axis_iarg_119_tstrb(ap_axis_iarg_119_tstrb),
        .ap_axis_iarg_119_tdata(ap_axis_iarg_119_tdata),
        .ap_axis_iarg_119_tready(ap_axis_iarg_119_tready),
        .s_axis_iarg_120_aclk(s_axis_iarg_120_aclk),
        .s_axis_iarg_120_aresetn(s_axis_iarg_120_aresetn),
        .s_axis_iarg_120_tlast(s_axis_iarg_120_tlast),
        .s_axis_iarg_120_tvalid(s_axis_iarg_120_tvalid),
        .s_axis_iarg_120_tkeep(s_axis_iarg_120_tkeep),
        .s_axis_iarg_120_tstrb(s_axis_iarg_120_tstrb),
        .s_axis_iarg_120_tdata(s_axis_iarg_120_tdata),
        .s_axis_iarg_120_tready(s_axis_iarg_120_tready),
        .ap_axis_iarg_120_tlast(ap_axis_iarg_120_tlast),
        .ap_axis_iarg_120_tvalid(ap_axis_iarg_120_tvalid),
        .ap_axis_iarg_120_tkeep(ap_axis_iarg_120_tkeep),
        .ap_axis_iarg_120_tstrb(ap_axis_iarg_120_tstrb),
        .ap_axis_iarg_120_tdata(ap_axis_iarg_120_tdata),
        .ap_axis_iarg_120_tready(ap_axis_iarg_120_tready),
        .s_axis_iarg_121_aclk(s_axis_iarg_121_aclk),
        .s_axis_iarg_121_aresetn(s_axis_iarg_121_aresetn),
        .s_axis_iarg_121_tlast(s_axis_iarg_121_tlast),
        .s_axis_iarg_121_tvalid(s_axis_iarg_121_tvalid),
        .s_axis_iarg_121_tkeep(s_axis_iarg_121_tkeep),
        .s_axis_iarg_121_tstrb(s_axis_iarg_121_tstrb),
        .s_axis_iarg_121_tdata(s_axis_iarg_121_tdata),
        .s_axis_iarg_121_tready(s_axis_iarg_121_tready),
        .ap_axis_iarg_121_tlast(ap_axis_iarg_121_tlast),
        .ap_axis_iarg_121_tvalid(ap_axis_iarg_121_tvalid),
        .ap_axis_iarg_121_tkeep(ap_axis_iarg_121_tkeep),
        .ap_axis_iarg_121_tstrb(ap_axis_iarg_121_tstrb),
        .ap_axis_iarg_121_tdata(ap_axis_iarg_121_tdata),
        .ap_axis_iarg_121_tready(ap_axis_iarg_121_tready),
        .s_axis_iarg_122_aclk(s_axis_iarg_122_aclk),
        .s_axis_iarg_122_aresetn(s_axis_iarg_122_aresetn),
        .s_axis_iarg_122_tlast(s_axis_iarg_122_tlast),
        .s_axis_iarg_122_tvalid(s_axis_iarg_122_tvalid),
        .s_axis_iarg_122_tkeep(s_axis_iarg_122_tkeep),
        .s_axis_iarg_122_tstrb(s_axis_iarg_122_tstrb),
        .s_axis_iarg_122_tdata(s_axis_iarg_122_tdata),
        .s_axis_iarg_122_tready(s_axis_iarg_122_tready),
        .ap_axis_iarg_122_tlast(ap_axis_iarg_122_tlast),
        .ap_axis_iarg_122_tvalid(ap_axis_iarg_122_tvalid),
        .ap_axis_iarg_122_tkeep(ap_axis_iarg_122_tkeep),
        .ap_axis_iarg_122_tstrb(ap_axis_iarg_122_tstrb),
        .ap_axis_iarg_122_tdata(ap_axis_iarg_122_tdata),
        .ap_axis_iarg_122_tready(ap_axis_iarg_122_tready),
        .s_axis_iarg_123_aclk(s_axis_iarg_123_aclk),
        .s_axis_iarg_123_aresetn(s_axis_iarg_123_aresetn),
        .s_axis_iarg_123_tlast(s_axis_iarg_123_tlast),
        .s_axis_iarg_123_tvalid(s_axis_iarg_123_tvalid),
        .s_axis_iarg_123_tkeep(s_axis_iarg_123_tkeep),
        .s_axis_iarg_123_tstrb(s_axis_iarg_123_tstrb),
        .s_axis_iarg_123_tdata(s_axis_iarg_123_tdata),
        .s_axis_iarg_123_tready(s_axis_iarg_123_tready),
        .ap_axis_iarg_123_tlast(ap_axis_iarg_123_tlast),
        .ap_axis_iarg_123_tvalid(ap_axis_iarg_123_tvalid),
        .ap_axis_iarg_123_tkeep(ap_axis_iarg_123_tkeep),
        .ap_axis_iarg_123_tstrb(ap_axis_iarg_123_tstrb),
        .ap_axis_iarg_123_tdata(ap_axis_iarg_123_tdata),
        .ap_axis_iarg_123_tready(ap_axis_iarg_123_tready),
        .s_axis_iarg_124_aclk(s_axis_iarg_124_aclk),
        .s_axis_iarg_124_aresetn(s_axis_iarg_124_aresetn),
        .s_axis_iarg_124_tlast(s_axis_iarg_124_tlast),
        .s_axis_iarg_124_tvalid(s_axis_iarg_124_tvalid),
        .s_axis_iarg_124_tkeep(s_axis_iarg_124_tkeep),
        .s_axis_iarg_124_tstrb(s_axis_iarg_124_tstrb),
        .s_axis_iarg_124_tdata(s_axis_iarg_124_tdata),
        .s_axis_iarg_124_tready(s_axis_iarg_124_tready),
        .ap_axis_iarg_124_tlast(ap_axis_iarg_124_tlast),
        .ap_axis_iarg_124_tvalid(ap_axis_iarg_124_tvalid),
        .ap_axis_iarg_124_tkeep(ap_axis_iarg_124_tkeep),
        .ap_axis_iarg_124_tstrb(ap_axis_iarg_124_tstrb),
        .ap_axis_iarg_124_tdata(ap_axis_iarg_124_tdata),
        .ap_axis_iarg_124_tready(ap_axis_iarg_124_tready),
        .s_axis_iarg_125_aclk(s_axis_iarg_125_aclk),
        .s_axis_iarg_125_aresetn(s_axis_iarg_125_aresetn),
        .s_axis_iarg_125_tlast(s_axis_iarg_125_tlast),
        .s_axis_iarg_125_tvalid(s_axis_iarg_125_tvalid),
        .s_axis_iarg_125_tkeep(s_axis_iarg_125_tkeep),
        .s_axis_iarg_125_tstrb(s_axis_iarg_125_tstrb),
        .s_axis_iarg_125_tdata(s_axis_iarg_125_tdata),
        .s_axis_iarg_125_tready(s_axis_iarg_125_tready),
        .ap_axis_iarg_125_tlast(ap_axis_iarg_125_tlast),
        .ap_axis_iarg_125_tvalid(ap_axis_iarg_125_tvalid),
        .ap_axis_iarg_125_tkeep(ap_axis_iarg_125_tkeep),
        .ap_axis_iarg_125_tstrb(ap_axis_iarg_125_tstrb),
        .ap_axis_iarg_125_tdata(ap_axis_iarg_125_tdata),
        .ap_axis_iarg_125_tready(ap_axis_iarg_125_tready),
        .s_axis_iarg_126_aclk(s_axis_iarg_126_aclk),
        .s_axis_iarg_126_aresetn(s_axis_iarg_126_aresetn),
        .s_axis_iarg_126_tlast(s_axis_iarg_126_tlast),
        .s_axis_iarg_126_tvalid(s_axis_iarg_126_tvalid),
        .s_axis_iarg_126_tkeep(s_axis_iarg_126_tkeep),
        .s_axis_iarg_126_tstrb(s_axis_iarg_126_tstrb),
        .s_axis_iarg_126_tdata(s_axis_iarg_126_tdata),
        .s_axis_iarg_126_tready(s_axis_iarg_126_tready),
        .ap_axis_iarg_126_tlast(ap_axis_iarg_126_tlast),
        .ap_axis_iarg_126_tvalid(ap_axis_iarg_126_tvalid),
        .ap_axis_iarg_126_tkeep(ap_axis_iarg_126_tkeep),
        .ap_axis_iarg_126_tstrb(ap_axis_iarg_126_tstrb),
        .ap_axis_iarg_126_tdata(ap_axis_iarg_126_tdata),
        .ap_axis_iarg_126_tready(ap_axis_iarg_126_tready),
        .s_axis_iarg_127_aclk(s_axis_iarg_127_aclk),
        .s_axis_iarg_127_aresetn(s_axis_iarg_127_aresetn),
        .s_axis_iarg_127_tlast(s_axis_iarg_127_tlast),
        .s_axis_iarg_127_tvalid(s_axis_iarg_127_tvalid),
        .s_axis_iarg_127_tkeep(s_axis_iarg_127_tkeep),
        .s_axis_iarg_127_tstrb(s_axis_iarg_127_tstrb),
        .s_axis_iarg_127_tdata(s_axis_iarg_127_tdata),
        .s_axis_iarg_127_tready(s_axis_iarg_127_tready),
        .ap_axis_iarg_127_tlast(ap_axis_iarg_127_tlast),
        .ap_axis_iarg_127_tvalid(ap_axis_iarg_127_tvalid),
        .ap_axis_iarg_127_tkeep(ap_axis_iarg_127_tkeep),
        .ap_axis_iarg_127_tstrb(ap_axis_iarg_127_tstrb),
        .ap_axis_iarg_127_tdata(ap_axis_iarg_127_tdata),
        .ap_axis_iarg_127_tready(ap_axis_iarg_127_tready)
    );
        
    out_axis_args #(
        .C_NUM_OUTPUT_AXISs(C_NUM_OUTPUT_AXISs),
        .M_AXIS_OARG_0_WIDTH(M_AXIS_OARG_0_WIDTH),
        .M_AXIS_OARG_1_WIDTH(M_AXIS_OARG_1_WIDTH),
        .M_AXIS_OARG_2_WIDTH(M_AXIS_OARG_2_WIDTH),
        .M_AXIS_OARG_3_WIDTH(M_AXIS_OARG_3_WIDTH),
        .M_AXIS_OARG_4_WIDTH(M_AXIS_OARG_4_WIDTH),
        .M_AXIS_OARG_5_WIDTH(M_AXIS_OARG_5_WIDTH),
        .M_AXIS_OARG_6_WIDTH(M_AXIS_OARG_6_WIDTH),
        .M_AXIS_OARG_7_WIDTH(M_AXIS_OARG_7_WIDTH),
        .M_AXIS_OARG_8_WIDTH(M_AXIS_OARG_8_WIDTH),
        .M_AXIS_OARG_9_WIDTH(M_AXIS_OARG_9_WIDTH),
        .M_AXIS_OARG_10_WIDTH(M_AXIS_OARG_10_WIDTH),
        .M_AXIS_OARG_11_WIDTH(M_AXIS_OARG_11_WIDTH),
        .M_AXIS_OARG_12_WIDTH(M_AXIS_OARG_12_WIDTH),
        .M_AXIS_OARG_13_WIDTH(M_AXIS_OARG_13_WIDTH),
        .M_AXIS_OARG_14_WIDTH(M_AXIS_OARG_14_WIDTH),
        .M_AXIS_OARG_15_WIDTH(M_AXIS_OARG_15_WIDTH),
        .M_AXIS_OARG_16_WIDTH(M_AXIS_OARG_16_WIDTH),
        .M_AXIS_OARG_17_WIDTH(M_AXIS_OARG_17_WIDTH),
        .M_AXIS_OARG_18_WIDTH(M_AXIS_OARG_18_WIDTH),
        .M_AXIS_OARG_19_WIDTH(M_AXIS_OARG_19_WIDTH),
        .M_AXIS_OARG_20_WIDTH(M_AXIS_OARG_20_WIDTH),
        .M_AXIS_OARG_21_WIDTH(M_AXIS_OARG_21_WIDTH),
        .M_AXIS_OARG_22_WIDTH(M_AXIS_OARG_22_WIDTH),
        .M_AXIS_OARG_23_WIDTH(M_AXIS_OARG_23_WIDTH),
        .M_AXIS_OARG_24_WIDTH(M_AXIS_OARG_24_WIDTH),
        .M_AXIS_OARG_25_WIDTH(M_AXIS_OARG_25_WIDTH),
        .M_AXIS_OARG_26_WIDTH(M_AXIS_OARG_26_WIDTH),
        .M_AXIS_OARG_27_WIDTH(M_AXIS_OARG_27_WIDTH),
        .M_AXIS_OARG_28_WIDTH(M_AXIS_OARG_28_WIDTH),
        .M_AXIS_OARG_29_WIDTH(M_AXIS_OARG_29_WIDTH),
        .M_AXIS_OARG_30_WIDTH(M_AXIS_OARG_30_WIDTH),
        .M_AXIS_OARG_31_WIDTH(M_AXIS_OARG_31_WIDTH),
        .M_AXIS_OARG_32_WIDTH(M_AXIS_OARG_32_WIDTH),
        .M_AXIS_OARG_33_WIDTH(M_AXIS_OARG_33_WIDTH),
        .M_AXIS_OARG_34_WIDTH(M_AXIS_OARG_34_WIDTH),
        .M_AXIS_OARG_35_WIDTH(M_AXIS_OARG_35_WIDTH),
        .M_AXIS_OARG_36_WIDTH(M_AXIS_OARG_36_WIDTH),
        .M_AXIS_OARG_37_WIDTH(M_AXIS_OARG_37_WIDTH),
        .M_AXIS_OARG_38_WIDTH(M_AXIS_OARG_38_WIDTH),
        .M_AXIS_OARG_39_WIDTH(M_AXIS_OARG_39_WIDTH),
        .M_AXIS_OARG_40_WIDTH(M_AXIS_OARG_40_WIDTH),
        .M_AXIS_OARG_41_WIDTH(M_AXIS_OARG_41_WIDTH),
        .M_AXIS_OARG_42_WIDTH(M_AXIS_OARG_42_WIDTH),
        .M_AXIS_OARG_43_WIDTH(M_AXIS_OARG_43_WIDTH),
        .M_AXIS_OARG_44_WIDTH(M_AXIS_OARG_44_WIDTH),
        .M_AXIS_OARG_45_WIDTH(M_AXIS_OARG_45_WIDTH),
        .M_AXIS_OARG_46_WIDTH(M_AXIS_OARG_46_WIDTH),
        .M_AXIS_OARG_47_WIDTH(M_AXIS_OARG_47_WIDTH),
        .M_AXIS_OARG_48_WIDTH(M_AXIS_OARG_48_WIDTH),
        .M_AXIS_OARG_49_WIDTH(M_AXIS_OARG_49_WIDTH),
        .M_AXIS_OARG_50_WIDTH(M_AXIS_OARG_50_WIDTH),
        .M_AXIS_OARG_51_WIDTH(M_AXIS_OARG_51_WIDTH),
        .M_AXIS_OARG_52_WIDTH(M_AXIS_OARG_52_WIDTH),
        .M_AXIS_OARG_53_WIDTH(M_AXIS_OARG_53_WIDTH),
        .M_AXIS_OARG_54_WIDTH(M_AXIS_OARG_54_WIDTH),
        .M_AXIS_OARG_55_WIDTH(M_AXIS_OARG_55_WIDTH),
        .M_AXIS_OARG_56_WIDTH(M_AXIS_OARG_56_WIDTH),
        .M_AXIS_OARG_57_WIDTH(M_AXIS_OARG_57_WIDTH),
        .M_AXIS_OARG_58_WIDTH(M_AXIS_OARG_58_WIDTH),
        .M_AXIS_OARG_59_WIDTH(M_AXIS_OARG_59_WIDTH),
        .M_AXIS_OARG_60_WIDTH(M_AXIS_OARG_60_WIDTH),
        .M_AXIS_OARG_61_WIDTH(M_AXIS_OARG_61_WIDTH),
        .M_AXIS_OARG_62_WIDTH(M_AXIS_OARG_62_WIDTH),
        .M_AXIS_OARG_63_WIDTH(M_AXIS_OARG_63_WIDTH),
        .M_AXIS_OARG_64_WIDTH(M_AXIS_OARG_64_WIDTH),
        .M_AXIS_OARG_65_WIDTH(M_AXIS_OARG_65_WIDTH),
        .M_AXIS_OARG_66_WIDTH(M_AXIS_OARG_66_WIDTH),
        .M_AXIS_OARG_67_WIDTH(M_AXIS_OARG_67_WIDTH),
        .M_AXIS_OARG_68_WIDTH(M_AXIS_OARG_68_WIDTH),
        .M_AXIS_OARG_69_WIDTH(M_AXIS_OARG_69_WIDTH),
        .M_AXIS_OARG_70_WIDTH(M_AXIS_OARG_70_WIDTH),
        .M_AXIS_OARG_71_WIDTH(M_AXIS_OARG_71_WIDTH),
        .M_AXIS_OARG_72_WIDTH(M_AXIS_OARG_72_WIDTH),
        .M_AXIS_OARG_73_WIDTH(M_AXIS_OARG_73_WIDTH),
        .M_AXIS_OARG_74_WIDTH(M_AXIS_OARG_74_WIDTH),
        .M_AXIS_OARG_75_WIDTH(M_AXIS_OARG_75_WIDTH),
        .M_AXIS_OARG_76_WIDTH(M_AXIS_OARG_76_WIDTH),
        .M_AXIS_OARG_77_WIDTH(M_AXIS_OARG_77_WIDTH),
        .M_AXIS_OARG_78_WIDTH(M_AXIS_OARG_78_WIDTH),
        .M_AXIS_OARG_79_WIDTH(M_AXIS_OARG_79_WIDTH),
        .M_AXIS_OARG_80_WIDTH(M_AXIS_OARG_80_WIDTH),
        .M_AXIS_OARG_81_WIDTH(M_AXIS_OARG_81_WIDTH),
        .M_AXIS_OARG_82_WIDTH(M_AXIS_OARG_82_WIDTH),
        .M_AXIS_OARG_83_WIDTH(M_AXIS_OARG_83_WIDTH),
        .M_AXIS_OARG_84_WIDTH(M_AXIS_OARG_84_WIDTH),
        .M_AXIS_OARG_85_WIDTH(M_AXIS_OARG_85_WIDTH),
        .M_AXIS_OARG_86_WIDTH(M_AXIS_OARG_86_WIDTH),
        .M_AXIS_OARG_87_WIDTH(M_AXIS_OARG_87_WIDTH),
        .M_AXIS_OARG_88_WIDTH(M_AXIS_OARG_88_WIDTH),
        .M_AXIS_OARG_89_WIDTH(M_AXIS_OARG_89_WIDTH),
        .M_AXIS_OARG_90_WIDTH(M_AXIS_OARG_90_WIDTH),
        .M_AXIS_OARG_91_WIDTH(M_AXIS_OARG_91_WIDTH),
        .M_AXIS_OARG_92_WIDTH(M_AXIS_OARG_92_WIDTH),
        .M_AXIS_OARG_93_WIDTH(M_AXIS_OARG_93_WIDTH),
        .M_AXIS_OARG_94_WIDTH(M_AXIS_OARG_94_WIDTH),
        .M_AXIS_OARG_95_WIDTH(M_AXIS_OARG_95_WIDTH),
        .M_AXIS_OARG_96_WIDTH(M_AXIS_OARG_96_WIDTH),
        .M_AXIS_OARG_97_WIDTH(M_AXIS_OARG_97_WIDTH),
        .M_AXIS_OARG_98_WIDTH(M_AXIS_OARG_98_WIDTH),
        .M_AXIS_OARG_99_WIDTH(M_AXIS_OARG_99_WIDTH),
        .M_AXIS_OARG_100_WIDTH(M_AXIS_OARG_100_WIDTH),
        .M_AXIS_OARG_101_WIDTH(M_AXIS_OARG_101_WIDTH),
        .M_AXIS_OARG_102_WIDTH(M_AXIS_OARG_102_WIDTH),
        .M_AXIS_OARG_103_WIDTH(M_AXIS_OARG_103_WIDTH),
        .M_AXIS_OARG_104_WIDTH(M_AXIS_OARG_104_WIDTH),
        .M_AXIS_OARG_105_WIDTH(M_AXIS_OARG_105_WIDTH),
        .M_AXIS_OARG_106_WIDTH(M_AXIS_OARG_106_WIDTH),
        .M_AXIS_OARG_107_WIDTH(M_AXIS_OARG_107_WIDTH),
        .M_AXIS_OARG_108_WIDTH(M_AXIS_OARG_108_WIDTH),
        .M_AXIS_OARG_109_WIDTH(M_AXIS_OARG_109_WIDTH),
        .M_AXIS_OARG_110_WIDTH(M_AXIS_OARG_110_WIDTH),
        .M_AXIS_OARG_111_WIDTH(M_AXIS_OARG_111_WIDTH),
        .M_AXIS_OARG_112_WIDTH(M_AXIS_OARG_112_WIDTH),
        .M_AXIS_OARG_113_WIDTH(M_AXIS_OARG_113_WIDTH),
        .M_AXIS_OARG_114_WIDTH(M_AXIS_OARG_114_WIDTH),
        .M_AXIS_OARG_115_WIDTH(M_AXIS_OARG_115_WIDTH),
        .M_AXIS_OARG_116_WIDTH(M_AXIS_OARG_116_WIDTH),
        .M_AXIS_OARG_117_WIDTH(M_AXIS_OARG_117_WIDTH),
        .M_AXIS_OARG_118_WIDTH(M_AXIS_OARG_118_WIDTH),
        .M_AXIS_OARG_119_WIDTH(M_AXIS_OARG_119_WIDTH),
        .M_AXIS_OARG_120_WIDTH(M_AXIS_OARG_120_WIDTH),
        .M_AXIS_OARG_121_WIDTH(M_AXIS_OARG_121_WIDTH),
        .M_AXIS_OARG_122_WIDTH(M_AXIS_OARG_122_WIDTH),
        .M_AXIS_OARG_123_WIDTH(M_AXIS_OARG_123_WIDTH),
        .M_AXIS_OARG_124_WIDTH(M_AXIS_OARG_124_WIDTH),
        .M_AXIS_OARG_125_WIDTH(M_AXIS_OARG_125_WIDTH),
        .M_AXIS_OARG_126_WIDTH(M_AXIS_OARG_126_WIDTH),
        .M_AXIS_OARG_127_WIDTH(M_AXIS_OARG_127_WIDTH),
        .M_AXIS_OARG_0_DEPTH(M_AXIS_OARG_0_DEPTH),
        .M_AXIS_OARG_1_DEPTH(M_AXIS_OARG_1_DEPTH),
        .M_AXIS_OARG_2_DEPTH(M_AXIS_OARG_2_DEPTH),
        .M_AXIS_OARG_3_DEPTH(M_AXIS_OARG_3_DEPTH),
        .M_AXIS_OARG_4_DEPTH(M_AXIS_OARG_4_DEPTH),
        .M_AXIS_OARG_5_DEPTH(M_AXIS_OARG_5_DEPTH),
        .M_AXIS_OARG_6_DEPTH(M_AXIS_OARG_6_DEPTH),
        .M_AXIS_OARG_7_DEPTH(M_AXIS_OARG_7_DEPTH),
        .M_AXIS_OARG_8_DEPTH(M_AXIS_OARG_8_DEPTH),
        .M_AXIS_OARG_9_DEPTH(M_AXIS_OARG_9_DEPTH),
        .M_AXIS_OARG_10_DEPTH(M_AXIS_OARG_10_DEPTH),
        .M_AXIS_OARG_11_DEPTH(M_AXIS_OARG_11_DEPTH),
        .M_AXIS_OARG_12_DEPTH(M_AXIS_OARG_12_DEPTH),
        .M_AXIS_OARG_13_DEPTH(M_AXIS_OARG_13_DEPTH),
        .M_AXIS_OARG_14_DEPTH(M_AXIS_OARG_14_DEPTH),
        .M_AXIS_OARG_15_DEPTH(M_AXIS_OARG_15_DEPTH),
        .M_AXIS_OARG_16_DEPTH(M_AXIS_OARG_16_DEPTH),
        .M_AXIS_OARG_17_DEPTH(M_AXIS_OARG_17_DEPTH),
        .M_AXIS_OARG_18_DEPTH(M_AXIS_OARG_18_DEPTH),
        .M_AXIS_OARG_19_DEPTH(M_AXIS_OARG_19_DEPTH),
        .M_AXIS_OARG_20_DEPTH(M_AXIS_OARG_20_DEPTH),
        .M_AXIS_OARG_21_DEPTH(M_AXIS_OARG_21_DEPTH),
        .M_AXIS_OARG_22_DEPTH(M_AXIS_OARG_22_DEPTH),
        .M_AXIS_OARG_23_DEPTH(M_AXIS_OARG_23_DEPTH),
        .M_AXIS_OARG_24_DEPTH(M_AXIS_OARG_24_DEPTH),
        .M_AXIS_OARG_25_DEPTH(M_AXIS_OARG_25_DEPTH),
        .M_AXIS_OARG_26_DEPTH(M_AXIS_OARG_26_DEPTH),
        .M_AXIS_OARG_27_DEPTH(M_AXIS_OARG_27_DEPTH),
        .M_AXIS_OARG_28_DEPTH(M_AXIS_OARG_28_DEPTH),
        .M_AXIS_OARG_29_DEPTH(M_AXIS_OARG_29_DEPTH),
        .M_AXIS_OARG_30_DEPTH(M_AXIS_OARG_30_DEPTH),
        .M_AXIS_OARG_31_DEPTH(M_AXIS_OARG_31_DEPTH),
        .M_AXIS_OARG_32_DEPTH(M_AXIS_OARG_32_DEPTH),
        .M_AXIS_OARG_33_DEPTH(M_AXIS_OARG_33_DEPTH),
        .M_AXIS_OARG_34_DEPTH(M_AXIS_OARG_34_DEPTH),
        .M_AXIS_OARG_35_DEPTH(M_AXIS_OARG_35_DEPTH),
        .M_AXIS_OARG_36_DEPTH(M_AXIS_OARG_36_DEPTH),
        .M_AXIS_OARG_37_DEPTH(M_AXIS_OARG_37_DEPTH),
        .M_AXIS_OARG_38_DEPTH(M_AXIS_OARG_38_DEPTH),
        .M_AXIS_OARG_39_DEPTH(M_AXIS_OARG_39_DEPTH),
        .M_AXIS_OARG_40_DEPTH(M_AXIS_OARG_40_DEPTH),
        .M_AXIS_OARG_41_DEPTH(M_AXIS_OARG_41_DEPTH),
        .M_AXIS_OARG_42_DEPTH(M_AXIS_OARG_42_DEPTH),
        .M_AXIS_OARG_43_DEPTH(M_AXIS_OARG_43_DEPTH),
        .M_AXIS_OARG_44_DEPTH(M_AXIS_OARG_44_DEPTH),
        .M_AXIS_OARG_45_DEPTH(M_AXIS_OARG_45_DEPTH),
        .M_AXIS_OARG_46_DEPTH(M_AXIS_OARG_46_DEPTH),
        .M_AXIS_OARG_47_DEPTH(M_AXIS_OARG_47_DEPTH),
        .M_AXIS_OARG_48_DEPTH(M_AXIS_OARG_48_DEPTH),
        .M_AXIS_OARG_49_DEPTH(M_AXIS_OARG_49_DEPTH),
        .M_AXIS_OARG_50_DEPTH(M_AXIS_OARG_50_DEPTH),
        .M_AXIS_OARG_51_DEPTH(M_AXIS_OARG_51_DEPTH),
        .M_AXIS_OARG_52_DEPTH(M_AXIS_OARG_52_DEPTH),
        .M_AXIS_OARG_53_DEPTH(M_AXIS_OARG_53_DEPTH),
        .M_AXIS_OARG_54_DEPTH(M_AXIS_OARG_54_DEPTH),
        .M_AXIS_OARG_55_DEPTH(M_AXIS_OARG_55_DEPTH),
        .M_AXIS_OARG_56_DEPTH(M_AXIS_OARG_56_DEPTH),
        .M_AXIS_OARG_57_DEPTH(M_AXIS_OARG_57_DEPTH),
        .M_AXIS_OARG_58_DEPTH(M_AXIS_OARG_58_DEPTH),
        .M_AXIS_OARG_59_DEPTH(M_AXIS_OARG_59_DEPTH),
        .M_AXIS_OARG_60_DEPTH(M_AXIS_OARG_60_DEPTH),
        .M_AXIS_OARG_61_DEPTH(M_AXIS_OARG_61_DEPTH),
        .M_AXIS_OARG_62_DEPTH(M_AXIS_OARG_62_DEPTH),
        .M_AXIS_OARG_63_DEPTH(M_AXIS_OARG_63_DEPTH),
        .M_AXIS_OARG_64_DEPTH(M_AXIS_OARG_64_DEPTH),
        .M_AXIS_OARG_65_DEPTH(M_AXIS_OARG_65_DEPTH),
        .M_AXIS_OARG_66_DEPTH(M_AXIS_OARG_66_DEPTH),
        .M_AXIS_OARG_67_DEPTH(M_AXIS_OARG_67_DEPTH),
        .M_AXIS_OARG_68_DEPTH(M_AXIS_OARG_68_DEPTH),
        .M_AXIS_OARG_69_DEPTH(M_AXIS_OARG_69_DEPTH),
        .M_AXIS_OARG_70_DEPTH(M_AXIS_OARG_70_DEPTH),
        .M_AXIS_OARG_71_DEPTH(M_AXIS_OARG_71_DEPTH),
        .M_AXIS_OARG_72_DEPTH(M_AXIS_OARG_72_DEPTH),
        .M_AXIS_OARG_73_DEPTH(M_AXIS_OARG_73_DEPTH),
        .M_AXIS_OARG_74_DEPTH(M_AXIS_OARG_74_DEPTH),
        .M_AXIS_OARG_75_DEPTH(M_AXIS_OARG_75_DEPTH),
        .M_AXIS_OARG_76_DEPTH(M_AXIS_OARG_76_DEPTH),
        .M_AXIS_OARG_77_DEPTH(M_AXIS_OARG_77_DEPTH),
        .M_AXIS_OARG_78_DEPTH(M_AXIS_OARG_78_DEPTH),
        .M_AXIS_OARG_79_DEPTH(M_AXIS_OARG_79_DEPTH),
        .M_AXIS_OARG_80_DEPTH(M_AXIS_OARG_80_DEPTH),
        .M_AXIS_OARG_81_DEPTH(M_AXIS_OARG_81_DEPTH),
        .M_AXIS_OARG_82_DEPTH(M_AXIS_OARG_82_DEPTH),
        .M_AXIS_OARG_83_DEPTH(M_AXIS_OARG_83_DEPTH),
        .M_AXIS_OARG_84_DEPTH(M_AXIS_OARG_84_DEPTH),
        .M_AXIS_OARG_85_DEPTH(M_AXIS_OARG_85_DEPTH),
        .M_AXIS_OARG_86_DEPTH(M_AXIS_OARG_86_DEPTH),
        .M_AXIS_OARG_87_DEPTH(M_AXIS_OARG_87_DEPTH),
        .M_AXIS_OARG_88_DEPTH(M_AXIS_OARG_88_DEPTH),
        .M_AXIS_OARG_89_DEPTH(M_AXIS_OARG_89_DEPTH),
        .M_AXIS_OARG_90_DEPTH(M_AXIS_OARG_90_DEPTH),
        .M_AXIS_OARG_91_DEPTH(M_AXIS_OARG_91_DEPTH),
        .M_AXIS_OARG_92_DEPTH(M_AXIS_OARG_92_DEPTH),
        .M_AXIS_OARG_93_DEPTH(M_AXIS_OARG_93_DEPTH),
        .M_AXIS_OARG_94_DEPTH(M_AXIS_OARG_94_DEPTH),
        .M_AXIS_OARG_95_DEPTH(M_AXIS_OARG_95_DEPTH),
        .M_AXIS_OARG_96_DEPTH(M_AXIS_OARG_96_DEPTH),
        .M_AXIS_OARG_97_DEPTH(M_AXIS_OARG_97_DEPTH),
        .M_AXIS_OARG_98_DEPTH(M_AXIS_OARG_98_DEPTH),
        .M_AXIS_OARG_99_DEPTH(M_AXIS_OARG_99_DEPTH),
        .M_AXIS_OARG_100_DEPTH(M_AXIS_OARG_100_DEPTH),
        .M_AXIS_OARG_101_DEPTH(M_AXIS_OARG_101_DEPTH),
        .M_AXIS_OARG_102_DEPTH(M_AXIS_OARG_102_DEPTH),
        .M_AXIS_OARG_103_DEPTH(M_AXIS_OARG_103_DEPTH),
        .M_AXIS_OARG_104_DEPTH(M_AXIS_OARG_104_DEPTH),
        .M_AXIS_OARG_105_DEPTH(M_AXIS_OARG_105_DEPTH),
        .M_AXIS_OARG_106_DEPTH(M_AXIS_OARG_106_DEPTH),
        .M_AXIS_OARG_107_DEPTH(M_AXIS_OARG_107_DEPTH),
        .M_AXIS_OARG_108_DEPTH(M_AXIS_OARG_108_DEPTH),
        .M_AXIS_OARG_109_DEPTH(M_AXIS_OARG_109_DEPTH),
        .M_AXIS_OARG_110_DEPTH(M_AXIS_OARG_110_DEPTH),
        .M_AXIS_OARG_111_DEPTH(M_AXIS_OARG_111_DEPTH),
        .M_AXIS_OARG_112_DEPTH(M_AXIS_OARG_112_DEPTH),
        .M_AXIS_OARG_113_DEPTH(M_AXIS_OARG_113_DEPTH),
        .M_AXIS_OARG_114_DEPTH(M_AXIS_OARG_114_DEPTH),
        .M_AXIS_OARG_115_DEPTH(M_AXIS_OARG_115_DEPTH),
        .M_AXIS_OARG_116_DEPTH(M_AXIS_OARG_116_DEPTH),
        .M_AXIS_OARG_117_DEPTH(M_AXIS_OARG_117_DEPTH),
        .M_AXIS_OARG_118_DEPTH(M_AXIS_OARG_118_DEPTH),
        .M_AXIS_OARG_119_DEPTH(M_AXIS_OARG_119_DEPTH),
        .M_AXIS_OARG_120_DEPTH(M_AXIS_OARG_120_DEPTH),
        .M_AXIS_OARG_121_DEPTH(M_AXIS_OARG_121_DEPTH),
        .M_AXIS_OARG_122_DEPTH(M_AXIS_OARG_122_DEPTH),
        .M_AXIS_OARG_123_DEPTH(M_AXIS_OARG_123_DEPTH),
        .M_AXIS_OARG_124_DEPTH(M_AXIS_OARG_124_DEPTH),
        .M_AXIS_OARG_125_DEPTH(M_AXIS_OARG_125_DEPTH),
        .M_AXIS_OARG_126_DEPTH(M_AXIS_OARG_126_DEPTH),
        .M_AXIS_OARG_127_DEPTH(M_AXIS_OARG_127_DEPTH),
        .M_AXIS_OARG_0_IS_ASYNC(M_AXIS_OARG_0_IS_ASYNC),
        .M_AXIS_OARG_1_IS_ASYNC(M_AXIS_OARG_1_IS_ASYNC),
        .M_AXIS_OARG_2_IS_ASYNC(M_AXIS_OARG_2_IS_ASYNC),
        .M_AXIS_OARG_3_IS_ASYNC(M_AXIS_OARG_3_IS_ASYNC),
        .M_AXIS_OARG_4_IS_ASYNC(M_AXIS_OARG_4_IS_ASYNC),
        .M_AXIS_OARG_5_IS_ASYNC(M_AXIS_OARG_5_IS_ASYNC),
        .M_AXIS_OARG_6_IS_ASYNC(M_AXIS_OARG_6_IS_ASYNC),
        .M_AXIS_OARG_7_IS_ASYNC(M_AXIS_OARG_7_IS_ASYNC),
        .M_AXIS_OARG_8_IS_ASYNC(M_AXIS_OARG_8_IS_ASYNC),
        .M_AXIS_OARG_9_IS_ASYNC(M_AXIS_OARG_9_IS_ASYNC),
        .M_AXIS_OARG_10_IS_ASYNC(M_AXIS_OARG_10_IS_ASYNC),
        .M_AXIS_OARG_11_IS_ASYNC(M_AXIS_OARG_11_IS_ASYNC),
        .M_AXIS_OARG_12_IS_ASYNC(M_AXIS_OARG_12_IS_ASYNC),
        .M_AXIS_OARG_13_IS_ASYNC(M_AXIS_OARG_13_IS_ASYNC),
        .M_AXIS_OARG_14_IS_ASYNC(M_AXIS_OARG_14_IS_ASYNC),
        .M_AXIS_OARG_15_IS_ASYNC(M_AXIS_OARG_15_IS_ASYNC),
        .M_AXIS_OARG_16_IS_ASYNC(M_AXIS_OARG_16_IS_ASYNC),
        .M_AXIS_OARG_17_IS_ASYNC(M_AXIS_OARG_17_IS_ASYNC),
        .M_AXIS_OARG_18_IS_ASYNC(M_AXIS_OARG_18_IS_ASYNC),
        .M_AXIS_OARG_19_IS_ASYNC(M_AXIS_OARG_19_IS_ASYNC),
        .M_AXIS_OARG_20_IS_ASYNC(M_AXIS_OARG_20_IS_ASYNC),
        .M_AXIS_OARG_21_IS_ASYNC(M_AXIS_OARG_21_IS_ASYNC),
        .M_AXIS_OARG_22_IS_ASYNC(M_AXIS_OARG_22_IS_ASYNC),
        .M_AXIS_OARG_23_IS_ASYNC(M_AXIS_OARG_23_IS_ASYNC),
        .M_AXIS_OARG_24_IS_ASYNC(M_AXIS_OARG_24_IS_ASYNC),
        .M_AXIS_OARG_25_IS_ASYNC(M_AXIS_OARG_25_IS_ASYNC),
        .M_AXIS_OARG_26_IS_ASYNC(M_AXIS_OARG_26_IS_ASYNC),
        .M_AXIS_OARG_27_IS_ASYNC(M_AXIS_OARG_27_IS_ASYNC),
        .M_AXIS_OARG_28_IS_ASYNC(M_AXIS_OARG_28_IS_ASYNC),
        .M_AXIS_OARG_29_IS_ASYNC(M_AXIS_OARG_29_IS_ASYNC),
        .M_AXIS_OARG_30_IS_ASYNC(M_AXIS_OARG_30_IS_ASYNC),
        .M_AXIS_OARG_31_IS_ASYNC(M_AXIS_OARG_31_IS_ASYNC),
        .M_AXIS_OARG_32_IS_ASYNC(M_AXIS_OARG_32_IS_ASYNC),
        .M_AXIS_OARG_33_IS_ASYNC(M_AXIS_OARG_33_IS_ASYNC),
        .M_AXIS_OARG_34_IS_ASYNC(M_AXIS_OARG_34_IS_ASYNC),
        .M_AXIS_OARG_35_IS_ASYNC(M_AXIS_OARG_35_IS_ASYNC),
        .M_AXIS_OARG_36_IS_ASYNC(M_AXIS_OARG_36_IS_ASYNC),
        .M_AXIS_OARG_37_IS_ASYNC(M_AXIS_OARG_37_IS_ASYNC),
        .M_AXIS_OARG_38_IS_ASYNC(M_AXIS_OARG_38_IS_ASYNC),
        .M_AXIS_OARG_39_IS_ASYNC(M_AXIS_OARG_39_IS_ASYNC),
        .M_AXIS_OARG_40_IS_ASYNC(M_AXIS_OARG_40_IS_ASYNC),
        .M_AXIS_OARG_41_IS_ASYNC(M_AXIS_OARG_41_IS_ASYNC),
        .M_AXIS_OARG_42_IS_ASYNC(M_AXIS_OARG_42_IS_ASYNC),
        .M_AXIS_OARG_43_IS_ASYNC(M_AXIS_OARG_43_IS_ASYNC),
        .M_AXIS_OARG_44_IS_ASYNC(M_AXIS_OARG_44_IS_ASYNC),
        .M_AXIS_OARG_45_IS_ASYNC(M_AXIS_OARG_45_IS_ASYNC),
        .M_AXIS_OARG_46_IS_ASYNC(M_AXIS_OARG_46_IS_ASYNC),
        .M_AXIS_OARG_47_IS_ASYNC(M_AXIS_OARG_47_IS_ASYNC),
        .M_AXIS_OARG_48_IS_ASYNC(M_AXIS_OARG_48_IS_ASYNC),
        .M_AXIS_OARG_49_IS_ASYNC(M_AXIS_OARG_49_IS_ASYNC),
        .M_AXIS_OARG_50_IS_ASYNC(M_AXIS_OARG_50_IS_ASYNC),
        .M_AXIS_OARG_51_IS_ASYNC(M_AXIS_OARG_51_IS_ASYNC),
        .M_AXIS_OARG_52_IS_ASYNC(M_AXIS_OARG_52_IS_ASYNC),
        .M_AXIS_OARG_53_IS_ASYNC(M_AXIS_OARG_53_IS_ASYNC),
        .M_AXIS_OARG_54_IS_ASYNC(M_AXIS_OARG_54_IS_ASYNC),
        .M_AXIS_OARG_55_IS_ASYNC(M_AXIS_OARG_55_IS_ASYNC),
        .M_AXIS_OARG_56_IS_ASYNC(M_AXIS_OARG_56_IS_ASYNC),
        .M_AXIS_OARG_57_IS_ASYNC(M_AXIS_OARG_57_IS_ASYNC),
        .M_AXIS_OARG_58_IS_ASYNC(M_AXIS_OARG_58_IS_ASYNC),
        .M_AXIS_OARG_59_IS_ASYNC(M_AXIS_OARG_59_IS_ASYNC),
        .M_AXIS_OARG_60_IS_ASYNC(M_AXIS_OARG_60_IS_ASYNC),
        .M_AXIS_OARG_61_IS_ASYNC(M_AXIS_OARG_61_IS_ASYNC),
        .M_AXIS_OARG_62_IS_ASYNC(M_AXIS_OARG_62_IS_ASYNC),
        .M_AXIS_OARG_63_IS_ASYNC(M_AXIS_OARG_63_IS_ASYNC),
        .M_AXIS_OARG_64_IS_ASYNC(M_AXIS_OARG_64_IS_ASYNC),
        .M_AXIS_OARG_65_IS_ASYNC(M_AXIS_OARG_65_IS_ASYNC),
        .M_AXIS_OARG_66_IS_ASYNC(M_AXIS_OARG_66_IS_ASYNC),
        .M_AXIS_OARG_67_IS_ASYNC(M_AXIS_OARG_67_IS_ASYNC),
        .M_AXIS_OARG_68_IS_ASYNC(M_AXIS_OARG_68_IS_ASYNC),
        .M_AXIS_OARG_69_IS_ASYNC(M_AXIS_OARG_69_IS_ASYNC),
        .M_AXIS_OARG_70_IS_ASYNC(M_AXIS_OARG_70_IS_ASYNC),
        .M_AXIS_OARG_71_IS_ASYNC(M_AXIS_OARG_71_IS_ASYNC),
        .M_AXIS_OARG_72_IS_ASYNC(M_AXIS_OARG_72_IS_ASYNC),
        .M_AXIS_OARG_73_IS_ASYNC(M_AXIS_OARG_73_IS_ASYNC),
        .M_AXIS_OARG_74_IS_ASYNC(M_AXIS_OARG_74_IS_ASYNC),
        .M_AXIS_OARG_75_IS_ASYNC(M_AXIS_OARG_75_IS_ASYNC),
        .M_AXIS_OARG_76_IS_ASYNC(M_AXIS_OARG_76_IS_ASYNC),
        .M_AXIS_OARG_77_IS_ASYNC(M_AXIS_OARG_77_IS_ASYNC),
        .M_AXIS_OARG_78_IS_ASYNC(M_AXIS_OARG_78_IS_ASYNC),
        .M_AXIS_OARG_79_IS_ASYNC(M_AXIS_OARG_79_IS_ASYNC),
        .M_AXIS_OARG_80_IS_ASYNC(M_AXIS_OARG_80_IS_ASYNC),
        .M_AXIS_OARG_81_IS_ASYNC(M_AXIS_OARG_81_IS_ASYNC),
        .M_AXIS_OARG_82_IS_ASYNC(M_AXIS_OARG_82_IS_ASYNC),
        .M_AXIS_OARG_83_IS_ASYNC(M_AXIS_OARG_83_IS_ASYNC),
        .M_AXIS_OARG_84_IS_ASYNC(M_AXIS_OARG_84_IS_ASYNC),
        .M_AXIS_OARG_85_IS_ASYNC(M_AXIS_OARG_85_IS_ASYNC),
        .M_AXIS_OARG_86_IS_ASYNC(M_AXIS_OARG_86_IS_ASYNC),
        .M_AXIS_OARG_87_IS_ASYNC(M_AXIS_OARG_87_IS_ASYNC),
        .M_AXIS_OARG_88_IS_ASYNC(M_AXIS_OARG_88_IS_ASYNC),
        .M_AXIS_OARG_89_IS_ASYNC(M_AXIS_OARG_89_IS_ASYNC),
        .M_AXIS_OARG_90_IS_ASYNC(M_AXIS_OARG_90_IS_ASYNC),
        .M_AXIS_OARG_91_IS_ASYNC(M_AXIS_OARG_91_IS_ASYNC),
        .M_AXIS_OARG_92_IS_ASYNC(M_AXIS_OARG_92_IS_ASYNC),
        .M_AXIS_OARG_93_IS_ASYNC(M_AXIS_OARG_93_IS_ASYNC),
        .M_AXIS_OARG_94_IS_ASYNC(M_AXIS_OARG_94_IS_ASYNC),
        .M_AXIS_OARG_95_IS_ASYNC(M_AXIS_OARG_95_IS_ASYNC),
        .M_AXIS_OARG_96_IS_ASYNC(M_AXIS_OARG_96_IS_ASYNC),
        .M_AXIS_OARG_97_IS_ASYNC(M_AXIS_OARG_97_IS_ASYNC),
        .M_AXIS_OARG_98_IS_ASYNC(M_AXIS_OARG_98_IS_ASYNC),
        .M_AXIS_OARG_99_IS_ASYNC(M_AXIS_OARG_99_IS_ASYNC),
        .M_AXIS_OARG_100_IS_ASYNC(M_AXIS_OARG_100_IS_ASYNC),
        .M_AXIS_OARG_101_IS_ASYNC(M_AXIS_OARG_101_IS_ASYNC),
        .M_AXIS_OARG_102_IS_ASYNC(M_AXIS_OARG_102_IS_ASYNC),
        .M_AXIS_OARG_103_IS_ASYNC(M_AXIS_OARG_103_IS_ASYNC),
        .M_AXIS_OARG_104_IS_ASYNC(M_AXIS_OARG_104_IS_ASYNC),
        .M_AXIS_OARG_105_IS_ASYNC(M_AXIS_OARG_105_IS_ASYNC),
        .M_AXIS_OARG_106_IS_ASYNC(M_AXIS_OARG_106_IS_ASYNC),
        .M_AXIS_OARG_107_IS_ASYNC(M_AXIS_OARG_107_IS_ASYNC),
        .M_AXIS_OARG_108_IS_ASYNC(M_AXIS_OARG_108_IS_ASYNC),
        .M_AXIS_OARG_109_IS_ASYNC(M_AXIS_OARG_109_IS_ASYNC),
        .M_AXIS_OARG_110_IS_ASYNC(M_AXIS_OARG_110_IS_ASYNC),
        .M_AXIS_OARG_111_IS_ASYNC(M_AXIS_OARG_111_IS_ASYNC),
        .M_AXIS_OARG_112_IS_ASYNC(M_AXIS_OARG_112_IS_ASYNC),
        .M_AXIS_OARG_113_IS_ASYNC(M_AXIS_OARG_113_IS_ASYNC),
        .M_AXIS_OARG_114_IS_ASYNC(M_AXIS_OARG_114_IS_ASYNC),
        .M_AXIS_OARG_115_IS_ASYNC(M_AXIS_OARG_115_IS_ASYNC),
        .M_AXIS_OARG_116_IS_ASYNC(M_AXIS_OARG_116_IS_ASYNC),
        .M_AXIS_OARG_117_IS_ASYNC(M_AXIS_OARG_117_IS_ASYNC),
        .M_AXIS_OARG_118_IS_ASYNC(M_AXIS_OARG_118_IS_ASYNC),
        .M_AXIS_OARG_119_IS_ASYNC(M_AXIS_OARG_119_IS_ASYNC),
        .M_AXIS_OARG_120_IS_ASYNC(M_AXIS_OARG_120_IS_ASYNC),
        .M_AXIS_OARG_121_IS_ASYNC(M_AXIS_OARG_121_IS_ASYNC),
        .M_AXIS_OARG_122_IS_ASYNC(M_AXIS_OARG_122_IS_ASYNC),
        .M_AXIS_OARG_123_IS_ASYNC(M_AXIS_OARG_123_IS_ASYNC),
        .M_AXIS_OARG_124_IS_ASYNC(M_AXIS_OARG_124_IS_ASYNC),
        .M_AXIS_OARG_125_IS_ASYNC(M_AXIS_OARG_125_IS_ASYNC),
        .M_AXIS_OARG_126_IS_ASYNC(M_AXIS_OARG_126_IS_ASYNC),
        .M_AXIS_OARG_127_IS_ASYNC(M_AXIS_OARG_127_IS_ASYNC),
        .M_AXIS_OARG_0_GEN_TLAST(M_AXIS_OARG_0_GEN_TLAST),
        .M_AXIS_OARG_1_GEN_TLAST(M_AXIS_OARG_1_GEN_TLAST),
        .M_AXIS_OARG_2_GEN_TLAST(M_AXIS_OARG_2_GEN_TLAST),
        .M_AXIS_OARG_3_GEN_TLAST(M_AXIS_OARG_3_GEN_TLAST),
        .M_AXIS_OARG_4_GEN_TLAST(M_AXIS_OARG_4_GEN_TLAST),
        .M_AXIS_OARG_5_GEN_TLAST(M_AXIS_OARG_5_GEN_TLAST),
        .M_AXIS_OARG_6_GEN_TLAST(M_AXIS_OARG_6_GEN_TLAST),
        .M_AXIS_OARG_7_GEN_TLAST(M_AXIS_OARG_7_GEN_TLAST),
        .M_AXIS_OARG_8_GEN_TLAST(M_AXIS_OARG_8_GEN_TLAST),
        .M_AXIS_OARG_9_GEN_TLAST(M_AXIS_OARG_9_GEN_TLAST),
        .M_AXIS_OARG_10_GEN_TLAST(M_AXIS_OARG_10_GEN_TLAST),
        .M_AXIS_OARG_11_GEN_TLAST(M_AXIS_OARG_11_GEN_TLAST),
        .M_AXIS_OARG_12_GEN_TLAST(M_AXIS_OARG_12_GEN_TLAST),
        .M_AXIS_OARG_13_GEN_TLAST(M_AXIS_OARG_13_GEN_TLAST),
        .M_AXIS_OARG_14_GEN_TLAST(M_AXIS_OARG_14_GEN_TLAST),
        .M_AXIS_OARG_15_GEN_TLAST(M_AXIS_OARG_15_GEN_TLAST),
        .M_AXIS_OARG_16_GEN_TLAST(M_AXIS_OARG_16_GEN_TLAST),
        .M_AXIS_OARG_17_GEN_TLAST(M_AXIS_OARG_17_GEN_TLAST),
        .M_AXIS_OARG_18_GEN_TLAST(M_AXIS_OARG_18_GEN_TLAST),
        .M_AXIS_OARG_19_GEN_TLAST(M_AXIS_OARG_19_GEN_TLAST),
        .M_AXIS_OARG_20_GEN_TLAST(M_AXIS_OARG_20_GEN_TLAST),
        .M_AXIS_OARG_21_GEN_TLAST(M_AXIS_OARG_21_GEN_TLAST),
        .M_AXIS_OARG_22_GEN_TLAST(M_AXIS_OARG_22_GEN_TLAST),
        .M_AXIS_OARG_23_GEN_TLAST(M_AXIS_OARG_23_GEN_TLAST),
        .M_AXIS_OARG_24_GEN_TLAST(M_AXIS_OARG_24_GEN_TLAST),
        .M_AXIS_OARG_25_GEN_TLAST(M_AXIS_OARG_25_GEN_TLAST),
        .M_AXIS_OARG_26_GEN_TLAST(M_AXIS_OARG_26_GEN_TLAST),
        .M_AXIS_OARG_27_GEN_TLAST(M_AXIS_OARG_27_GEN_TLAST),
        .M_AXIS_OARG_28_GEN_TLAST(M_AXIS_OARG_28_GEN_TLAST),
        .M_AXIS_OARG_29_GEN_TLAST(M_AXIS_OARG_29_GEN_TLAST),
        .M_AXIS_OARG_30_GEN_TLAST(M_AXIS_OARG_30_GEN_TLAST),
        .M_AXIS_OARG_31_GEN_TLAST(M_AXIS_OARG_31_GEN_TLAST),
        .M_AXIS_OARG_32_GEN_TLAST(M_AXIS_OARG_32_GEN_TLAST),
        .M_AXIS_OARG_33_GEN_TLAST(M_AXIS_OARG_33_GEN_TLAST),
        .M_AXIS_OARG_34_GEN_TLAST(M_AXIS_OARG_34_GEN_TLAST),
        .M_AXIS_OARG_35_GEN_TLAST(M_AXIS_OARG_35_GEN_TLAST),
        .M_AXIS_OARG_36_GEN_TLAST(M_AXIS_OARG_36_GEN_TLAST),
        .M_AXIS_OARG_37_GEN_TLAST(M_AXIS_OARG_37_GEN_TLAST),
        .M_AXIS_OARG_38_GEN_TLAST(M_AXIS_OARG_38_GEN_TLAST),
        .M_AXIS_OARG_39_GEN_TLAST(M_AXIS_OARG_39_GEN_TLAST),
        .M_AXIS_OARG_40_GEN_TLAST(M_AXIS_OARG_40_GEN_TLAST),
        .M_AXIS_OARG_41_GEN_TLAST(M_AXIS_OARG_41_GEN_TLAST),
        .M_AXIS_OARG_42_GEN_TLAST(M_AXIS_OARG_42_GEN_TLAST),
        .M_AXIS_OARG_43_GEN_TLAST(M_AXIS_OARG_43_GEN_TLAST),
        .M_AXIS_OARG_44_GEN_TLAST(M_AXIS_OARG_44_GEN_TLAST),
        .M_AXIS_OARG_45_GEN_TLAST(M_AXIS_OARG_45_GEN_TLAST),
        .M_AXIS_OARG_46_GEN_TLAST(M_AXIS_OARG_46_GEN_TLAST),
        .M_AXIS_OARG_47_GEN_TLAST(M_AXIS_OARG_47_GEN_TLAST),
        .M_AXIS_OARG_48_GEN_TLAST(M_AXIS_OARG_48_GEN_TLAST),
        .M_AXIS_OARG_49_GEN_TLAST(M_AXIS_OARG_49_GEN_TLAST),
        .M_AXIS_OARG_50_GEN_TLAST(M_AXIS_OARG_50_GEN_TLAST),
        .M_AXIS_OARG_51_GEN_TLAST(M_AXIS_OARG_51_GEN_TLAST),
        .M_AXIS_OARG_52_GEN_TLAST(M_AXIS_OARG_52_GEN_TLAST),
        .M_AXIS_OARG_53_GEN_TLAST(M_AXIS_OARG_53_GEN_TLAST),
        .M_AXIS_OARG_54_GEN_TLAST(M_AXIS_OARG_54_GEN_TLAST),
        .M_AXIS_OARG_55_GEN_TLAST(M_AXIS_OARG_55_GEN_TLAST),
        .M_AXIS_OARG_56_GEN_TLAST(M_AXIS_OARG_56_GEN_TLAST),
        .M_AXIS_OARG_57_GEN_TLAST(M_AXIS_OARG_57_GEN_TLAST),
        .M_AXIS_OARG_58_GEN_TLAST(M_AXIS_OARG_58_GEN_TLAST),
        .M_AXIS_OARG_59_GEN_TLAST(M_AXIS_OARG_59_GEN_TLAST),
        .M_AXIS_OARG_60_GEN_TLAST(M_AXIS_OARG_60_GEN_TLAST),
        .M_AXIS_OARG_61_GEN_TLAST(M_AXIS_OARG_61_GEN_TLAST),
        .M_AXIS_OARG_62_GEN_TLAST(M_AXIS_OARG_62_GEN_TLAST),
        .M_AXIS_OARG_63_GEN_TLAST(M_AXIS_OARG_63_GEN_TLAST),
        .M_AXIS_OARG_64_GEN_TLAST(M_AXIS_OARG_64_GEN_TLAST),
        .M_AXIS_OARG_65_GEN_TLAST(M_AXIS_OARG_65_GEN_TLAST),
        .M_AXIS_OARG_66_GEN_TLAST(M_AXIS_OARG_66_GEN_TLAST),
        .M_AXIS_OARG_67_GEN_TLAST(M_AXIS_OARG_67_GEN_TLAST),
        .M_AXIS_OARG_68_GEN_TLAST(M_AXIS_OARG_68_GEN_TLAST),
        .M_AXIS_OARG_69_GEN_TLAST(M_AXIS_OARG_69_GEN_TLAST),
        .M_AXIS_OARG_70_GEN_TLAST(M_AXIS_OARG_70_GEN_TLAST),
        .M_AXIS_OARG_71_GEN_TLAST(M_AXIS_OARG_71_GEN_TLAST),
        .M_AXIS_OARG_72_GEN_TLAST(M_AXIS_OARG_72_GEN_TLAST),
        .M_AXIS_OARG_73_GEN_TLAST(M_AXIS_OARG_73_GEN_TLAST),
        .M_AXIS_OARG_74_GEN_TLAST(M_AXIS_OARG_74_GEN_TLAST),
        .M_AXIS_OARG_75_GEN_TLAST(M_AXIS_OARG_75_GEN_TLAST),
        .M_AXIS_OARG_76_GEN_TLAST(M_AXIS_OARG_76_GEN_TLAST),
        .M_AXIS_OARG_77_GEN_TLAST(M_AXIS_OARG_77_GEN_TLAST),
        .M_AXIS_OARG_78_GEN_TLAST(M_AXIS_OARG_78_GEN_TLAST),
        .M_AXIS_OARG_79_GEN_TLAST(M_AXIS_OARG_79_GEN_TLAST),
        .M_AXIS_OARG_80_GEN_TLAST(M_AXIS_OARG_80_GEN_TLAST),
        .M_AXIS_OARG_81_GEN_TLAST(M_AXIS_OARG_81_GEN_TLAST),
        .M_AXIS_OARG_82_GEN_TLAST(M_AXIS_OARG_82_GEN_TLAST),
        .M_AXIS_OARG_83_GEN_TLAST(M_AXIS_OARG_83_GEN_TLAST),
        .M_AXIS_OARG_84_GEN_TLAST(M_AXIS_OARG_84_GEN_TLAST),
        .M_AXIS_OARG_85_GEN_TLAST(M_AXIS_OARG_85_GEN_TLAST),
        .M_AXIS_OARG_86_GEN_TLAST(M_AXIS_OARG_86_GEN_TLAST),
        .M_AXIS_OARG_87_GEN_TLAST(M_AXIS_OARG_87_GEN_TLAST),
        .M_AXIS_OARG_88_GEN_TLAST(M_AXIS_OARG_88_GEN_TLAST),
        .M_AXIS_OARG_89_GEN_TLAST(M_AXIS_OARG_89_GEN_TLAST),
        .M_AXIS_OARG_90_GEN_TLAST(M_AXIS_OARG_90_GEN_TLAST),
        .M_AXIS_OARG_91_GEN_TLAST(M_AXIS_OARG_91_GEN_TLAST),
        .M_AXIS_OARG_92_GEN_TLAST(M_AXIS_OARG_92_GEN_TLAST),
        .M_AXIS_OARG_93_GEN_TLAST(M_AXIS_OARG_93_GEN_TLAST),
        .M_AXIS_OARG_94_GEN_TLAST(M_AXIS_OARG_94_GEN_TLAST),
        .M_AXIS_OARG_95_GEN_TLAST(M_AXIS_OARG_95_GEN_TLAST),
        .M_AXIS_OARG_96_GEN_TLAST(M_AXIS_OARG_96_GEN_TLAST),
        .M_AXIS_OARG_97_GEN_TLAST(M_AXIS_OARG_97_GEN_TLAST),
        .M_AXIS_OARG_98_GEN_TLAST(M_AXIS_OARG_98_GEN_TLAST),
        .M_AXIS_OARG_99_GEN_TLAST(M_AXIS_OARG_99_GEN_TLAST),
        .M_AXIS_OARG_100_GEN_TLAST(M_AXIS_OARG_100_GEN_TLAST),
        .M_AXIS_OARG_101_GEN_TLAST(M_AXIS_OARG_101_GEN_TLAST),
        .M_AXIS_OARG_102_GEN_TLAST(M_AXIS_OARG_102_GEN_TLAST),
        .M_AXIS_OARG_103_GEN_TLAST(M_AXIS_OARG_103_GEN_TLAST),
        .M_AXIS_OARG_104_GEN_TLAST(M_AXIS_OARG_104_GEN_TLAST),
        .M_AXIS_OARG_105_GEN_TLAST(M_AXIS_OARG_105_GEN_TLAST),
        .M_AXIS_OARG_106_GEN_TLAST(M_AXIS_OARG_106_GEN_TLAST),
        .M_AXIS_OARG_107_GEN_TLAST(M_AXIS_OARG_107_GEN_TLAST),
        .M_AXIS_OARG_108_GEN_TLAST(M_AXIS_OARG_108_GEN_TLAST),
        .M_AXIS_OARG_109_GEN_TLAST(M_AXIS_OARG_109_GEN_TLAST),
        .M_AXIS_OARG_110_GEN_TLAST(M_AXIS_OARG_110_GEN_TLAST),
        .M_AXIS_OARG_111_GEN_TLAST(M_AXIS_OARG_111_GEN_TLAST),
        .M_AXIS_OARG_112_GEN_TLAST(M_AXIS_OARG_112_GEN_TLAST),
        .M_AXIS_OARG_113_GEN_TLAST(M_AXIS_OARG_113_GEN_TLAST),
        .M_AXIS_OARG_114_GEN_TLAST(M_AXIS_OARG_114_GEN_TLAST),
        .M_AXIS_OARG_115_GEN_TLAST(M_AXIS_OARG_115_GEN_TLAST),
        .M_AXIS_OARG_116_GEN_TLAST(M_AXIS_OARG_116_GEN_TLAST),
        .M_AXIS_OARG_117_GEN_TLAST(M_AXIS_OARG_117_GEN_TLAST),
        .M_AXIS_OARG_118_GEN_TLAST(M_AXIS_OARG_118_GEN_TLAST),
        .M_AXIS_OARG_119_GEN_TLAST(M_AXIS_OARG_119_GEN_TLAST),
        .M_AXIS_OARG_120_GEN_TLAST(M_AXIS_OARG_120_GEN_TLAST),
        .M_AXIS_OARG_121_GEN_TLAST(M_AXIS_OARG_121_GEN_TLAST),
        .M_AXIS_OARG_122_GEN_TLAST(M_AXIS_OARG_122_GEN_TLAST),
        .M_AXIS_OARG_123_GEN_TLAST(M_AXIS_OARG_123_GEN_TLAST),
        .M_AXIS_OARG_124_GEN_TLAST(M_AXIS_OARG_124_GEN_TLAST),
        .M_AXIS_OARG_125_GEN_TLAST(M_AXIS_OARG_125_GEN_TLAST),
        .M_AXIS_OARG_126_GEN_TLAST(M_AXIS_OARG_126_GEN_TLAST),
        .M_AXIS_OARG_127_GEN_TLAST(M_AXIS_OARG_127_GEN_TLAST),
        .M_AXIS_OARG_0_DMWIDTH(M_AXIS_OARG_0_DMWIDTH),
        .M_AXIS_OARG_1_DMWIDTH(M_AXIS_OARG_1_DMWIDTH),
        .M_AXIS_OARG_2_DMWIDTH(M_AXIS_OARG_2_DMWIDTH),
        .M_AXIS_OARG_3_DMWIDTH(M_AXIS_OARG_3_DMWIDTH),
        .M_AXIS_OARG_4_DMWIDTH(M_AXIS_OARG_4_DMWIDTH),
        .M_AXIS_OARG_5_DMWIDTH(M_AXIS_OARG_5_DMWIDTH),
        .M_AXIS_OARG_6_DMWIDTH(M_AXIS_OARG_6_DMWIDTH),
        .M_AXIS_OARG_7_DMWIDTH(M_AXIS_OARG_7_DMWIDTH),
        .M_AXIS_OARG_8_DMWIDTH(M_AXIS_OARG_8_DMWIDTH),
        .M_AXIS_OARG_9_DMWIDTH(M_AXIS_OARG_9_DMWIDTH),
        .M_AXIS_OARG_10_DMWIDTH(M_AXIS_OARG_10_DMWIDTH),
        .M_AXIS_OARG_11_DMWIDTH(M_AXIS_OARG_11_DMWIDTH),
        .M_AXIS_OARG_12_DMWIDTH(M_AXIS_OARG_12_DMWIDTH),
        .M_AXIS_OARG_13_DMWIDTH(M_AXIS_OARG_13_DMWIDTH),
        .M_AXIS_OARG_14_DMWIDTH(M_AXIS_OARG_14_DMWIDTH),
        .M_AXIS_OARG_15_DMWIDTH(M_AXIS_OARG_15_DMWIDTH),
        .M_AXIS_OARG_16_DMWIDTH(M_AXIS_OARG_16_DMWIDTH),
        .M_AXIS_OARG_17_DMWIDTH(M_AXIS_OARG_17_DMWIDTH),
        .M_AXIS_OARG_18_DMWIDTH(M_AXIS_OARG_18_DMWIDTH),
        .M_AXIS_OARG_19_DMWIDTH(M_AXIS_OARG_19_DMWIDTH),
        .M_AXIS_OARG_20_DMWIDTH(M_AXIS_OARG_20_DMWIDTH),
        .M_AXIS_OARG_21_DMWIDTH(M_AXIS_OARG_21_DMWIDTH),
        .M_AXIS_OARG_22_DMWIDTH(M_AXIS_OARG_22_DMWIDTH),
        .M_AXIS_OARG_23_DMWIDTH(M_AXIS_OARG_23_DMWIDTH),
        .M_AXIS_OARG_24_DMWIDTH(M_AXIS_OARG_24_DMWIDTH),
        .M_AXIS_OARG_25_DMWIDTH(M_AXIS_OARG_25_DMWIDTH),
        .M_AXIS_OARG_26_DMWIDTH(M_AXIS_OARG_26_DMWIDTH),
        .M_AXIS_OARG_27_DMWIDTH(M_AXIS_OARG_27_DMWIDTH),
        .M_AXIS_OARG_28_DMWIDTH(M_AXIS_OARG_28_DMWIDTH),
        .M_AXIS_OARG_29_DMWIDTH(M_AXIS_OARG_29_DMWIDTH),
        .M_AXIS_OARG_30_DMWIDTH(M_AXIS_OARG_30_DMWIDTH),
        .M_AXIS_OARG_31_DMWIDTH(M_AXIS_OARG_31_DMWIDTH),
        .M_AXIS_OARG_32_DMWIDTH(M_AXIS_OARG_32_DMWIDTH),
        .M_AXIS_OARG_33_DMWIDTH(M_AXIS_OARG_33_DMWIDTH),
        .M_AXIS_OARG_34_DMWIDTH(M_AXIS_OARG_34_DMWIDTH),
        .M_AXIS_OARG_35_DMWIDTH(M_AXIS_OARG_35_DMWIDTH),
        .M_AXIS_OARG_36_DMWIDTH(M_AXIS_OARG_36_DMWIDTH),
        .M_AXIS_OARG_37_DMWIDTH(M_AXIS_OARG_37_DMWIDTH),
        .M_AXIS_OARG_38_DMWIDTH(M_AXIS_OARG_38_DMWIDTH),
        .M_AXIS_OARG_39_DMWIDTH(M_AXIS_OARG_39_DMWIDTH),
        .M_AXIS_OARG_40_DMWIDTH(M_AXIS_OARG_40_DMWIDTH),
        .M_AXIS_OARG_41_DMWIDTH(M_AXIS_OARG_41_DMWIDTH),
        .M_AXIS_OARG_42_DMWIDTH(M_AXIS_OARG_42_DMWIDTH),
        .M_AXIS_OARG_43_DMWIDTH(M_AXIS_OARG_43_DMWIDTH),
        .M_AXIS_OARG_44_DMWIDTH(M_AXIS_OARG_44_DMWIDTH),
        .M_AXIS_OARG_45_DMWIDTH(M_AXIS_OARG_45_DMWIDTH),
        .M_AXIS_OARG_46_DMWIDTH(M_AXIS_OARG_46_DMWIDTH),
        .M_AXIS_OARG_47_DMWIDTH(M_AXIS_OARG_47_DMWIDTH),
        .M_AXIS_OARG_48_DMWIDTH(M_AXIS_OARG_48_DMWIDTH),
        .M_AXIS_OARG_49_DMWIDTH(M_AXIS_OARG_49_DMWIDTH),
        .M_AXIS_OARG_50_DMWIDTH(M_AXIS_OARG_50_DMWIDTH),
        .M_AXIS_OARG_51_DMWIDTH(M_AXIS_OARG_51_DMWIDTH),
        .M_AXIS_OARG_52_DMWIDTH(M_AXIS_OARG_52_DMWIDTH),
        .M_AXIS_OARG_53_DMWIDTH(M_AXIS_OARG_53_DMWIDTH),
        .M_AXIS_OARG_54_DMWIDTH(M_AXIS_OARG_54_DMWIDTH),
        .M_AXIS_OARG_55_DMWIDTH(M_AXIS_OARG_55_DMWIDTH),
        .M_AXIS_OARG_56_DMWIDTH(M_AXIS_OARG_56_DMWIDTH),
        .M_AXIS_OARG_57_DMWIDTH(M_AXIS_OARG_57_DMWIDTH),
        .M_AXIS_OARG_58_DMWIDTH(M_AXIS_OARG_58_DMWIDTH),
        .M_AXIS_OARG_59_DMWIDTH(M_AXIS_OARG_59_DMWIDTH),
        .M_AXIS_OARG_60_DMWIDTH(M_AXIS_OARG_60_DMWIDTH),
        .M_AXIS_OARG_61_DMWIDTH(M_AXIS_OARG_61_DMWIDTH),
        .M_AXIS_OARG_62_DMWIDTH(M_AXIS_OARG_62_DMWIDTH),
        .M_AXIS_OARG_63_DMWIDTH(M_AXIS_OARG_63_DMWIDTH),
        .M_AXIS_OARG_64_DMWIDTH(M_AXIS_OARG_64_DMWIDTH),
        .M_AXIS_OARG_65_DMWIDTH(M_AXIS_OARG_65_DMWIDTH),
        .M_AXIS_OARG_66_DMWIDTH(M_AXIS_OARG_66_DMWIDTH),
        .M_AXIS_OARG_67_DMWIDTH(M_AXIS_OARG_67_DMWIDTH),
        .M_AXIS_OARG_68_DMWIDTH(M_AXIS_OARG_68_DMWIDTH),
        .M_AXIS_OARG_69_DMWIDTH(M_AXIS_OARG_69_DMWIDTH),
        .M_AXIS_OARG_70_DMWIDTH(M_AXIS_OARG_70_DMWIDTH),
        .M_AXIS_OARG_71_DMWIDTH(M_AXIS_OARG_71_DMWIDTH),
        .M_AXIS_OARG_72_DMWIDTH(M_AXIS_OARG_72_DMWIDTH),
        .M_AXIS_OARG_73_DMWIDTH(M_AXIS_OARG_73_DMWIDTH),
        .M_AXIS_OARG_74_DMWIDTH(M_AXIS_OARG_74_DMWIDTH),
        .M_AXIS_OARG_75_DMWIDTH(M_AXIS_OARG_75_DMWIDTH),
        .M_AXIS_OARG_76_DMWIDTH(M_AXIS_OARG_76_DMWIDTH),
        .M_AXIS_OARG_77_DMWIDTH(M_AXIS_OARG_77_DMWIDTH),
        .M_AXIS_OARG_78_DMWIDTH(M_AXIS_OARG_78_DMWIDTH),
        .M_AXIS_OARG_79_DMWIDTH(M_AXIS_OARG_79_DMWIDTH),
        .M_AXIS_OARG_80_DMWIDTH(M_AXIS_OARG_80_DMWIDTH),
        .M_AXIS_OARG_81_DMWIDTH(M_AXIS_OARG_81_DMWIDTH),
        .M_AXIS_OARG_82_DMWIDTH(M_AXIS_OARG_82_DMWIDTH),
        .M_AXIS_OARG_83_DMWIDTH(M_AXIS_OARG_83_DMWIDTH),
        .M_AXIS_OARG_84_DMWIDTH(M_AXIS_OARG_84_DMWIDTH),
        .M_AXIS_OARG_85_DMWIDTH(M_AXIS_OARG_85_DMWIDTH),
        .M_AXIS_OARG_86_DMWIDTH(M_AXIS_OARG_86_DMWIDTH),
        .M_AXIS_OARG_87_DMWIDTH(M_AXIS_OARG_87_DMWIDTH),
        .M_AXIS_OARG_88_DMWIDTH(M_AXIS_OARG_88_DMWIDTH),
        .M_AXIS_OARG_89_DMWIDTH(M_AXIS_OARG_89_DMWIDTH),
        .M_AXIS_OARG_90_DMWIDTH(M_AXIS_OARG_90_DMWIDTH),
        .M_AXIS_OARG_91_DMWIDTH(M_AXIS_OARG_91_DMWIDTH),
        .M_AXIS_OARG_92_DMWIDTH(M_AXIS_OARG_92_DMWIDTH),
        .M_AXIS_OARG_93_DMWIDTH(M_AXIS_OARG_93_DMWIDTH),
        .M_AXIS_OARG_94_DMWIDTH(M_AXIS_OARG_94_DMWIDTH),
        .M_AXIS_OARG_95_DMWIDTH(M_AXIS_OARG_95_DMWIDTH),
        .M_AXIS_OARG_96_DMWIDTH(M_AXIS_OARG_96_DMWIDTH),
        .M_AXIS_OARG_97_DMWIDTH(M_AXIS_OARG_97_DMWIDTH),
        .M_AXIS_OARG_98_DMWIDTH(M_AXIS_OARG_98_DMWIDTH),
        .M_AXIS_OARG_99_DMWIDTH(M_AXIS_OARG_99_DMWIDTH),
        .M_AXIS_OARG_100_DMWIDTH(M_AXIS_OARG_100_DMWIDTH),
        .M_AXIS_OARG_101_DMWIDTH(M_AXIS_OARG_101_DMWIDTH),
        .M_AXIS_OARG_102_DMWIDTH(M_AXIS_OARG_102_DMWIDTH),
        .M_AXIS_OARG_103_DMWIDTH(M_AXIS_OARG_103_DMWIDTH),
        .M_AXIS_OARG_104_DMWIDTH(M_AXIS_OARG_104_DMWIDTH),
        .M_AXIS_OARG_105_DMWIDTH(M_AXIS_OARG_105_DMWIDTH),
        .M_AXIS_OARG_106_DMWIDTH(M_AXIS_OARG_106_DMWIDTH),
        .M_AXIS_OARG_107_DMWIDTH(M_AXIS_OARG_107_DMWIDTH),
        .M_AXIS_OARG_108_DMWIDTH(M_AXIS_OARG_108_DMWIDTH),
        .M_AXIS_OARG_109_DMWIDTH(M_AXIS_OARG_109_DMWIDTH),
        .M_AXIS_OARG_110_DMWIDTH(M_AXIS_OARG_110_DMWIDTH),
        .M_AXIS_OARG_111_DMWIDTH(M_AXIS_OARG_111_DMWIDTH),
        .M_AXIS_OARG_112_DMWIDTH(M_AXIS_OARG_112_DMWIDTH),
        .M_AXIS_OARG_113_DMWIDTH(M_AXIS_OARG_113_DMWIDTH),
        .M_AXIS_OARG_114_DMWIDTH(M_AXIS_OARG_114_DMWIDTH),
        .M_AXIS_OARG_115_DMWIDTH(M_AXIS_OARG_115_DMWIDTH),
        .M_AXIS_OARG_116_DMWIDTH(M_AXIS_OARG_116_DMWIDTH),
        .M_AXIS_OARG_117_DMWIDTH(M_AXIS_OARG_117_DMWIDTH),
        .M_AXIS_OARG_118_DMWIDTH(M_AXIS_OARG_118_DMWIDTH),
        .M_AXIS_OARG_119_DMWIDTH(M_AXIS_OARG_119_DMWIDTH),
        .M_AXIS_OARG_120_DMWIDTH(M_AXIS_OARG_120_DMWIDTH),
        .M_AXIS_OARG_121_DMWIDTH(M_AXIS_OARG_121_DMWIDTH),
        .M_AXIS_OARG_122_DMWIDTH(M_AXIS_OARG_122_DMWIDTH),
        .M_AXIS_OARG_123_DMWIDTH(M_AXIS_OARG_123_DMWIDTH),
        .M_AXIS_OARG_124_DMWIDTH(M_AXIS_OARG_124_DMWIDTH),
        .M_AXIS_OARG_125_DMWIDTH(M_AXIS_OARG_125_DMWIDTH),
        .M_AXIS_OARG_126_DMWIDTH(M_AXIS_OARG_126_DMWIDTH),
        .M_AXIS_OARG_127_DMWIDTH(M_AXIS_OARG_127_DMWIDTH)
    ) out_axis_args_i (
        .acc_clk(acc_aclk),
        .acc_aresetn(acc_aresetn),
        .out_axis_allow(outaxis_ctrl_allow),
        .m_axis_oarg_0_aclk(m_axis_oarg_0_aclk),
        .m_axis_oarg_0_aresetn(m_axis_oarg_0_aresetn),
        .m_axis_oarg_0_tlast(m_axis_oarg_0_tlast),
        .m_axis_oarg_0_tvalid(m_axis_oarg_0_tvalid),
        .m_axis_oarg_0_tkeep(m_axis_oarg_0_tkeep),
        .m_axis_oarg_0_tstrb(m_axis_oarg_0_tstrb),
        .m_axis_oarg_0_tdata(m_axis_oarg_0_tdata),
        .m_axis_oarg_0_tready(m_axis_oarg_0_tready),
        .ap_axis_oarg_0_tlast(ap_axis_oarg_0_tlast),
        .ap_axis_oarg_0_tvalid(ap_axis_oarg_0_tvalid),
        .ap_axis_oarg_0_tkeep(ap_axis_oarg_0_tkeep),
        .ap_axis_oarg_0_tstrb(ap_axis_oarg_0_tstrb),
        .ap_axis_oarg_0_tdata(ap_axis_oarg_0_tdata),
        .ap_axis_oarg_0_tready(ap_axis_oarg_0_tready),
        .m_axis_oarg_1_aclk(m_axis_oarg_1_aclk),
        .m_axis_oarg_1_aresetn(m_axis_oarg_1_aresetn),
        .m_axis_oarg_1_tlast(m_axis_oarg_1_tlast),
        .m_axis_oarg_1_tvalid(m_axis_oarg_1_tvalid),
        .m_axis_oarg_1_tkeep(m_axis_oarg_1_tkeep),
        .m_axis_oarg_1_tstrb(m_axis_oarg_1_tstrb),
        .m_axis_oarg_1_tdata(m_axis_oarg_1_tdata),
        .m_axis_oarg_1_tready(m_axis_oarg_1_tready),
        .ap_axis_oarg_1_tlast(ap_axis_oarg_1_tlast),
        .ap_axis_oarg_1_tvalid(ap_axis_oarg_1_tvalid),
        .ap_axis_oarg_1_tkeep(ap_axis_oarg_1_tkeep),
        .ap_axis_oarg_1_tstrb(ap_axis_oarg_1_tstrb),
        .ap_axis_oarg_1_tdata(ap_axis_oarg_1_tdata),
        .ap_axis_oarg_1_tready(ap_axis_oarg_1_tready),
        .m_axis_oarg_2_aclk(m_axis_oarg_2_aclk),
        .m_axis_oarg_2_aresetn(m_axis_oarg_2_aresetn),
        .m_axis_oarg_2_tlast(m_axis_oarg_2_tlast),
        .m_axis_oarg_2_tvalid(m_axis_oarg_2_tvalid),
        .m_axis_oarg_2_tkeep(m_axis_oarg_2_tkeep),
        .m_axis_oarg_2_tstrb(m_axis_oarg_2_tstrb),
        .m_axis_oarg_2_tdata(m_axis_oarg_2_tdata),
        .m_axis_oarg_2_tready(m_axis_oarg_2_tready),
        .ap_axis_oarg_2_tlast(ap_axis_oarg_2_tlast),
        .ap_axis_oarg_2_tvalid(ap_axis_oarg_2_tvalid),
        .ap_axis_oarg_2_tkeep(ap_axis_oarg_2_tkeep),
        .ap_axis_oarg_2_tstrb(ap_axis_oarg_2_tstrb),
        .ap_axis_oarg_2_tdata(ap_axis_oarg_2_tdata),
        .ap_axis_oarg_2_tready(ap_axis_oarg_2_tready),
        .m_axis_oarg_3_aclk(m_axis_oarg_3_aclk),
        .m_axis_oarg_3_aresetn(m_axis_oarg_3_aresetn),
        .m_axis_oarg_3_tlast(m_axis_oarg_3_tlast),
        .m_axis_oarg_3_tvalid(m_axis_oarg_3_tvalid),
        .m_axis_oarg_3_tkeep(m_axis_oarg_3_tkeep),
        .m_axis_oarg_3_tstrb(m_axis_oarg_3_tstrb),
        .m_axis_oarg_3_tdata(m_axis_oarg_3_tdata),
        .m_axis_oarg_3_tready(m_axis_oarg_3_tready),
        .ap_axis_oarg_3_tlast(ap_axis_oarg_3_tlast),
        .ap_axis_oarg_3_tvalid(ap_axis_oarg_3_tvalid),
        .ap_axis_oarg_3_tkeep(ap_axis_oarg_3_tkeep),
        .ap_axis_oarg_3_tstrb(ap_axis_oarg_3_tstrb),
        .ap_axis_oarg_3_tdata(ap_axis_oarg_3_tdata),
        .ap_axis_oarg_3_tready(ap_axis_oarg_3_tready),
        .m_axis_oarg_4_aclk(m_axis_oarg_4_aclk),
        .m_axis_oarg_4_aresetn(m_axis_oarg_4_aresetn),
        .m_axis_oarg_4_tlast(m_axis_oarg_4_tlast),
        .m_axis_oarg_4_tvalid(m_axis_oarg_4_tvalid),
        .m_axis_oarg_4_tkeep(m_axis_oarg_4_tkeep),
        .m_axis_oarg_4_tstrb(m_axis_oarg_4_tstrb),
        .m_axis_oarg_4_tdata(m_axis_oarg_4_tdata),
        .m_axis_oarg_4_tready(m_axis_oarg_4_tready),
        .ap_axis_oarg_4_tlast(ap_axis_oarg_4_tlast),
        .ap_axis_oarg_4_tvalid(ap_axis_oarg_4_tvalid),
        .ap_axis_oarg_4_tkeep(ap_axis_oarg_4_tkeep),
        .ap_axis_oarg_4_tstrb(ap_axis_oarg_4_tstrb),
        .ap_axis_oarg_4_tdata(ap_axis_oarg_4_tdata),
        .ap_axis_oarg_4_tready(ap_axis_oarg_4_tready),
        .m_axis_oarg_5_aclk(m_axis_oarg_5_aclk),
        .m_axis_oarg_5_aresetn(m_axis_oarg_5_aresetn),
        .m_axis_oarg_5_tlast(m_axis_oarg_5_tlast),
        .m_axis_oarg_5_tvalid(m_axis_oarg_5_tvalid),
        .m_axis_oarg_5_tkeep(m_axis_oarg_5_tkeep),
        .m_axis_oarg_5_tstrb(m_axis_oarg_5_tstrb),
        .m_axis_oarg_5_tdata(m_axis_oarg_5_tdata),
        .m_axis_oarg_5_tready(m_axis_oarg_5_tready),
        .ap_axis_oarg_5_tlast(ap_axis_oarg_5_tlast),
        .ap_axis_oarg_5_tvalid(ap_axis_oarg_5_tvalid),
        .ap_axis_oarg_5_tkeep(ap_axis_oarg_5_tkeep),
        .ap_axis_oarg_5_tstrb(ap_axis_oarg_5_tstrb),
        .ap_axis_oarg_5_tdata(ap_axis_oarg_5_tdata),
        .ap_axis_oarg_5_tready(ap_axis_oarg_5_tready),
        .m_axis_oarg_6_aclk(m_axis_oarg_6_aclk),
        .m_axis_oarg_6_aresetn(m_axis_oarg_6_aresetn),
        .m_axis_oarg_6_tlast(m_axis_oarg_6_tlast),
        .m_axis_oarg_6_tvalid(m_axis_oarg_6_tvalid),
        .m_axis_oarg_6_tkeep(m_axis_oarg_6_tkeep),
        .m_axis_oarg_6_tstrb(m_axis_oarg_6_tstrb),
        .m_axis_oarg_6_tdata(m_axis_oarg_6_tdata),
        .m_axis_oarg_6_tready(m_axis_oarg_6_tready),
        .ap_axis_oarg_6_tlast(ap_axis_oarg_6_tlast),
        .ap_axis_oarg_6_tvalid(ap_axis_oarg_6_tvalid),
        .ap_axis_oarg_6_tkeep(ap_axis_oarg_6_tkeep),
        .ap_axis_oarg_6_tstrb(ap_axis_oarg_6_tstrb),
        .ap_axis_oarg_6_tdata(ap_axis_oarg_6_tdata),
        .ap_axis_oarg_6_tready(ap_axis_oarg_6_tready),
        .m_axis_oarg_7_aclk(m_axis_oarg_7_aclk),
        .m_axis_oarg_7_aresetn(m_axis_oarg_7_aresetn),
        .m_axis_oarg_7_tlast(m_axis_oarg_7_tlast),
        .m_axis_oarg_7_tvalid(m_axis_oarg_7_tvalid),
        .m_axis_oarg_7_tkeep(m_axis_oarg_7_tkeep),
        .m_axis_oarg_7_tstrb(m_axis_oarg_7_tstrb),
        .m_axis_oarg_7_tdata(m_axis_oarg_7_tdata),
        .m_axis_oarg_7_tready(m_axis_oarg_7_tready),
        .ap_axis_oarg_7_tlast(ap_axis_oarg_7_tlast),
        .ap_axis_oarg_7_tvalid(ap_axis_oarg_7_tvalid),
        .ap_axis_oarg_7_tkeep(ap_axis_oarg_7_tkeep),
        .ap_axis_oarg_7_tstrb(ap_axis_oarg_7_tstrb),
        .ap_axis_oarg_7_tdata(ap_axis_oarg_7_tdata),
        .ap_axis_oarg_7_tready(ap_axis_oarg_7_tready),
        .m_axis_oarg_8_aclk(m_axis_oarg_8_aclk),
        .m_axis_oarg_8_aresetn(m_axis_oarg_8_aresetn),
        .m_axis_oarg_8_tlast(m_axis_oarg_8_tlast),
        .m_axis_oarg_8_tvalid(m_axis_oarg_8_tvalid),
        .m_axis_oarg_8_tkeep(m_axis_oarg_8_tkeep),
        .m_axis_oarg_8_tstrb(m_axis_oarg_8_tstrb),
        .m_axis_oarg_8_tdata(m_axis_oarg_8_tdata),
        .m_axis_oarg_8_tready(m_axis_oarg_8_tready),
        .ap_axis_oarg_8_tlast(ap_axis_oarg_8_tlast),
        .ap_axis_oarg_8_tvalid(ap_axis_oarg_8_tvalid),
        .ap_axis_oarg_8_tkeep(ap_axis_oarg_8_tkeep),
        .ap_axis_oarg_8_tstrb(ap_axis_oarg_8_tstrb),
        .ap_axis_oarg_8_tdata(ap_axis_oarg_8_tdata),
        .ap_axis_oarg_8_tready(ap_axis_oarg_8_tready),
        .m_axis_oarg_9_aclk(m_axis_oarg_9_aclk),
        .m_axis_oarg_9_aresetn(m_axis_oarg_9_aresetn),
        .m_axis_oarg_9_tlast(m_axis_oarg_9_tlast),
        .m_axis_oarg_9_tvalid(m_axis_oarg_9_tvalid),
        .m_axis_oarg_9_tkeep(m_axis_oarg_9_tkeep),
        .m_axis_oarg_9_tstrb(m_axis_oarg_9_tstrb),
        .m_axis_oarg_9_tdata(m_axis_oarg_9_tdata),
        .m_axis_oarg_9_tready(m_axis_oarg_9_tready),
        .ap_axis_oarg_9_tlast(ap_axis_oarg_9_tlast),
        .ap_axis_oarg_9_tvalid(ap_axis_oarg_9_tvalid),
        .ap_axis_oarg_9_tkeep(ap_axis_oarg_9_tkeep),
        .ap_axis_oarg_9_tstrb(ap_axis_oarg_9_tstrb),
        .ap_axis_oarg_9_tdata(ap_axis_oarg_9_tdata),
        .ap_axis_oarg_9_tready(ap_axis_oarg_9_tready),
        .m_axis_oarg_10_aclk(m_axis_oarg_10_aclk),
        .m_axis_oarg_10_aresetn(m_axis_oarg_10_aresetn),
        .m_axis_oarg_10_tlast(m_axis_oarg_10_tlast),
        .m_axis_oarg_10_tvalid(m_axis_oarg_10_tvalid),
        .m_axis_oarg_10_tkeep(m_axis_oarg_10_tkeep),
        .m_axis_oarg_10_tstrb(m_axis_oarg_10_tstrb),
        .m_axis_oarg_10_tdata(m_axis_oarg_10_tdata),
        .m_axis_oarg_10_tready(m_axis_oarg_10_tready),
        .ap_axis_oarg_10_tlast(ap_axis_oarg_10_tlast),
        .ap_axis_oarg_10_tvalid(ap_axis_oarg_10_tvalid),
        .ap_axis_oarg_10_tkeep(ap_axis_oarg_10_tkeep),
        .ap_axis_oarg_10_tstrb(ap_axis_oarg_10_tstrb),
        .ap_axis_oarg_10_tdata(ap_axis_oarg_10_tdata),
        .ap_axis_oarg_10_tready(ap_axis_oarg_10_tready),
        .m_axis_oarg_11_aclk(m_axis_oarg_11_aclk),
        .m_axis_oarg_11_aresetn(m_axis_oarg_11_aresetn),
        .m_axis_oarg_11_tlast(m_axis_oarg_11_tlast),
        .m_axis_oarg_11_tvalid(m_axis_oarg_11_tvalid),
        .m_axis_oarg_11_tkeep(m_axis_oarg_11_tkeep),
        .m_axis_oarg_11_tstrb(m_axis_oarg_11_tstrb),
        .m_axis_oarg_11_tdata(m_axis_oarg_11_tdata),
        .m_axis_oarg_11_tready(m_axis_oarg_11_tready),
        .ap_axis_oarg_11_tlast(ap_axis_oarg_11_tlast),
        .ap_axis_oarg_11_tvalid(ap_axis_oarg_11_tvalid),
        .ap_axis_oarg_11_tkeep(ap_axis_oarg_11_tkeep),
        .ap_axis_oarg_11_tstrb(ap_axis_oarg_11_tstrb),
        .ap_axis_oarg_11_tdata(ap_axis_oarg_11_tdata),
        .ap_axis_oarg_11_tready(ap_axis_oarg_11_tready),
        .m_axis_oarg_12_aclk(m_axis_oarg_12_aclk),
        .m_axis_oarg_12_aresetn(m_axis_oarg_12_aresetn),
        .m_axis_oarg_12_tlast(m_axis_oarg_12_tlast),
        .m_axis_oarg_12_tvalid(m_axis_oarg_12_tvalid),
        .m_axis_oarg_12_tkeep(m_axis_oarg_12_tkeep),
        .m_axis_oarg_12_tstrb(m_axis_oarg_12_tstrb),
        .m_axis_oarg_12_tdata(m_axis_oarg_12_tdata),
        .m_axis_oarg_12_tready(m_axis_oarg_12_tready),
        .ap_axis_oarg_12_tlast(ap_axis_oarg_12_tlast),
        .ap_axis_oarg_12_tvalid(ap_axis_oarg_12_tvalid),
        .ap_axis_oarg_12_tkeep(ap_axis_oarg_12_tkeep),
        .ap_axis_oarg_12_tstrb(ap_axis_oarg_12_tstrb),
        .ap_axis_oarg_12_tdata(ap_axis_oarg_12_tdata),
        .ap_axis_oarg_12_tready(ap_axis_oarg_12_tready),
        .m_axis_oarg_13_aclk(m_axis_oarg_13_aclk),
        .m_axis_oarg_13_aresetn(m_axis_oarg_13_aresetn),
        .m_axis_oarg_13_tlast(m_axis_oarg_13_tlast),
        .m_axis_oarg_13_tvalid(m_axis_oarg_13_tvalid),
        .m_axis_oarg_13_tkeep(m_axis_oarg_13_tkeep),
        .m_axis_oarg_13_tstrb(m_axis_oarg_13_tstrb),
        .m_axis_oarg_13_tdata(m_axis_oarg_13_tdata),
        .m_axis_oarg_13_tready(m_axis_oarg_13_tready),
        .ap_axis_oarg_13_tlast(ap_axis_oarg_13_tlast),
        .ap_axis_oarg_13_tvalid(ap_axis_oarg_13_tvalid),
        .ap_axis_oarg_13_tkeep(ap_axis_oarg_13_tkeep),
        .ap_axis_oarg_13_tstrb(ap_axis_oarg_13_tstrb),
        .ap_axis_oarg_13_tdata(ap_axis_oarg_13_tdata),
        .ap_axis_oarg_13_tready(ap_axis_oarg_13_tready),
        .m_axis_oarg_14_aclk(m_axis_oarg_14_aclk),
        .m_axis_oarg_14_aresetn(m_axis_oarg_14_aresetn),
        .m_axis_oarg_14_tlast(m_axis_oarg_14_tlast),
        .m_axis_oarg_14_tvalid(m_axis_oarg_14_tvalid),
        .m_axis_oarg_14_tkeep(m_axis_oarg_14_tkeep),
        .m_axis_oarg_14_tstrb(m_axis_oarg_14_tstrb),
        .m_axis_oarg_14_tdata(m_axis_oarg_14_tdata),
        .m_axis_oarg_14_tready(m_axis_oarg_14_tready),
        .ap_axis_oarg_14_tlast(ap_axis_oarg_14_tlast),
        .ap_axis_oarg_14_tvalid(ap_axis_oarg_14_tvalid),
        .ap_axis_oarg_14_tkeep(ap_axis_oarg_14_tkeep),
        .ap_axis_oarg_14_tstrb(ap_axis_oarg_14_tstrb),
        .ap_axis_oarg_14_tdata(ap_axis_oarg_14_tdata),
        .ap_axis_oarg_14_tready(ap_axis_oarg_14_tready),
        .m_axis_oarg_15_aclk(m_axis_oarg_15_aclk),
        .m_axis_oarg_15_aresetn(m_axis_oarg_15_aresetn),
        .m_axis_oarg_15_tlast(m_axis_oarg_15_tlast),
        .m_axis_oarg_15_tvalid(m_axis_oarg_15_tvalid),
        .m_axis_oarg_15_tkeep(m_axis_oarg_15_tkeep),
        .m_axis_oarg_15_tstrb(m_axis_oarg_15_tstrb),
        .m_axis_oarg_15_tdata(m_axis_oarg_15_tdata),
        .m_axis_oarg_15_tready(m_axis_oarg_15_tready),
        .ap_axis_oarg_15_tlast(ap_axis_oarg_15_tlast),
        .ap_axis_oarg_15_tvalid(ap_axis_oarg_15_tvalid),
        .ap_axis_oarg_15_tkeep(ap_axis_oarg_15_tkeep),
        .ap_axis_oarg_15_tstrb(ap_axis_oarg_15_tstrb),
        .ap_axis_oarg_15_tdata(ap_axis_oarg_15_tdata),
        .ap_axis_oarg_15_tready(ap_axis_oarg_15_tready),
        .m_axis_oarg_16_aclk(m_axis_oarg_16_aclk),
        .m_axis_oarg_16_aresetn(m_axis_oarg_16_aresetn),
        .m_axis_oarg_16_tlast(m_axis_oarg_16_tlast),
        .m_axis_oarg_16_tvalid(m_axis_oarg_16_tvalid),
        .m_axis_oarg_16_tkeep(m_axis_oarg_16_tkeep),
        .m_axis_oarg_16_tstrb(m_axis_oarg_16_tstrb),
        .m_axis_oarg_16_tdata(m_axis_oarg_16_tdata),
        .m_axis_oarg_16_tready(m_axis_oarg_16_tready),
        .ap_axis_oarg_16_tlast(ap_axis_oarg_16_tlast),
        .ap_axis_oarg_16_tvalid(ap_axis_oarg_16_tvalid),
        .ap_axis_oarg_16_tkeep(ap_axis_oarg_16_tkeep),
        .ap_axis_oarg_16_tstrb(ap_axis_oarg_16_tstrb),
        .ap_axis_oarg_16_tdata(ap_axis_oarg_16_tdata),
        .ap_axis_oarg_16_tready(ap_axis_oarg_16_tready),
        .m_axis_oarg_17_aclk(m_axis_oarg_17_aclk),
        .m_axis_oarg_17_aresetn(m_axis_oarg_17_aresetn),
        .m_axis_oarg_17_tlast(m_axis_oarg_17_tlast),
        .m_axis_oarg_17_tvalid(m_axis_oarg_17_tvalid),
        .m_axis_oarg_17_tkeep(m_axis_oarg_17_tkeep),
        .m_axis_oarg_17_tstrb(m_axis_oarg_17_tstrb),
        .m_axis_oarg_17_tdata(m_axis_oarg_17_tdata),
        .m_axis_oarg_17_tready(m_axis_oarg_17_tready),
        .ap_axis_oarg_17_tlast(ap_axis_oarg_17_tlast),
        .ap_axis_oarg_17_tvalid(ap_axis_oarg_17_tvalid),
        .ap_axis_oarg_17_tkeep(ap_axis_oarg_17_tkeep),
        .ap_axis_oarg_17_tstrb(ap_axis_oarg_17_tstrb),
        .ap_axis_oarg_17_tdata(ap_axis_oarg_17_tdata),
        .ap_axis_oarg_17_tready(ap_axis_oarg_17_tready),
        .m_axis_oarg_18_aclk(m_axis_oarg_18_aclk),
        .m_axis_oarg_18_aresetn(m_axis_oarg_18_aresetn),
        .m_axis_oarg_18_tlast(m_axis_oarg_18_tlast),
        .m_axis_oarg_18_tvalid(m_axis_oarg_18_tvalid),
        .m_axis_oarg_18_tkeep(m_axis_oarg_18_tkeep),
        .m_axis_oarg_18_tstrb(m_axis_oarg_18_tstrb),
        .m_axis_oarg_18_tdata(m_axis_oarg_18_tdata),
        .m_axis_oarg_18_tready(m_axis_oarg_18_tready),
        .ap_axis_oarg_18_tlast(ap_axis_oarg_18_tlast),
        .ap_axis_oarg_18_tvalid(ap_axis_oarg_18_tvalid),
        .ap_axis_oarg_18_tkeep(ap_axis_oarg_18_tkeep),
        .ap_axis_oarg_18_tstrb(ap_axis_oarg_18_tstrb),
        .ap_axis_oarg_18_tdata(ap_axis_oarg_18_tdata),
        .ap_axis_oarg_18_tready(ap_axis_oarg_18_tready),
        .m_axis_oarg_19_aclk(m_axis_oarg_19_aclk),
        .m_axis_oarg_19_aresetn(m_axis_oarg_19_aresetn),
        .m_axis_oarg_19_tlast(m_axis_oarg_19_tlast),
        .m_axis_oarg_19_tvalid(m_axis_oarg_19_tvalid),
        .m_axis_oarg_19_tkeep(m_axis_oarg_19_tkeep),
        .m_axis_oarg_19_tstrb(m_axis_oarg_19_tstrb),
        .m_axis_oarg_19_tdata(m_axis_oarg_19_tdata),
        .m_axis_oarg_19_tready(m_axis_oarg_19_tready),
        .ap_axis_oarg_19_tlast(ap_axis_oarg_19_tlast),
        .ap_axis_oarg_19_tvalid(ap_axis_oarg_19_tvalid),
        .ap_axis_oarg_19_tkeep(ap_axis_oarg_19_tkeep),
        .ap_axis_oarg_19_tstrb(ap_axis_oarg_19_tstrb),
        .ap_axis_oarg_19_tdata(ap_axis_oarg_19_tdata),
        .ap_axis_oarg_19_tready(ap_axis_oarg_19_tready),
        .m_axis_oarg_20_aclk(m_axis_oarg_20_aclk),
        .m_axis_oarg_20_aresetn(m_axis_oarg_20_aresetn),
        .m_axis_oarg_20_tlast(m_axis_oarg_20_tlast),
        .m_axis_oarg_20_tvalid(m_axis_oarg_20_tvalid),
        .m_axis_oarg_20_tkeep(m_axis_oarg_20_tkeep),
        .m_axis_oarg_20_tstrb(m_axis_oarg_20_tstrb),
        .m_axis_oarg_20_tdata(m_axis_oarg_20_tdata),
        .m_axis_oarg_20_tready(m_axis_oarg_20_tready),
        .ap_axis_oarg_20_tlast(ap_axis_oarg_20_tlast),
        .ap_axis_oarg_20_tvalid(ap_axis_oarg_20_tvalid),
        .ap_axis_oarg_20_tkeep(ap_axis_oarg_20_tkeep),
        .ap_axis_oarg_20_tstrb(ap_axis_oarg_20_tstrb),
        .ap_axis_oarg_20_tdata(ap_axis_oarg_20_tdata),
        .ap_axis_oarg_20_tready(ap_axis_oarg_20_tready),
        .m_axis_oarg_21_aclk(m_axis_oarg_21_aclk),
        .m_axis_oarg_21_aresetn(m_axis_oarg_21_aresetn),
        .m_axis_oarg_21_tlast(m_axis_oarg_21_tlast),
        .m_axis_oarg_21_tvalid(m_axis_oarg_21_tvalid),
        .m_axis_oarg_21_tkeep(m_axis_oarg_21_tkeep),
        .m_axis_oarg_21_tstrb(m_axis_oarg_21_tstrb),
        .m_axis_oarg_21_tdata(m_axis_oarg_21_tdata),
        .m_axis_oarg_21_tready(m_axis_oarg_21_tready),
        .ap_axis_oarg_21_tlast(ap_axis_oarg_21_tlast),
        .ap_axis_oarg_21_tvalid(ap_axis_oarg_21_tvalid),
        .ap_axis_oarg_21_tkeep(ap_axis_oarg_21_tkeep),
        .ap_axis_oarg_21_tstrb(ap_axis_oarg_21_tstrb),
        .ap_axis_oarg_21_tdata(ap_axis_oarg_21_tdata),
        .ap_axis_oarg_21_tready(ap_axis_oarg_21_tready),
        .m_axis_oarg_22_aclk(m_axis_oarg_22_aclk),
        .m_axis_oarg_22_aresetn(m_axis_oarg_22_aresetn),
        .m_axis_oarg_22_tlast(m_axis_oarg_22_tlast),
        .m_axis_oarg_22_tvalid(m_axis_oarg_22_tvalid),
        .m_axis_oarg_22_tkeep(m_axis_oarg_22_tkeep),
        .m_axis_oarg_22_tstrb(m_axis_oarg_22_tstrb),
        .m_axis_oarg_22_tdata(m_axis_oarg_22_tdata),
        .m_axis_oarg_22_tready(m_axis_oarg_22_tready),
        .ap_axis_oarg_22_tlast(ap_axis_oarg_22_tlast),
        .ap_axis_oarg_22_tvalid(ap_axis_oarg_22_tvalid),
        .ap_axis_oarg_22_tkeep(ap_axis_oarg_22_tkeep),
        .ap_axis_oarg_22_tstrb(ap_axis_oarg_22_tstrb),
        .ap_axis_oarg_22_tdata(ap_axis_oarg_22_tdata),
        .ap_axis_oarg_22_tready(ap_axis_oarg_22_tready),
        .m_axis_oarg_23_aclk(m_axis_oarg_23_aclk),
        .m_axis_oarg_23_aresetn(m_axis_oarg_23_aresetn),
        .m_axis_oarg_23_tlast(m_axis_oarg_23_tlast),
        .m_axis_oarg_23_tvalid(m_axis_oarg_23_tvalid),
        .m_axis_oarg_23_tkeep(m_axis_oarg_23_tkeep),
        .m_axis_oarg_23_tstrb(m_axis_oarg_23_tstrb),
        .m_axis_oarg_23_tdata(m_axis_oarg_23_tdata),
        .m_axis_oarg_23_tready(m_axis_oarg_23_tready),
        .ap_axis_oarg_23_tlast(ap_axis_oarg_23_tlast),
        .ap_axis_oarg_23_tvalid(ap_axis_oarg_23_tvalid),
        .ap_axis_oarg_23_tkeep(ap_axis_oarg_23_tkeep),
        .ap_axis_oarg_23_tstrb(ap_axis_oarg_23_tstrb),
        .ap_axis_oarg_23_tdata(ap_axis_oarg_23_tdata),
        .ap_axis_oarg_23_tready(ap_axis_oarg_23_tready),
        .m_axis_oarg_24_aclk(m_axis_oarg_24_aclk),
        .m_axis_oarg_24_aresetn(m_axis_oarg_24_aresetn),
        .m_axis_oarg_24_tlast(m_axis_oarg_24_tlast),
        .m_axis_oarg_24_tvalid(m_axis_oarg_24_tvalid),
        .m_axis_oarg_24_tkeep(m_axis_oarg_24_tkeep),
        .m_axis_oarg_24_tstrb(m_axis_oarg_24_tstrb),
        .m_axis_oarg_24_tdata(m_axis_oarg_24_tdata),
        .m_axis_oarg_24_tready(m_axis_oarg_24_tready),
        .ap_axis_oarg_24_tlast(ap_axis_oarg_24_tlast),
        .ap_axis_oarg_24_tvalid(ap_axis_oarg_24_tvalid),
        .ap_axis_oarg_24_tkeep(ap_axis_oarg_24_tkeep),
        .ap_axis_oarg_24_tstrb(ap_axis_oarg_24_tstrb),
        .ap_axis_oarg_24_tdata(ap_axis_oarg_24_tdata),
        .ap_axis_oarg_24_tready(ap_axis_oarg_24_tready),
        .m_axis_oarg_25_aclk(m_axis_oarg_25_aclk),
        .m_axis_oarg_25_aresetn(m_axis_oarg_25_aresetn),
        .m_axis_oarg_25_tlast(m_axis_oarg_25_tlast),
        .m_axis_oarg_25_tvalid(m_axis_oarg_25_tvalid),
        .m_axis_oarg_25_tkeep(m_axis_oarg_25_tkeep),
        .m_axis_oarg_25_tstrb(m_axis_oarg_25_tstrb),
        .m_axis_oarg_25_tdata(m_axis_oarg_25_tdata),
        .m_axis_oarg_25_tready(m_axis_oarg_25_tready),
        .ap_axis_oarg_25_tlast(ap_axis_oarg_25_tlast),
        .ap_axis_oarg_25_tvalid(ap_axis_oarg_25_tvalid),
        .ap_axis_oarg_25_tkeep(ap_axis_oarg_25_tkeep),
        .ap_axis_oarg_25_tstrb(ap_axis_oarg_25_tstrb),
        .ap_axis_oarg_25_tdata(ap_axis_oarg_25_tdata),
        .ap_axis_oarg_25_tready(ap_axis_oarg_25_tready),
        .m_axis_oarg_26_aclk(m_axis_oarg_26_aclk),
        .m_axis_oarg_26_aresetn(m_axis_oarg_26_aresetn),
        .m_axis_oarg_26_tlast(m_axis_oarg_26_tlast),
        .m_axis_oarg_26_tvalid(m_axis_oarg_26_tvalid),
        .m_axis_oarg_26_tkeep(m_axis_oarg_26_tkeep),
        .m_axis_oarg_26_tstrb(m_axis_oarg_26_tstrb),
        .m_axis_oarg_26_tdata(m_axis_oarg_26_tdata),
        .m_axis_oarg_26_tready(m_axis_oarg_26_tready),
        .ap_axis_oarg_26_tlast(ap_axis_oarg_26_tlast),
        .ap_axis_oarg_26_tvalid(ap_axis_oarg_26_tvalid),
        .ap_axis_oarg_26_tkeep(ap_axis_oarg_26_tkeep),
        .ap_axis_oarg_26_tstrb(ap_axis_oarg_26_tstrb),
        .ap_axis_oarg_26_tdata(ap_axis_oarg_26_tdata),
        .ap_axis_oarg_26_tready(ap_axis_oarg_26_tready),
        .m_axis_oarg_27_aclk(m_axis_oarg_27_aclk),
        .m_axis_oarg_27_aresetn(m_axis_oarg_27_aresetn),
        .m_axis_oarg_27_tlast(m_axis_oarg_27_tlast),
        .m_axis_oarg_27_tvalid(m_axis_oarg_27_tvalid),
        .m_axis_oarg_27_tkeep(m_axis_oarg_27_tkeep),
        .m_axis_oarg_27_tstrb(m_axis_oarg_27_tstrb),
        .m_axis_oarg_27_tdata(m_axis_oarg_27_tdata),
        .m_axis_oarg_27_tready(m_axis_oarg_27_tready),
        .ap_axis_oarg_27_tlast(ap_axis_oarg_27_tlast),
        .ap_axis_oarg_27_tvalid(ap_axis_oarg_27_tvalid),
        .ap_axis_oarg_27_tkeep(ap_axis_oarg_27_tkeep),
        .ap_axis_oarg_27_tstrb(ap_axis_oarg_27_tstrb),
        .ap_axis_oarg_27_tdata(ap_axis_oarg_27_tdata),
        .ap_axis_oarg_27_tready(ap_axis_oarg_27_tready),
        .m_axis_oarg_28_aclk(m_axis_oarg_28_aclk),
        .m_axis_oarg_28_aresetn(m_axis_oarg_28_aresetn),
        .m_axis_oarg_28_tlast(m_axis_oarg_28_tlast),
        .m_axis_oarg_28_tvalid(m_axis_oarg_28_tvalid),
        .m_axis_oarg_28_tkeep(m_axis_oarg_28_tkeep),
        .m_axis_oarg_28_tstrb(m_axis_oarg_28_tstrb),
        .m_axis_oarg_28_tdata(m_axis_oarg_28_tdata),
        .m_axis_oarg_28_tready(m_axis_oarg_28_tready),
        .ap_axis_oarg_28_tlast(ap_axis_oarg_28_tlast),
        .ap_axis_oarg_28_tvalid(ap_axis_oarg_28_tvalid),
        .ap_axis_oarg_28_tkeep(ap_axis_oarg_28_tkeep),
        .ap_axis_oarg_28_tstrb(ap_axis_oarg_28_tstrb),
        .ap_axis_oarg_28_tdata(ap_axis_oarg_28_tdata),
        .ap_axis_oarg_28_tready(ap_axis_oarg_28_tready),
        .m_axis_oarg_29_aclk(m_axis_oarg_29_aclk),
        .m_axis_oarg_29_aresetn(m_axis_oarg_29_aresetn),
        .m_axis_oarg_29_tlast(m_axis_oarg_29_tlast),
        .m_axis_oarg_29_tvalid(m_axis_oarg_29_tvalid),
        .m_axis_oarg_29_tkeep(m_axis_oarg_29_tkeep),
        .m_axis_oarg_29_tstrb(m_axis_oarg_29_tstrb),
        .m_axis_oarg_29_tdata(m_axis_oarg_29_tdata),
        .m_axis_oarg_29_tready(m_axis_oarg_29_tready),
        .ap_axis_oarg_29_tlast(ap_axis_oarg_29_tlast),
        .ap_axis_oarg_29_tvalid(ap_axis_oarg_29_tvalid),
        .ap_axis_oarg_29_tkeep(ap_axis_oarg_29_tkeep),
        .ap_axis_oarg_29_tstrb(ap_axis_oarg_29_tstrb),
        .ap_axis_oarg_29_tdata(ap_axis_oarg_29_tdata),
        .ap_axis_oarg_29_tready(ap_axis_oarg_29_tready),
        .m_axis_oarg_30_aclk(m_axis_oarg_30_aclk),
        .m_axis_oarg_30_aresetn(m_axis_oarg_30_aresetn),
        .m_axis_oarg_30_tlast(m_axis_oarg_30_tlast),
        .m_axis_oarg_30_tvalid(m_axis_oarg_30_tvalid),
        .m_axis_oarg_30_tkeep(m_axis_oarg_30_tkeep),
        .m_axis_oarg_30_tstrb(m_axis_oarg_30_tstrb),
        .m_axis_oarg_30_tdata(m_axis_oarg_30_tdata),
        .m_axis_oarg_30_tready(m_axis_oarg_30_tready),
        .ap_axis_oarg_30_tlast(ap_axis_oarg_30_tlast),
        .ap_axis_oarg_30_tvalid(ap_axis_oarg_30_tvalid),
        .ap_axis_oarg_30_tkeep(ap_axis_oarg_30_tkeep),
        .ap_axis_oarg_30_tstrb(ap_axis_oarg_30_tstrb),
        .ap_axis_oarg_30_tdata(ap_axis_oarg_30_tdata),
        .ap_axis_oarg_30_tready(ap_axis_oarg_30_tready),
        .m_axis_oarg_31_aclk(m_axis_oarg_31_aclk),
        .m_axis_oarg_31_aresetn(m_axis_oarg_31_aresetn),
        .m_axis_oarg_31_tlast(m_axis_oarg_31_tlast),
        .m_axis_oarg_31_tvalid(m_axis_oarg_31_tvalid),
        .m_axis_oarg_31_tkeep(m_axis_oarg_31_tkeep),
        .m_axis_oarg_31_tstrb(m_axis_oarg_31_tstrb),
        .m_axis_oarg_31_tdata(m_axis_oarg_31_tdata),
        .m_axis_oarg_31_tready(m_axis_oarg_31_tready),
        .ap_axis_oarg_31_tlast(ap_axis_oarg_31_tlast),
        .ap_axis_oarg_31_tvalid(ap_axis_oarg_31_tvalid),
        .ap_axis_oarg_31_tkeep(ap_axis_oarg_31_tkeep),
        .ap_axis_oarg_31_tstrb(ap_axis_oarg_31_tstrb),
        .ap_axis_oarg_31_tdata(ap_axis_oarg_31_tdata),
        .ap_axis_oarg_31_tready(ap_axis_oarg_31_tready),
        .m_axis_oarg_32_aclk(m_axis_oarg_32_aclk),
        .m_axis_oarg_32_aresetn(m_axis_oarg_32_aresetn),
        .m_axis_oarg_32_tlast(m_axis_oarg_32_tlast),
        .m_axis_oarg_32_tvalid(m_axis_oarg_32_tvalid),
        .m_axis_oarg_32_tkeep(m_axis_oarg_32_tkeep),
        .m_axis_oarg_32_tstrb(m_axis_oarg_32_tstrb),
        .m_axis_oarg_32_tdata(m_axis_oarg_32_tdata),
        .m_axis_oarg_32_tready(m_axis_oarg_32_tready),
        .ap_axis_oarg_32_tlast(ap_axis_oarg_32_tlast),
        .ap_axis_oarg_32_tvalid(ap_axis_oarg_32_tvalid),
        .ap_axis_oarg_32_tkeep(ap_axis_oarg_32_tkeep),
        .ap_axis_oarg_32_tstrb(ap_axis_oarg_32_tstrb),
        .ap_axis_oarg_32_tdata(ap_axis_oarg_32_tdata),
        .ap_axis_oarg_32_tready(ap_axis_oarg_32_tready),
        .m_axis_oarg_33_aclk(m_axis_oarg_33_aclk),
        .m_axis_oarg_33_aresetn(m_axis_oarg_33_aresetn),
        .m_axis_oarg_33_tlast(m_axis_oarg_33_tlast),
        .m_axis_oarg_33_tvalid(m_axis_oarg_33_tvalid),
        .m_axis_oarg_33_tkeep(m_axis_oarg_33_tkeep),
        .m_axis_oarg_33_tstrb(m_axis_oarg_33_tstrb),
        .m_axis_oarg_33_tdata(m_axis_oarg_33_tdata),
        .m_axis_oarg_33_tready(m_axis_oarg_33_tready),
        .ap_axis_oarg_33_tlast(ap_axis_oarg_33_tlast),
        .ap_axis_oarg_33_tvalid(ap_axis_oarg_33_tvalid),
        .ap_axis_oarg_33_tkeep(ap_axis_oarg_33_tkeep),
        .ap_axis_oarg_33_tstrb(ap_axis_oarg_33_tstrb),
        .ap_axis_oarg_33_tdata(ap_axis_oarg_33_tdata),
        .ap_axis_oarg_33_tready(ap_axis_oarg_33_tready),
        .m_axis_oarg_34_aclk(m_axis_oarg_34_aclk),
        .m_axis_oarg_34_aresetn(m_axis_oarg_34_aresetn),
        .m_axis_oarg_34_tlast(m_axis_oarg_34_tlast),
        .m_axis_oarg_34_tvalid(m_axis_oarg_34_tvalid),
        .m_axis_oarg_34_tkeep(m_axis_oarg_34_tkeep),
        .m_axis_oarg_34_tstrb(m_axis_oarg_34_tstrb),
        .m_axis_oarg_34_tdata(m_axis_oarg_34_tdata),
        .m_axis_oarg_34_tready(m_axis_oarg_34_tready),
        .ap_axis_oarg_34_tlast(ap_axis_oarg_34_tlast),
        .ap_axis_oarg_34_tvalid(ap_axis_oarg_34_tvalid),
        .ap_axis_oarg_34_tkeep(ap_axis_oarg_34_tkeep),
        .ap_axis_oarg_34_tstrb(ap_axis_oarg_34_tstrb),
        .ap_axis_oarg_34_tdata(ap_axis_oarg_34_tdata),
        .ap_axis_oarg_34_tready(ap_axis_oarg_34_tready),
        .m_axis_oarg_35_aclk(m_axis_oarg_35_aclk),
        .m_axis_oarg_35_aresetn(m_axis_oarg_35_aresetn),
        .m_axis_oarg_35_tlast(m_axis_oarg_35_tlast),
        .m_axis_oarg_35_tvalid(m_axis_oarg_35_tvalid),
        .m_axis_oarg_35_tkeep(m_axis_oarg_35_tkeep),
        .m_axis_oarg_35_tstrb(m_axis_oarg_35_tstrb),
        .m_axis_oarg_35_tdata(m_axis_oarg_35_tdata),
        .m_axis_oarg_35_tready(m_axis_oarg_35_tready),
        .ap_axis_oarg_35_tlast(ap_axis_oarg_35_tlast),
        .ap_axis_oarg_35_tvalid(ap_axis_oarg_35_tvalid),
        .ap_axis_oarg_35_tkeep(ap_axis_oarg_35_tkeep),
        .ap_axis_oarg_35_tstrb(ap_axis_oarg_35_tstrb),
        .ap_axis_oarg_35_tdata(ap_axis_oarg_35_tdata),
        .ap_axis_oarg_35_tready(ap_axis_oarg_35_tready),
        .m_axis_oarg_36_aclk(m_axis_oarg_36_aclk),
        .m_axis_oarg_36_aresetn(m_axis_oarg_36_aresetn),
        .m_axis_oarg_36_tlast(m_axis_oarg_36_tlast),
        .m_axis_oarg_36_tvalid(m_axis_oarg_36_tvalid),
        .m_axis_oarg_36_tkeep(m_axis_oarg_36_tkeep),
        .m_axis_oarg_36_tstrb(m_axis_oarg_36_tstrb),
        .m_axis_oarg_36_tdata(m_axis_oarg_36_tdata),
        .m_axis_oarg_36_tready(m_axis_oarg_36_tready),
        .ap_axis_oarg_36_tlast(ap_axis_oarg_36_tlast),
        .ap_axis_oarg_36_tvalid(ap_axis_oarg_36_tvalid),
        .ap_axis_oarg_36_tkeep(ap_axis_oarg_36_tkeep),
        .ap_axis_oarg_36_tstrb(ap_axis_oarg_36_tstrb),
        .ap_axis_oarg_36_tdata(ap_axis_oarg_36_tdata),
        .ap_axis_oarg_36_tready(ap_axis_oarg_36_tready),
        .m_axis_oarg_37_aclk(m_axis_oarg_37_aclk),
        .m_axis_oarg_37_aresetn(m_axis_oarg_37_aresetn),
        .m_axis_oarg_37_tlast(m_axis_oarg_37_tlast),
        .m_axis_oarg_37_tvalid(m_axis_oarg_37_tvalid),
        .m_axis_oarg_37_tkeep(m_axis_oarg_37_tkeep),
        .m_axis_oarg_37_tstrb(m_axis_oarg_37_tstrb),
        .m_axis_oarg_37_tdata(m_axis_oarg_37_tdata),
        .m_axis_oarg_37_tready(m_axis_oarg_37_tready),
        .ap_axis_oarg_37_tlast(ap_axis_oarg_37_tlast),
        .ap_axis_oarg_37_tvalid(ap_axis_oarg_37_tvalid),
        .ap_axis_oarg_37_tkeep(ap_axis_oarg_37_tkeep),
        .ap_axis_oarg_37_tstrb(ap_axis_oarg_37_tstrb),
        .ap_axis_oarg_37_tdata(ap_axis_oarg_37_tdata),
        .ap_axis_oarg_37_tready(ap_axis_oarg_37_tready),
        .m_axis_oarg_38_aclk(m_axis_oarg_38_aclk),
        .m_axis_oarg_38_aresetn(m_axis_oarg_38_aresetn),
        .m_axis_oarg_38_tlast(m_axis_oarg_38_tlast),
        .m_axis_oarg_38_tvalid(m_axis_oarg_38_tvalid),
        .m_axis_oarg_38_tkeep(m_axis_oarg_38_tkeep),
        .m_axis_oarg_38_tstrb(m_axis_oarg_38_tstrb),
        .m_axis_oarg_38_tdata(m_axis_oarg_38_tdata),
        .m_axis_oarg_38_tready(m_axis_oarg_38_tready),
        .ap_axis_oarg_38_tlast(ap_axis_oarg_38_tlast),
        .ap_axis_oarg_38_tvalid(ap_axis_oarg_38_tvalid),
        .ap_axis_oarg_38_tkeep(ap_axis_oarg_38_tkeep),
        .ap_axis_oarg_38_tstrb(ap_axis_oarg_38_tstrb),
        .ap_axis_oarg_38_tdata(ap_axis_oarg_38_tdata),
        .ap_axis_oarg_38_tready(ap_axis_oarg_38_tready),
        .m_axis_oarg_39_aclk(m_axis_oarg_39_aclk),
        .m_axis_oarg_39_aresetn(m_axis_oarg_39_aresetn),
        .m_axis_oarg_39_tlast(m_axis_oarg_39_tlast),
        .m_axis_oarg_39_tvalid(m_axis_oarg_39_tvalid),
        .m_axis_oarg_39_tkeep(m_axis_oarg_39_tkeep),
        .m_axis_oarg_39_tstrb(m_axis_oarg_39_tstrb),
        .m_axis_oarg_39_tdata(m_axis_oarg_39_tdata),
        .m_axis_oarg_39_tready(m_axis_oarg_39_tready),
        .ap_axis_oarg_39_tlast(ap_axis_oarg_39_tlast),
        .ap_axis_oarg_39_tvalid(ap_axis_oarg_39_tvalid),
        .ap_axis_oarg_39_tkeep(ap_axis_oarg_39_tkeep),
        .ap_axis_oarg_39_tstrb(ap_axis_oarg_39_tstrb),
        .ap_axis_oarg_39_tdata(ap_axis_oarg_39_tdata),
        .ap_axis_oarg_39_tready(ap_axis_oarg_39_tready),
        .m_axis_oarg_40_aclk(m_axis_oarg_40_aclk),
        .m_axis_oarg_40_aresetn(m_axis_oarg_40_aresetn),
        .m_axis_oarg_40_tlast(m_axis_oarg_40_tlast),
        .m_axis_oarg_40_tvalid(m_axis_oarg_40_tvalid),
        .m_axis_oarg_40_tkeep(m_axis_oarg_40_tkeep),
        .m_axis_oarg_40_tstrb(m_axis_oarg_40_tstrb),
        .m_axis_oarg_40_tdata(m_axis_oarg_40_tdata),
        .m_axis_oarg_40_tready(m_axis_oarg_40_tready),
        .ap_axis_oarg_40_tlast(ap_axis_oarg_40_tlast),
        .ap_axis_oarg_40_tvalid(ap_axis_oarg_40_tvalid),
        .ap_axis_oarg_40_tkeep(ap_axis_oarg_40_tkeep),
        .ap_axis_oarg_40_tstrb(ap_axis_oarg_40_tstrb),
        .ap_axis_oarg_40_tdata(ap_axis_oarg_40_tdata),
        .ap_axis_oarg_40_tready(ap_axis_oarg_40_tready),
        .m_axis_oarg_41_aclk(m_axis_oarg_41_aclk),
        .m_axis_oarg_41_aresetn(m_axis_oarg_41_aresetn),
        .m_axis_oarg_41_tlast(m_axis_oarg_41_tlast),
        .m_axis_oarg_41_tvalid(m_axis_oarg_41_tvalid),
        .m_axis_oarg_41_tkeep(m_axis_oarg_41_tkeep),
        .m_axis_oarg_41_tstrb(m_axis_oarg_41_tstrb),
        .m_axis_oarg_41_tdata(m_axis_oarg_41_tdata),
        .m_axis_oarg_41_tready(m_axis_oarg_41_tready),
        .ap_axis_oarg_41_tlast(ap_axis_oarg_41_tlast),
        .ap_axis_oarg_41_tvalid(ap_axis_oarg_41_tvalid),
        .ap_axis_oarg_41_tkeep(ap_axis_oarg_41_tkeep),
        .ap_axis_oarg_41_tstrb(ap_axis_oarg_41_tstrb),
        .ap_axis_oarg_41_tdata(ap_axis_oarg_41_tdata),
        .ap_axis_oarg_41_tready(ap_axis_oarg_41_tready),
        .m_axis_oarg_42_aclk(m_axis_oarg_42_aclk),
        .m_axis_oarg_42_aresetn(m_axis_oarg_42_aresetn),
        .m_axis_oarg_42_tlast(m_axis_oarg_42_tlast),
        .m_axis_oarg_42_tvalid(m_axis_oarg_42_tvalid),
        .m_axis_oarg_42_tkeep(m_axis_oarg_42_tkeep),
        .m_axis_oarg_42_tstrb(m_axis_oarg_42_tstrb),
        .m_axis_oarg_42_tdata(m_axis_oarg_42_tdata),
        .m_axis_oarg_42_tready(m_axis_oarg_42_tready),
        .ap_axis_oarg_42_tlast(ap_axis_oarg_42_tlast),
        .ap_axis_oarg_42_tvalid(ap_axis_oarg_42_tvalid),
        .ap_axis_oarg_42_tkeep(ap_axis_oarg_42_tkeep),
        .ap_axis_oarg_42_tstrb(ap_axis_oarg_42_tstrb),
        .ap_axis_oarg_42_tdata(ap_axis_oarg_42_tdata),
        .ap_axis_oarg_42_tready(ap_axis_oarg_42_tready),
        .m_axis_oarg_43_aclk(m_axis_oarg_43_aclk),
        .m_axis_oarg_43_aresetn(m_axis_oarg_43_aresetn),
        .m_axis_oarg_43_tlast(m_axis_oarg_43_tlast),
        .m_axis_oarg_43_tvalid(m_axis_oarg_43_tvalid),
        .m_axis_oarg_43_tkeep(m_axis_oarg_43_tkeep),
        .m_axis_oarg_43_tstrb(m_axis_oarg_43_tstrb),
        .m_axis_oarg_43_tdata(m_axis_oarg_43_tdata),
        .m_axis_oarg_43_tready(m_axis_oarg_43_tready),
        .ap_axis_oarg_43_tlast(ap_axis_oarg_43_tlast),
        .ap_axis_oarg_43_tvalid(ap_axis_oarg_43_tvalid),
        .ap_axis_oarg_43_tkeep(ap_axis_oarg_43_tkeep),
        .ap_axis_oarg_43_tstrb(ap_axis_oarg_43_tstrb),
        .ap_axis_oarg_43_tdata(ap_axis_oarg_43_tdata),
        .ap_axis_oarg_43_tready(ap_axis_oarg_43_tready),
        .m_axis_oarg_44_aclk(m_axis_oarg_44_aclk),
        .m_axis_oarg_44_aresetn(m_axis_oarg_44_aresetn),
        .m_axis_oarg_44_tlast(m_axis_oarg_44_tlast),
        .m_axis_oarg_44_tvalid(m_axis_oarg_44_tvalid),
        .m_axis_oarg_44_tkeep(m_axis_oarg_44_tkeep),
        .m_axis_oarg_44_tstrb(m_axis_oarg_44_tstrb),
        .m_axis_oarg_44_tdata(m_axis_oarg_44_tdata),
        .m_axis_oarg_44_tready(m_axis_oarg_44_tready),
        .ap_axis_oarg_44_tlast(ap_axis_oarg_44_tlast),
        .ap_axis_oarg_44_tvalid(ap_axis_oarg_44_tvalid),
        .ap_axis_oarg_44_tkeep(ap_axis_oarg_44_tkeep),
        .ap_axis_oarg_44_tstrb(ap_axis_oarg_44_tstrb),
        .ap_axis_oarg_44_tdata(ap_axis_oarg_44_tdata),
        .ap_axis_oarg_44_tready(ap_axis_oarg_44_tready),
        .m_axis_oarg_45_aclk(m_axis_oarg_45_aclk),
        .m_axis_oarg_45_aresetn(m_axis_oarg_45_aresetn),
        .m_axis_oarg_45_tlast(m_axis_oarg_45_tlast),
        .m_axis_oarg_45_tvalid(m_axis_oarg_45_tvalid),
        .m_axis_oarg_45_tkeep(m_axis_oarg_45_tkeep),
        .m_axis_oarg_45_tstrb(m_axis_oarg_45_tstrb),
        .m_axis_oarg_45_tdata(m_axis_oarg_45_tdata),
        .m_axis_oarg_45_tready(m_axis_oarg_45_tready),
        .ap_axis_oarg_45_tlast(ap_axis_oarg_45_tlast),
        .ap_axis_oarg_45_tvalid(ap_axis_oarg_45_tvalid),
        .ap_axis_oarg_45_tkeep(ap_axis_oarg_45_tkeep),
        .ap_axis_oarg_45_tstrb(ap_axis_oarg_45_tstrb),
        .ap_axis_oarg_45_tdata(ap_axis_oarg_45_tdata),
        .ap_axis_oarg_45_tready(ap_axis_oarg_45_tready),
        .m_axis_oarg_46_aclk(m_axis_oarg_46_aclk),
        .m_axis_oarg_46_aresetn(m_axis_oarg_46_aresetn),
        .m_axis_oarg_46_tlast(m_axis_oarg_46_tlast),
        .m_axis_oarg_46_tvalid(m_axis_oarg_46_tvalid),
        .m_axis_oarg_46_tkeep(m_axis_oarg_46_tkeep),
        .m_axis_oarg_46_tstrb(m_axis_oarg_46_tstrb),
        .m_axis_oarg_46_tdata(m_axis_oarg_46_tdata),
        .m_axis_oarg_46_tready(m_axis_oarg_46_tready),
        .ap_axis_oarg_46_tlast(ap_axis_oarg_46_tlast),
        .ap_axis_oarg_46_tvalid(ap_axis_oarg_46_tvalid),
        .ap_axis_oarg_46_tkeep(ap_axis_oarg_46_tkeep),
        .ap_axis_oarg_46_tstrb(ap_axis_oarg_46_tstrb),
        .ap_axis_oarg_46_tdata(ap_axis_oarg_46_tdata),
        .ap_axis_oarg_46_tready(ap_axis_oarg_46_tready),
        .m_axis_oarg_47_aclk(m_axis_oarg_47_aclk),
        .m_axis_oarg_47_aresetn(m_axis_oarg_47_aresetn),
        .m_axis_oarg_47_tlast(m_axis_oarg_47_tlast),
        .m_axis_oarg_47_tvalid(m_axis_oarg_47_tvalid),
        .m_axis_oarg_47_tkeep(m_axis_oarg_47_tkeep),
        .m_axis_oarg_47_tstrb(m_axis_oarg_47_tstrb),
        .m_axis_oarg_47_tdata(m_axis_oarg_47_tdata),
        .m_axis_oarg_47_tready(m_axis_oarg_47_tready),
        .ap_axis_oarg_47_tlast(ap_axis_oarg_47_tlast),
        .ap_axis_oarg_47_tvalid(ap_axis_oarg_47_tvalid),
        .ap_axis_oarg_47_tkeep(ap_axis_oarg_47_tkeep),
        .ap_axis_oarg_47_tstrb(ap_axis_oarg_47_tstrb),
        .ap_axis_oarg_47_tdata(ap_axis_oarg_47_tdata),
        .ap_axis_oarg_47_tready(ap_axis_oarg_47_tready),
        .m_axis_oarg_48_aclk(m_axis_oarg_48_aclk),
        .m_axis_oarg_48_aresetn(m_axis_oarg_48_aresetn),
        .m_axis_oarg_48_tlast(m_axis_oarg_48_tlast),
        .m_axis_oarg_48_tvalid(m_axis_oarg_48_tvalid),
        .m_axis_oarg_48_tkeep(m_axis_oarg_48_tkeep),
        .m_axis_oarg_48_tstrb(m_axis_oarg_48_tstrb),
        .m_axis_oarg_48_tdata(m_axis_oarg_48_tdata),
        .m_axis_oarg_48_tready(m_axis_oarg_48_tready),
        .ap_axis_oarg_48_tlast(ap_axis_oarg_48_tlast),
        .ap_axis_oarg_48_tvalid(ap_axis_oarg_48_tvalid),
        .ap_axis_oarg_48_tkeep(ap_axis_oarg_48_tkeep),
        .ap_axis_oarg_48_tstrb(ap_axis_oarg_48_tstrb),
        .ap_axis_oarg_48_tdata(ap_axis_oarg_48_tdata),
        .ap_axis_oarg_48_tready(ap_axis_oarg_48_tready),
        .m_axis_oarg_49_aclk(m_axis_oarg_49_aclk),
        .m_axis_oarg_49_aresetn(m_axis_oarg_49_aresetn),
        .m_axis_oarg_49_tlast(m_axis_oarg_49_tlast),
        .m_axis_oarg_49_tvalid(m_axis_oarg_49_tvalid),
        .m_axis_oarg_49_tkeep(m_axis_oarg_49_tkeep),
        .m_axis_oarg_49_tstrb(m_axis_oarg_49_tstrb),
        .m_axis_oarg_49_tdata(m_axis_oarg_49_tdata),
        .m_axis_oarg_49_tready(m_axis_oarg_49_tready),
        .ap_axis_oarg_49_tlast(ap_axis_oarg_49_tlast),
        .ap_axis_oarg_49_tvalid(ap_axis_oarg_49_tvalid),
        .ap_axis_oarg_49_tkeep(ap_axis_oarg_49_tkeep),
        .ap_axis_oarg_49_tstrb(ap_axis_oarg_49_tstrb),
        .ap_axis_oarg_49_tdata(ap_axis_oarg_49_tdata),
        .ap_axis_oarg_49_tready(ap_axis_oarg_49_tready),
        .m_axis_oarg_50_aclk(m_axis_oarg_50_aclk),
        .m_axis_oarg_50_aresetn(m_axis_oarg_50_aresetn),
        .m_axis_oarg_50_tlast(m_axis_oarg_50_tlast),
        .m_axis_oarg_50_tvalid(m_axis_oarg_50_tvalid),
        .m_axis_oarg_50_tkeep(m_axis_oarg_50_tkeep),
        .m_axis_oarg_50_tstrb(m_axis_oarg_50_tstrb),
        .m_axis_oarg_50_tdata(m_axis_oarg_50_tdata),
        .m_axis_oarg_50_tready(m_axis_oarg_50_tready),
        .ap_axis_oarg_50_tlast(ap_axis_oarg_50_tlast),
        .ap_axis_oarg_50_tvalid(ap_axis_oarg_50_tvalid),
        .ap_axis_oarg_50_tkeep(ap_axis_oarg_50_tkeep),
        .ap_axis_oarg_50_tstrb(ap_axis_oarg_50_tstrb),
        .ap_axis_oarg_50_tdata(ap_axis_oarg_50_tdata),
        .ap_axis_oarg_50_tready(ap_axis_oarg_50_tready),
        .m_axis_oarg_51_aclk(m_axis_oarg_51_aclk),
        .m_axis_oarg_51_aresetn(m_axis_oarg_51_aresetn),
        .m_axis_oarg_51_tlast(m_axis_oarg_51_tlast),
        .m_axis_oarg_51_tvalid(m_axis_oarg_51_tvalid),
        .m_axis_oarg_51_tkeep(m_axis_oarg_51_tkeep),
        .m_axis_oarg_51_tstrb(m_axis_oarg_51_tstrb),
        .m_axis_oarg_51_tdata(m_axis_oarg_51_tdata),
        .m_axis_oarg_51_tready(m_axis_oarg_51_tready),
        .ap_axis_oarg_51_tlast(ap_axis_oarg_51_tlast),
        .ap_axis_oarg_51_tvalid(ap_axis_oarg_51_tvalid),
        .ap_axis_oarg_51_tkeep(ap_axis_oarg_51_tkeep),
        .ap_axis_oarg_51_tstrb(ap_axis_oarg_51_tstrb),
        .ap_axis_oarg_51_tdata(ap_axis_oarg_51_tdata),
        .ap_axis_oarg_51_tready(ap_axis_oarg_51_tready),
        .m_axis_oarg_52_aclk(m_axis_oarg_52_aclk),
        .m_axis_oarg_52_aresetn(m_axis_oarg_52_aresetn),
        .m_axis_oarg_52_tlast(m_axis_oarg_52_tlast),
        .m_axis_oarg_52_tvalid(m_axis_oarg_52_tvalid),
        .m_axis_oarg_52_tkeep(m_axis_oarg_52_tkeep),
        .m_axis_oarg_52_tstrb(m_axis_oarg_52_tstrb),
        .m_axis_oarg_52_tdata(m_axis_oarg_52_tdata),
        .m_axis_oarg_52_tready(m_axis_oarg_52_tready),
        .ap_axis_oarg_52_tlast(ap_axis_oarg_52_tlast),
        .ap_axis_oarg_52_tvalid(ap_axis_oarg_52_tvalid),
        .ap_axis_oarg_52_tkeep(ap_axis_oarg_52_tkeep),
        .ap_axis_oarg_52_tstrb(ap_axis_oarg_52_tstrb),
        .ap_axis_oarg_52_tdata(ap_axis_oarg_52_tdata),
        .ap_axis_oarg_52_tready(ap_axis_oarg_52_tready),
        .m_axis_oarg_53_aclk(m_axis_oarg_53_aclk),
        .m_axis_oarg_53_aresetn(m_axis_oarg_53_aresetn),
        .m_axis_oarg_53_tlast(m_axis_oarg_53_tlast),
        .m_axis_oarg_53_tvalid(m_axis_oarg_53_tvalid),
        .m_axis_oarg_53_tkeep(m_axis_oarg_53_tkeep),
        .m_axis_oarg_53_tstrb(m_axis_oarg_53_tstrb),
        .m_axis_oarg_53_tdata(m_axis_oarg_53_tdata),
        .m_axis_oarg_53_tready(m_axis_oarg_53_tready),
        .ap_axis_oarg_53_tlast(ap_axis_oarg_53_tlast),
        .ap_axis_oarg_53_tvalid(ap_axis_oarg_53_tvalid),
        .ap_axis_oarg_53_tkeep(ap_axis_oarg_53_tkeep),
        .ap_axis_oarg_53_tstrb(ap_axis_oarg_53_tstrb),
        .ap_axis_oarg_53_tdata(ap_axis_oarg_53_tdata),
        .ap_axis_oarg_53_tready(ap_axis_oarg_53_tready),
        .m_axis_oarg_54_aclk(m_axis_oarg_54_aclk),
        .m_axis_oarg_54_aresetn(m_axis_oarg_54_aresetn),
        .m_axis_oarg_54_tlast(m_axis_oarg_54_tlast),
        .m_axis_oarg_54_tvalid(m_axis_oarg_54_tvalid),
        .m_axis_oarg_54_tkeep(m_axis_oarg_54_tkeep),
        .m_axis_oarg_54_tstrb(m_axis_oarg_54_tstrb),
        .m_axis_oarg_54_tdata(m_axis_oarg_54_tdata),
        .m_axis_oarg_54_tready(m_axis_oarg_54_tready),
        .ap_axis_oarg_54_tlast(ap_axis_oarg_54_tlast),
        .ap_axis_oarg_54_tvalid(ap_axis_oarg_54_tvalid),
        .ap_axis_oarg_54_tkeep(ap_axis_oarg_54_tkeep),
        .ap_axis_oarg_54_tstrb(ap_axis_oarg_54_tstrb),
        .ap_axis_oarg_54_tdata(ap_axis_oarg_54_tdata),
        .ap_axis_oarg_54_tready(ap_axis_oarg_54_tready),
        .m_axis_oarg_55_aclk(m_axis_oarg_55_aclk),
        .m_axis_oarg_55_aresetn(m_axis_oarg_55_aresetn),
        .m_axis_oarg_55_tlast(m_axis_oarg_55_tlast),
        .m_axis_oarg_55_tvalid(m_axis_oarg_55_tvalid),
        .m_axis_oarg_55_tkeep(m_axis_oarg_55_tkeep),
        .m_axis_oarg_55_tstrb(m_axis_oarg_55_tstrb),
        .m_axis_oarg_55_tdata(m_axis_oarg_55_tdata),
        .m_axis_oarg_55_tready(m_axis_oarg_55_tready),
        .ap_axis_oarg_55_tlast(ap_axis_oarg_55_tlast),
        .ap_axis_oarg_55_tvalid(ap_axis_oarg_55_tvalid),
        .ap_axis_oarg_55_tkeep(ap_axis_oarg_55_tkeep),
        .ap_axis_oarg_55_tstrb(ap_axis_oarg_55_tstrb),
        .ap_axis_oarg_55_tdata(ap_axis_oarg_55_tdata),
        .ap_axis_oarg_55_tready(ap_axis_oarg_55_tready),
        .m_axis_oarg_56_aclk(m_axis_oarg_56_aclk),
        .m_axis_oarg_56_aresetn(m_axis_oarg_56_aresetn),
        .m_axis_oarg_56_tlast(m_axis_oarg_56_tlast),
        .m_axis_oarg_56_tvalid(m_axis_oarg_56_tvalid),
        .m_axis_oarg_56_tkeep(m_axis_oarg_56_tkeep),
        .m_axis_oarg_56_tstrb(m_axis_oarg_56_tstrb),
        .m_axis_oarg_56_tdata(m_axis_oarg_56_tdata),
        .m_axis_oarg_56_tready(m_axis_oarg_56_tready),
        .ap_axis_oarg_56_tlast(ap_axis_oarg_56_tlast),
        .ap_axis_oarg_56_tvalid(ap_axis_oarg_56_tvalid),
        .ap_axis_oarg_56_tkeep(ap_axis_oarg_56_tkeep),
        .ap_axis_oarg_56_tstrb(ap_axis_oarg_56_tstrb),
        .ap_axis_oarg_56_tdata(ap_axis_oarg_56_tdata),
        .ap_axis_oarg_56_tready(ap_axis_oarg_56_tready),
        .m_axis_oarg_57_aclk(m_axis_oarg_57_aclk),
        .m_axis_oarg_57_aresetn(m_axis_oarg_57_aresetn),
        .m_axis_oarg_57_tlast(m_axis_oarg_57_tlast),
        .m_axis_oarg_57_tvalid(m_axis_oarg_57_tvalid),
        .m_axis_oarg_57_tkeep(m_axis_oarg_57_tkeep),
        .m_axis_oarg_57_tstrb(m_axis_oarg_57_tstrb),
        .m_axis_oarg_57_tdata(m_axis_oarg_57_tdata),
        .m_axis_oarg_57_tready(m_axis_oarg_57_tready),
        .ap_axis_oarg_57_tlast(ap_axis_oarg_57_tlast),
        .ap_axis_oarg_57_tvalid(ap_axis_oarg_57_tvalid),
        .ap_axis_oarg_57_tkeep(ap_axis_oarg_57_tkeep),
        .ap_axis_oarg_57_tstrb(ap_axis_oarg_57_tstrb),
        .ap_axis_oarg_57_tdata(ap_axis_oarg_57_tdata),
        .ap_axis_oarg_57_tready(ap_axis_oarg_57_tready),
        .m_axis_oarg_58_aclk(m_axis_oarg_58_aclk),
        .m_axis_oarg_58_aresetn(m_axis_oarg_58_aresetn),
        .m_axis_oarg_58_tlast(m_axis_oarg_58_tlast),
        .m_axis_oarg_58_tvalid(m_axis_oarg_58_tvalid),
        .m_axis_oarg_58_tkeep(m_axis_oarg_58_tkeep),
        .m_axis_oarg_58_tstrb(m_axis_oarg_58_tstrb),
        .m_axis_oarg_58_tdata(m_axis_oarg_58_tdata),
        .m_axis_oarg_58_tready(m_axis_oarg_58_tready),
        .ap_axis_oarg_58_tlast(ap_axis_oarg_58_tlast),
        .ap_axis_oarg_58_tvalid(ap_axis_oarg_58_tvalid),
        .ap_axis_oarg_58_tkeep(ap_axis_oarg_58_tkeep),
        .ap_axis_oarg_58_tstrb(ap_axis_oarg_58_tstrb),
        .ap_axis_oarg_58_tdata(ap_axis_oarg_58_tdata),
        .ap_axis_oarg_58_tready(ap_axis_oarg_58_tready),
        .m_axis_oarg_59_aclk(m_axis_oarg_59_aclk),
        .m_axis_oarg_59_aresetn(m_axis_oarg_59_aresetn),
        .m_axis_oarg_59_tlast(m_axis_oarg_59_tlast),
        .m_axis_oarg_59_tvalid(m_axis_oarg_59_tvalid),
        .m_axis_oarg_59_tkeep(m_axis_oarg_59_tkeep),
        .m_axis_oarg_59_tstrb(m_axis_oarg_59_tstrb),
        .m_axis_oarg_59_tdata(m_axis_oarg_59_tdata),
        .m_axis_oarg_59_tready(m_axis_oarg_59_tready),
        .ap_axis_oarg_59_tlast(ap_axis_oarg_59_tlast),
        .ap_axis_oarg_59_tvalid(ap_axis_oarg_59_tvalid),
        .ap_axis_oarg_59_tkeep(ap_axis_oarg_59_tkeep),
        .ap_axis_oarg_59_tstrb(ap_axis_oarg_59_tstrb),
        .ap_axis_oarg_59_tdata(ap_axis_oarg_59_tdata),
        .ap_axis_oarg_59_tready(ap_axis_oarg_59_tready),
        .m_axis_oarg_60_aclk(m_axis_oarg_60_aclk),
        .m_axis_oarg_60_aresetn(m_axis_oarg_60_aresetn),
        .m_axis_oarg_60_tlast(m_axis_oarg_60_tlast),
        .m_axis_oarg_60_tvalid(m_axis_oarg_60_tvalid),
        .m_axis_oarg_60_tkeep(m_axis_oarg_60_tkeep),
        .m_axis_oarg_60_tstrb(m_axis_oarg_60_tstrb),
        .m_axis_oarg_60_tdata(m_axis_oarg_60_tdata),
        .m_axis_oarg_60_tready(m_axis_oarg_60_tready),
        .ap_axis_oarg_60_tlast(ap_axis_oarg_60_tlast),
        .ap_axis_oarg_60_tvalid(ap_axis_oarg_60_tvalid),
        .ap_axis_oarg_60_tkeep(ap_axis_oarg_60_tkeep),
        .ap_axis_oarg_60_tstrb(ap_axis_oarg_60_tstrb),
        .ap_axis_oarg_60_tdata(ap_axis_oarg_60_tdata),
        .ap_axis_oarg_60_tready(ap_axis_oarg_60_tready),
        .m_axis_oarg_61_aclk(m_axis_oarg_61_aclk),
        .m_axis_oarg_61_aresetn(m_axis_oarg_61_aresetn),
        .m_axis_oarg_61_tlast(m_axis_oarg_61_tlast),
        .m_axis_oarg_61_tvalid(m_axis_oarg_61_tvalid),
        .m_axis_oarg_61_tkeep(m_axis_oarg_61_tkeep),
        .m_axis_oarg_61_tstrb(m_axis_oarg_61_tstrb),
        .m_axis_oarg_61_tdata(m_axis_oarg_61_tdata),
        .m_axis_oarg_61_tready(m_axis_oarg_61_tready),
        .ap_axis_oarg_61_tlast(ap_axis_oarg_61_tlast),
        .ap_axis_oarg_61_tvalid(ap_axis_oarg_61_tvalid),
        .ap_axis_oarg_61_tkeep(ap_axis_oarg_61_tkeep),
        .ap_axis_oarg_61_tstrb(ap_axis_oarg_61_tstrb),
        .ap_axis_oarg_61_tdata(ap_axis_oarg_61_tdata),
        .ap_axis_oarg_61_tready(ap_axis_oarg_61_tready),
        .m_axis_oarg_62_aclk(m_axis_oarg_62_aclk),
        .m_axis_oarg_62_aresetn(m_axis_oarg_62_aresetn),
        .m_axis_oarg_62_tlast(m_axis_oarg_62_tlast),
        .m_axis_oarg_62_tvalid(m_axis_oarg_62_tvalid),
        .m_axis_oarg_62_tkeep(m_axis_oarg_62_tkeep),
        .m_axis_oarg_62_tstrb(m_axis_oarg_62_tstrb),
        .m_axis_oarg_62_tdata(m_axis_oarg_62_tdata),
        .m_axis_oarg_62_tready(m_axis_oarg_62_tready),
        .ap_axis_oarg_62_tlast(ap_axis_oarg_62_tlast),
        .ap_axis_oarg_62_tvalid(ap_axis_oarg_62_tvalid),
        .ap_axis_oarg_62_tkeep(ap_axis_oarg_62_tkeep),
        .ap_axis_oarg_62_tstrb(ap_axis_oarg_62_tstrb),
        .ap_axis_oarg_62_tdata(ap_axis_oarg_62_tdata),
        .ap_axis_oarg_62_tready(ap_axis_oarg_62_tready),
        .m_axis_oarg_63_aclk(m_axis_oarg_63_aclk),
        .m_axis_oarg_63_aresetn(m_axis_oarg_63_aresetn),
        .m_axis_oarg_63_tlast(m_axis_oarg_63_tlast),
        .m_axis_oarg_63_tvalid(m_axis_oarg_63_tvalid),
        .m_axis_oarg_63_tkeep(m_axis_oarg_63_tkeep),
        .m_axis_oarg_63_tstrb(m_axis_oarg_63_tstrb),
        .m_axis_oarg_63_tdata(m_axis_oarg_63_tdata),
        .m_axis_oarg_63_tready(m_axis_oarg_63_tready),
        .ap_axis_oarg_63_tlast(ap_axis_oarg_63_tlast),
        .ap_axis_oarg_63_tvalid(ap_axis_oarg_63_tvalid),
        .ap_axis_oarg_63_tkeep(ap_axis_oarg_63_tkeep),
        .ap_axis_oarg_63_tstrb(ap_axis_oarg_63_tstrb),
        .ap_axis_oarg_63_tdata(ap_axis_oarg_63_tdata),
        .ap_axis_oarg_63_tready(ap_axis_oarg_63_tready),
        .m_axis_oarg_64_aclk(m_axis_oarg_64_aclk),
        .m_axis_oarg_64_aresetn(m_axis_oarg_64_aresetn),
        .m_axis_oarg_64_tlast(m_axis_oarg_64_tlast),
        .m_axis_oarg_64_tvalid(m_axis_oarg_64_tvalid),
        .m_axis_oarg_64_tkeep(m_axis_oarg_64_tkeep),
        .m_axis_oarg_64_tstrb(m_axis_oarg_64_tstrb),
        .m_axis_oarg_64_tdata(m_axis_oarg_64_tdata),
        .m_axis_oarg_64_tready(m_axis_oarg_64_tready),
        .ap_axis_oarg_64_tlast(ap_axis_oarg_64_tlast),
        .ap_axis_oarg_64_tvalid(ap_axis_oarg_64_tvalid),
        .ap_axis_oarg_64_tkeep(ap_axis_oarg_64_tkeep),
        .ap_axis_oarg_64_tstrb(ap_axis_oarg_64_tstrb),
        .ap_axis_oarg_64_tdata(ap_axis_oarg_64_tdata),
        .ap_axis_oarg_64_tready(ap_axis_oarg_64_tready),
        .m_axis_oarg_65_aclk(m_axis_oarg_65_aclk),
        .m_axis_oarg_65_aresetn(m_axis_oarg_65_aresetn),
        .m_axis_oarg_65_tlast(m_axis_oarg_65_tlast),
        .m_axis_oarg_65_tvalid(m_axis_oarg_65_tvalid),
        .m_axis_oarg_65_tkeep(m_axis_oarg_65_tkeep),
        .m_axis_oarg_65_tstrb(m_axis_oarg_65_tstrb),
        .m_axis_oarg_65_tdata(m_axis_oarg_65_tdata),
        .m_axis_oarg_65_tready(m_axis_oarg_65_tready),
        .ap_axis_oarg_65_tlast(ap_axis_oarg_65_tlast),
        .ap_axis_oarg_65_tvalid(ap_axis_oarg_65_tvalid),
        .ap_axis_oarg_65_tkeep(ap_axis_oarg_65_tkeep),
        .ap_axis_oarg_65_tstrb(ap_axis_oarg_65_tstrb),
        .ap_axis_oarg_65_tdata(ap_axis_oarg_65_tdata),
        .ap_axis_oarg_65_tready(ap_axis_oarg_65_tready),
        .m_axis_oarg_66_aclk(m_axis_oarg_66_aclk),
        .m_axis_oarg_66_aresetn(m_axis_oarg_66_aresetn),
        .m_axis_oarg_66_tlast(m_axis_oarg_66_tlast),
        .m_axis_oarg_66_tvalid(m_axis_oarg_66_tvalid),
        .m_axis_oarg_66_tkeep(m_axis_oarg_66_tkeep),
        .m_axis_oarg_66_tstrb(m_axis_oarg_66_tstrb),
        .m_axis_oarg_66_tdata(m_axis_oarg_66_tdata),
        .m_axis_oarg_66_tready(m_axis_oarg_66_tready),
        .ap_axis_oarg_66_tlast(ap_axis_oarg_66_tlast),
        .ap_axis_oarg_66_tvalid(ap_axis_oarg_66_tvalid),
        .ap_axis_oarg_66_tkeep(ap_axis_oarg_66_tkeep),
        .ap_axis_oarg_66_tstrb(ap_axis_oarg_66_tstrb),
        .ap_axis_oarg_66_tdata(ap_axis_oarg_66_tdata),
        .ap_axis_oarg_66_tready(ap_axis_oarg_66_tready),
        .m_axis_oarg_67_aclk(m_axis_oarg_67_aclk),
        .m_axis_oarg_67_aresetn(m_axis_oarg_67_aresetn),
        .m_axis_oarg_67_tlast(m_axis_oarg_67_tlast),
        .m_axis_oarg_67_tvalid(m_axis_oarg_67_tvalid),
        .m_axis_oarg_67_tkeep(m_axis_oarg_67_tkeep),
        .m_axis_oarg_67_tstrb(m_axis_oarg_67_tstrb),
        .m_axis_oarg_67_tdata(m_axis_oarg_67_tdata),
        .m_axis_oarg_67_tready(m_axis_oarg_67_tready),
        .ap_axis_oarg_67_tlast(ap_axis_oarg_67_tlast),
        .ap_axis_oarg_67_tvalid(ap_axis_oarg_67_tvalid),
        .ap_axis_oarg_67_tkeep(ap_axis_oarg_67_tkeep),
        .ap_axis_oarg_67_tstrb(ap_axis_oarg_67_tstrb),
        .ap_axis_oarg_67_tdata(ap_axis_oarg_67_tdata),
        .ap_axis_oarg_67_tready(ap_axis_oarg_67_tready),
        .m_axis_oarg_68_aclk(m_axis_oarg_68_aclk),
        .m_axis_oarg_68_aresetn(m_axis_oarg_68_aresetn),
        .m_axis_oarg_68_tlast(m_axis_oarg_68_tlast),
        .m_axis_oarg_68_tvalid(m_axis_oarg_68_tvalid),
        .m_axis_oarg_68_tkeep(m_axis_oarg_68_tkeep),
        .m_axis_oarg_68_tstrb(m_axis_oarg_68_tstrb),
        .m_axis_oarg_68_tdata(m_axis_oarg_68_tdata),
        .m_axis_oarg_68_tready(m_axis_oarg_68_tready),
        .ap_axis_oarg_68_tlast(ap_axis_oarg_68_tlast),
        .ap_axis_oarg_68_tvalid(ap_axis_oarg_68_tvalid),
        .ap_axis_oarg_68_tkeep(ap_axis_oarg_68_tkeep),
        .ap_axis_oarg_68_tstrb(ap_axis_oarg_68_tstrb),
        .ap_axis_oarg_68_tdata(ap_axis_oarg_68_tdata),
        .ap_axis_oarg_68_tready(ap_axis_oarg_68_tready),
        .m_axis_oarg_69_aclk(m_axis_oarg_69_aclk),
        .m_axis_oarg_69_aresetn(m_axis_oarg_69_aresetn),
        .m_axis_oarg_69_tlast(m_axis_oarg_69_tlast),
        .m_axis_oarg_69_tvalid(m_axis_oarg_69_tvalid),
        .m_axis_oarg_69_tkeep(m_axis_oarg_69_tkeep),
        .m_axis_oarg_69_tstrb(m_axis_oarg_69_tstrb),
        .m_axis_oarg_69_tdata(m_axis_oarg_69_tdata),
        .m_axis_oarg_69_tready(m_axis_oarg_69_tready),
        .ap_axis_oarg_69_tlast(ap_axis_oarg_69_tlast),
        .ap_axis_oarg_69_tvalid(ap_axis_oarg_69_tvalid),
        .ap_axis_oarg_69_tkeep(ap_axis_oarg_69_tkeep),
        .ap_axis_oarg_69_tstrb(ap_axis_oarg_69_tstrb),
        .ap_axis_oarg_69_tdata(ap_axis_oarg_69_tdata),
        .ap_axis_oarg_69_tready(ap_axis_oarg_69_tready),
        .m_axis_oarg_70_aclk(m_axis_oarg_70_aclk),
        .m_axis_oarg_70_aresetn(m_axis_oarg_70_aresetn),
        .m_axis_oarg_70_tlast(m_axis_oarg_70_tlast),
        .m_axis_oarg_70_tvalid(m_axis_oarg_70_tvalid),
        .m_axis_oarg_70_tkeep(m_axis_oarg_70_tkeep),
        .m_axis_oarg_70_tstrb(m_axis_oarg_70_tstrb),
        .m_axis_oarg_70_tdata(m_axis_oarg_70_tdata),
        .m_axis_oarg_70_tready(m_axis_oarg_70_tready),
        .ap_axis_oarg_70_tlast(ap_axis_oarg_70_tlast),
        .ap_axis_oarg_70_tvalid(ap_axis_oarg_70_tvalid),
        .ap_axis_oarg_70_tkeep(ap_axis_oarg_70_tkeep),
        .ap_axis_oarg_70_tstrb(ap_axis_oarg_70_tstrb),
        .ap_axis_oarg_70_tdata(ap_axis_oarg_70_tdata),
        .ap_axis_oarg_70_tready(ap_axis_oarg_70_tready),
        .m_axis_oarg_71_aclk(m_axis_oarg_71_aclk),
        .m_axis_oarg_71_aresetn(m_axis_oarg_71_aresetn),
        .m_axis_oarg_71_tlast(m_axis_oarg_71_tlast),
        .m_axis_oarg_71_tvalid(m_axis_oarg_71_tvalid),
        .m_axis_oarg_71_tkeep(m_axis_oarg_71_tkeep),
        .m_axis_oarg_71_tstrb(m_axis_oarg_71_tstrb),
        .m_axis_oarg_71_tdata(m_axis_oarg_71_tdata),
        .m_axis_oarg_71_tready(m_axis_oarg_71_tready),
        .ap_axis_oarg_71_tlast(ap_axis_oarg_71_tlast),
        .ap_axis_oarg_71_tvalid(ap_axis_oarg_71_tvalid),
        .ap_axis_oarg_71_tkeep(ap_axis_oarg_71_tkeep),
        .ap_axis_oarg_71_tstrb(ap_axis_oarg_71_tstrb),
        .ap_axis_oarg_71_tdata(ap_axis_oarg_71_tdata),
        .ap_axis_oarg_71_tready(ap_axis_oarg_71_tready),
        .m_axis_oarg_72_aclk(m_axis_oarg_72_aclk),
        .m_axis_oarg_72_aresetn(m_axis_oarg_72_aresetn),
        .m_axis_oarg_72_tlast(m_axis_oarg_72_tlast),
        .m_axis_oarg_72_tvalid(m_axis_oarg_72_tvalid),
        .m_axis_oarg_72_tkeep(m_axis_oarg_72_tkeep),
        .m_axis_oarg_72_tstrb(m_axis_oarg_72_tstrb),
        .m_axis_oarg_72_tdata(m_axis_oarg_72_tdata),
        .m_axis_oarg_72_tready(m_axis_oarg_72_tready),
        .ap_axis_oarg_72_tlast(ap_axis_oarg_72_tlast),
        .ap_axis_oarg_72_tvalid(ap_axis_oarg_72_tvalid),
        .ap_axis_oarg_72_tkeep(ap_axis_oarg_72_tkeep),
        .ap_axis_oarg_72_tstrb(ap_axis_oarg_72_tstrb),
        .ap_axis_oarg_72_tdata(ap_axis_oarg_72_tdata),
        .ap_axis_oarg_72_tready(ap_axis_oarg_72_tready),
        .m_axis_oarg_73_aclk(m_axis_oarg_73_aclk),
        .m_axis_oarg_73_aresetn(m_axis_oarg_73_aresetn),
        .m_axis_oarg_73_tlast(m_axis_oarg_73_tlast),
        .m_axis_oarg_73_tvalid(m_axis_oarg_73_tvalid),
        .m_axis_oarg_73_tkeep(m_axis_oarg_73_tkeep),
        .m_axis_oarg_73_tstrb(m_axis_oarg_73_tstrb),
        .m_axis_oarg_73_tdata(m_axis_oarg_73_tdata),
        .m_axis_oarg_73_tready(m_axis_oarg_73_tready),
        .ap_axis_oarg_73_tlast(ap_axis_oarg_73_tlast),
        .ap_axis_oarg_73_tvalid(ap_axis_oarg_73_tvalid),
        .ap_axis_oarg_73_tkeep(ap_axis_oarg_73_tkeep),
        .ap_axis_oarg_73_tstrb(ap_axis_oarg_73_tstrb),
        .ap_axis_oarg_73_tdata(ap_axis_oarg_73_tdata),
        .ap_axis_oarg_73_tready(ap_axis_oarg_73_tready),
        .m_axis_oarg_74_aclk(m_axis_oarg_74_aclk),
        .m_axis_oarg_74_aresetn(m_axis_oarg_74_aresetn),
        .m_axis_oarg_74_tlast(m_axis_oarg_74_tlast),
        .m_axis_oarg_74_tvalid(m_axis_oarg_74_tvalid),
        .m_axis_oarg_74_tkeep(m_axis_oarg_74_tkeep),
        .m_axis_oarg_74_tstrb(m_axis_oarg_74_tstrb),
        .m_axis_oarg_74_tdata(m_axis_oarg_74_tdata),
        .m_axis_oarg_74_tready(m_axis_oarg_74_tready),
        .ap_axis_oarg_74_tlast(ap_axis_oarg_74_tlast),
        .ap_axis_oarg_74_tvalid(ap_axis_oarg_74_tvalid),
        .ap_axis_oarg_74_tkeep(ap_axis_oarg_74_tkeep),
        .ap_axis_oarg_74_tstrb(ap_axis_oarg_74_tstrb),
        .ap_axis_oarg_74_tdata(ap_axis_oarg_74_tdata),
        .ap_axis_oarg_74_tready(ap_axis_oarg_74_tready),
        .m_axis_oarg_75_aclk(m_axis_oarg_75_aclk),
        .m_axis_oarg_75_aresetn(m_axis_oarg_75_aresetn),
        .m_axis_oarg_75_tlast(m_axis_oarg_75_tlast),
        .m_axis_oarg_75_tvalid(m_axis_oarg_75_tvalid),
        .m_axis_oarg_75_tkeep(m_axis_oarg_75_tkeep),
        .m_axis_oarg_75_tstrb(m_axis_oarg_75_tstrb),
        .m_axis_oarg_75_tdata(m_axis_oarg_75_tdata),
        .m_axis_oarg_75_tready(m_axis_oarg_75_tready),
        .ap_axis_oarg_75_tlast(ap_axis_oarg_75_tlast),
        .ap_axis_oarg_75_tvalid(ap_axis_oarg_75_tvalid),
        .ap_axis_oarg_75_tkeep(ap_axis_oarg_75_tkeep),
        .ap_axis_oarg_75_tstrb(ap_axis_oarg_75_tstrb),
        .ap_axis_oarg_75_tdata(ap_axis_oarg_75_tdata),
        .ap_axis_oarg_75_tready(ap_axis_oarg_75_tready),
        .m_axis_oarg_76_aclk(m_axis_oarg_76_aclk),
        .m_axis_oarg_76_aresetn(m_axis_oarg_76_aresetn),
        .m_axis_oarg_76_tlast(m_axis_oarg_76_tlast),
        .m_axis_oarg_76_tvalid(m_axis_oarg_76_tvalid),
        .m_axis_oarg_76_tkeep(m_axis_oarg_76_tkeep),
        .m_axis_oarg_76_tstrb(m_axis_oarg_76_tstrb),
        .m_axis_oarg_76_tdata(m_axis_oarg_76_tdata),
        .m_axis_oarg_76_tready(m_axis_oarg_76_tready),
        .ap_axis_oarg_76_tlast(ap_axis_oarg_76_tlast),
        .ap_axis_oarg_76_tvalid(ap_axis_oarg_76_tvalid),
        .ap_axis_oarg_76_tkeep(ap_axis_oarg_76_tkeep),
        .ap_axis_oarg_76_tstrb(ap_axis_oarg_76_tstrb),
        .ap_axis_oarg_76_tdata(ap_axis_oarg_76_tdata),
        .ap_axis_oarg_76_tready(ap_axis_oarg_76_tready),
        .m_axis_oarg_77_aclk(m_axis_oarg_77_aclk),
        .m_axis_oarg_77_aresetn(m_axis_oarg_77_aresetn),
        .m_axis_oarg_77_tlast(m_axis_oarg_77_tlast),
        .m_axis_oarg_77_tvalid(m_axis_oarg_77_tvalid),
        .m_axis_oarg_77_tkeep(m_axis_oarg_77_tkeep),
        .m_axis_oarg_77_tstrb(m_axis_oarg_77_tstrb),
        .m_axis_oarg_77_tdata(m_axis_oarg_77_tdata),
        .m_axis_oarg_77_tready(m_axis_oarg_77_tready),
        .ap_axis_oarg_77_tlast(ap_axis_oarg_77_tlast),
        .ap_axis_oarg_77_tvalid(ap_axis_oarg_77_tvalid),
        .ap_axis_oarg_77_tkeep(ap_axis_oarg_77_tkeep),
        .ap_axis_oarg_77_tstrb(ap_axis_oarg_77_tstrb),
        .ap_axis_oarg_77_tdata(ap_axis_oarg_77_tdata),
        .ap_axis_oarg_77_tready(ap_axis_oarg_77_tready),
        .m_axis_oarg_78_aclk(m_axis_oarg_78_aclk),
        .m_axis_oarg_78_aresetn(m_axis_oarg_78_aresetn),
        .m_axis_oarg_78_tlast(m_axis_oarg_78_tlast),
        .m_axis_oarg_78_tvalid(m_axis_oarg_78_tvalid),
        .m_axis_oarg_78_tkeep(m_axis_oarg_78_tkeep),
        .m_axis_oarg_78_tstrb(m_axis_oarg_78_tstrb),
        .m_axis_oarg_78_tdata(m_axis_oarg_78_tdata),
        .m_axis_oarg_78_tready(m_axis_oarg_78_tready),
        .ap_axis_oarg_78_tlast(ap_axis_oarg_78_tlast),
        .ap_axis_oarg_78_tvalid(ap_axis_oarg_78_tvalid),
        .ap_axis_oarg_78_tkeep(ap_axis_oarg_78_tkeep),
        .ap_axis_oarg_78_tstrb(ap_axis_oarg_78_tstrb),
        .ap_axis_oarg_78_tdata(ap_axis_oarg_78_tdata),
        .ap_axis_oarg_78_tready(ap_axis_oarg_78_tready),
        .m_axis_oarg_79_aclk(m_axis_oarg_79_aclk),
        .m_axis_oarg_79_aresetn(m_axis_oarg_79_aresetn),
        .m_axis_oarg_79_tlast(m_axis_oarg_79_tlast),
        .m_axis_oarg_79_tvalid(m_axis_oarg_79_tvalid),
        .m_axis_oarg_79_tkeep(m_axis_oarg_79_tkeep),
        .m_axis_oarg_79_tstrb(m_axis_oarg_79_tstrb),
        .m_axis_oarg_79_tdata(m_axis_oarg_79_tdata),
        .m_axis_oarg_79_tready(m_axis_oarg_79_tready),
        .ap_axis_oarg_79_tlast(ap_axis_oarg_79_tlast),
        .ap_axis_oarg_79_tvalid(ap_axis_oarg_79_tvalid),
        .ap_axis_oarg_79_tkeep(ap_axis_oarg_79_tkeep),
        .ap_axis_oarg_79_tstrb(ap_axis_oarg_79_tstrb),
        .ap_axis_oarg_79_tdata(ap_axis_oarg_79_tdata),
        .ap_axis_oarg_79_tready(ap_axis_oarg_79_tready),
        .m_axis_oarg_80_aclk(m_axis_oarg_80_aclk),
        .m_axis_oarg_80_aresetn(m_axis_oarg_80_aresetn),
        .m_axis_oarg_80_tlast(m_axis_oarg_80_tlast),
        .m_axis_oarg_80_tvalid(m_axis_oarg_80_tvalid),
        .m_axis_oarg_80_tkeep(m_axis_oarg_80_tkeep),
        .m_axis_oarg_80_tstrb(m_axis_oarg_80_tstrb),
        .m_axis_oarg_80_tdata(m_axis_oarg_80_tdata),
        .m_axis_oarg_80_tready(m_axis_oarg_80_tready),
        .ap_axis_oarg_80_tlast(ap_axis_oarg_80_tlast),
        .ap_axis_oarg_80_tvalid(ap_axis_oarg_80_tvalid),
        .ap_axis_oarg_80_tkeep(ap_axis_oarg_80_tkeep),
        .ap_axis_oarg_80_tstrb(ap_axis_oarg_80_tstrb),
        .ap_axis_oarg_80_tdata(ap_axis_oarg_80_tdata),
        .ap_axis_oarg_80_tready(ap_axis_oarg_80_tready),
        .m_axis_oarg_81_aclk(m_axis_oarg_81_aclk),
        .m_axis_oarg_81_aresetn(m_axis_oarg_81_aresetn),
        .m_axis_oarg_81_tlast(m_axis_oarg_81_tlast),
        .m_axis_oarg_81_tvalid(m_axis_oarg_81_tvalid),
        .m_axis_oarg_81_tkeep(m_axis_oarg_81_tkeep),
        .m_axis_oarg_81_tstrb(m_axis_oarg_81_tstrb),
        .m_axis_oarg_81_tdata(m_axis_oarg_81_tdata),
        .m_axis_oarg_81_tready(m_axis_oarg_81_tready),
        .ap_axis_oarg_81_tlast(ap_axis_oarg_81_tlast),
        .ap_axis_oarg_81_tvalid(ap_axis_oarg_81_tvalid),
        .ap_axis_oarg_81_tkeep(ap_axis_oarg_81_tkeep),
        .ap_axis_oarg_81_tstrb(ap_axis_oarg_81_tstrb),
        .ap_axis_oarg_81_tdata(ap_axis_oarg_81_tdata),
        .ap_axis_oarg_81_tready(ap_axis_oarg_81_tready),
        .m_axis_oarg_82_aclk(m_axis_oarg_82_aclk),
        .m_axis_oarg_82_aresetn(m_axis_oarg_82_aresetn),
        .m_axis_oarg_82_tlast(m_axis_oarg_82_tlast),
        .m_axis_oarg_82_tvalid(m_axis_oarg_82_tvalid),
        .m_axis_oarg_82_tkeep(m_axis_oarg_82_tkeep),
        .m_axis_oarg_82_tstrb(m_axis_oarg_82_tstrb),
        .m_axis_oarg_82_tdata(m_axis_oarg_82_tdata),
        .m_axis_oarg_82_tready(m_axis_oarg_82_tready),
        .ap_axis_oarg_82_tlast(ap_axis_oarg_82_tlast),
        .ap_axis_oarg_82_tvalid(ap_axis_oarg_82_tvalid),
        .ap_axis_oarg_82_tkeep(ap_axis_oarg_82_tkeep),
        .ap_axis_oarg_82_tstrb(ap_axis_oarg_82_tstrb),
        .ap_axis_oarg_82_tdata(ap_axis_oarg_82_tdata),
        .ap_axis_oarg_82_tready(ap_axis_oarg_82_tready),
        .m_axis_oarg_83_aclk(m_axis_oarg_83_aclk),
        .m_axis_oarg_83_aresetn(m_axis_oarg_83_aresetn),
        .m_axis_oarg_83_tlast(m_axis_oarg_83_tlast),
        .m_axis_oarg_83_tvalid(m_axis_oarg_83_tvalid),
        .m_axis_oarg_83_tkeep(m_axis_oarg_83_tkeep),
        .m_axis_oarg_83_tstrb(m_axis_oarg_83_tstrb),
        .m_axis_oarg_83_tdata(m_axis_oarg_83_tdata),
        .m_axis_oarg_83_tready(m_axis_oarg_83_tready),
        .ap_axis_oarg_83_tlast(ap_axis_oarg_83_tlast),
        .ap_axis_oarg_83_tvalid(ap_axis_oarg_83_tvalid),
        .ap_axis_oarg_83_tkeep(ap_axis_oarg_83_tkeep),
        .ap_axis_oarg_83_tstrb(ap_axis_oarg_83_tstrb),
        .ap_axis_oarg_83_tdata(ap_axis_oarg_83_tdata),
        .ap_axis_oarg_83_tready(ap_axis_oarg_83_tready),
        .m_axis_oarg_84_aclk(m_axis_oarg_84_aclk),
        .m_axis_oarg_84_aresetn(m_axis_oarg_84_aresetn),
        .m_axis_oarg_84_tlast(m_axis_oarg_84_tlast),
        .m_axis_oarg_84_tvalid(m_axis_oarg_84_tvalid),
        .m_axis_oarg_84_tkeep(m_axis_oarg_84_tkeep),
        .m_axis_oarg_84_tstrb(m_axis_oarg_84_tstrb),
        .m_axis_oarg_84_tdata(m_axis_oarg_84_tdata),
        .m_axis_oarg_84_tready(m_axis_oarg_84_tready),
        .ap_axis_oarg_84_tlast(ap_axis_oarg_84_tlast),
        .ap_axis_oarg_84_tvalid(ap_axis_oarg_84_tvalid),
        .ap_axis_oarg_84_tkeep(ap_axis_oarg_84_tkeep),
        .ap_axis_oarg_84_tstrb(ap_axis_oarg_84_tstrb),
        .ap_axis_oarg_84_tdata(ap_axis_oarg_84_tdata),
        .ap_axis_oarg_84_tready(ap_axis_oarg_84_tready),
        .m_axis_oarg_85_aclk(m_axis_oarg_85_aclk),
        .m_axis_oarg_85_aresetn(m_axis_oarg_85_aresetn),
        .m_axis_oarg_85_tlast(m_axis_oarg_85_tlast),
        .m_axis_oarg_85_tvalid(m_axis_oarg_85_tvalid),
        .m_axis_oarg_85_tkeep(m_axis_oarg_85_tkeep),
        .m_axis_oarg_85_tstrb(m_axis_oarg_85_tstrb),
        .m_axis_oarg_85_tdata(m_axis_oarg_85_tdata),
        .m_axis_oarg_85_tready(m_axis_oarg_85_tready),
        .ap_axis_oarg_85_tlast(ap_axis_oarg_85_tlast),
        .ap_axis_oarg_85_tvalid(ap_axis_oarg_85_tvalid),
        .ap_axis_oarg_85_tkeep(ap_axis_oarg_85_tkeep),
        .ap_axis_oarg_85_tstrb(ap_axis_oarg_85_tstrb),
        .ap_axis_oarg_85_tdata(ap_axis_oarg_85_tdata),
        .ap_axis_oarg_85_tready(ap_axis_oarg_85_tready),
        .m_axis_oarg_86_aclk(m_axis_oarg_86_aclk),
        .m_axis_oarg_86_aresetn(m_axis_oarg_86_aresetn),
        .m_axis_oarg_86_tlast(m_axis_oarg_86_tlast),
        .m_axis_oarg_86_tvalid(m_axis_oarg_86_tvalid),
        .m_axis_oarg_86_tkeep(m_axis_oarg_86_tkeep),
        .m_axis_oarg_86_tstrb(m_axis_oarg_86_tstrb),
        .m_axis_oarg_86_tdata(m_axis_oarg_86_tdata),
        .m_axis_oarg_86_tready(m_axis_oarg_86_tready),
        .ap_axis_oarg_86_tlast(ap_axis_oarg_86_tlast),
        .ap_axis_oarg_86_tvalid(ap_axis_oarg_86_tvalid),
        .ap_axis_oarg_86_tkeep(ap_axis_oarg_86_tkeep),
        .ap_axis_oarg_86_tstrb(ap_axis_oarg_86_tstrb),
        .ap_axis_oarg_86_tdata(ap_axis_oarg_86_tdata),
        .ap_axis_oarg_86_tready(ap_axis_oarg_86_tready),
        .m_axis_oarg_87_aclk(m_axis_oarg_87_aclk),
        .m_axis_oarg_87_aresetn(m_axis_oarg_87_aresetn),
        .m_axis_oarg_87_tlast(m_axis_oarg_87_tlast),
        .m_axis_oarg_87_tvalid(m_axis_oarg_87_tvalid),
        .m_axis_oarg_87_tkeep(m_axis_oarg_87_tkeep),
        .m_axis_oarg_87_tstrb(m_axis_oarg_87_tstrb),
        .m_axis_oarg_87_tdata(m_axis_oarg_87_tdata),
        .m_axis_oarg_87_tready(m_axis_oarg_87_tready),
        .ap_axis_oarg_87_tlast(ap_axis_oarg_87_tlast),
        .ap_axis_oarg_87_tvalid(ap_axis_oarg_87_tvalid),
        .ap_axis_oarg_87_tkeep(ap_axis_oarg_87_tkeep),
        .ap_axis_oarg_87_tstrb(ap_axis_oarg_87_tstrb),
        .ap_axis_oarg_87_tdata(ap_axis_oarg_87_tdata),
        .ap_axis_oarg_87_tready(ap_axis_oarg_87_tready),
        .m_axis_oarg_88_aclk(m_axis_oarg_88_aclk),
        .m_axis_oarg_88_aresetn(m_axis_oarg_88_aresetn),
        .m_axis_oarg_88_tlast(m_axis_oarg_88_tlast),
        .m_axis_oarg_88_tvalid(m_axis_oarg_88_tvalid),
        .m_axis_oarg_88_tkeep(m_axis_oarg_88_tkeep),
        .m_axis_oarg_88_tstrb(m_axis_oarg_88_tstrb),
        .m_axis_oarg_88_tdata(m_axis_oarg_88_tdata),
        .m_axis_oarg_88_tready(m_axis_oarg_88_tready),
        .ap_axis_oarg_88_tlast(ap_axis_oarg_88_tlast),
        .ap_axis_oarg_88_tvalid(ap_axis_oarg_88_tvalid),
        .ap_axis_oarg_88_tkeep(ap_axis_oarg_88_tkeep),
        .ap_axis_oarg_88_tstrb(ap_axis_oarg_88_tstrb),
        .ap_axis_oarg_88_tdata(ap_axis_oarg_88_tdata),
        .ap_axis_oarg_88_tready(ap_axis_oarg_88_tready),
        .m_axis_oarg_89_aclk(m_axis_oarg_89_aclk),
        .m_axis_oarg_89_aresetn(m_axis_oarg_89_aresetn),
        .m_axis_oarg_89_tlast(m_axis_oarg_89_tlast),
        .m_axis_oarg_89_tvalid(m_axis_oarg_89_tvalid),
        .m_axis_oarg_89_tkeep(m_axis_oarg_89_tkeep),
        .m_axis_oarg_89_tstrb(m_axis_oarg_89_tstrb),
        .m_axis_oarg_89_tdata(m_axis_oarg_89_tdata),
        .m_axis_oarg_89_tready(m_axis_oarg_89_tready),
        .ap_axis_oarg_89_tlast(ap_axis_oarg_89_tlast),
        .ap_axis_oarg_89_tvalid(ap_axis_oarg_89_tvalid),
        .ap_axis_oarg_89_tkeep(ap_axis_oarg_89_tkeep),
        .ap_axis_oarg_89_tstrb(ap_axis_oarg_89_tstrb),
        .ap_axis_oarg_89_tdata(ap_axis_oarg_89_tdata),
        .ap_axis_oarg_89_tready(ap_axis_oarg_89_tready),
        .m_axis_oarg_90_aclk(m_axis_oarg_90_aclk),
        .m_axis_oarg_90_aresetn(m_axis_oarg_90_aresetn),
        .m_axis_oarg_90_tlast(m_axis_oarg_90_tlast),
        .m_axis_oarg_90_tvalid(m_axis_oarg_90_tvalid),
        .m_axis_oarg_90_tkeep(m_axis_oarg_90_tkeep),
        .m_axis_oarg_90_tstrb(m_axis_oarg_90_tstrb),
        .m_axis_oarg_90_tdata(m_axis_oarg_90_tdata),
        .m_axis_oarg_90_tready(m_axis_oarg_90_tready),
        .ap_axis_oarg_90_tlast(ap_axis_oarg_90_tlast),
        .ap_axis_oarg_90_tvalid(ap_axis_oarg_90_tvalid),
        .ap_axis_oarg_90_tkeep(ap_axis_oarg_90_tkeep),
        .ap_axis_oarg_90_tstrb(ap_axis_oarg_90_tstrb),
        .ap_axis_oarg_90_tdata(ap_axis_oarg_90_tdata),
        .ap_axis_oarg_90_tready(ap_axis_oarg_90_tready),
        .m_axis_oarg_91_aclk(m_axis_oarg_91_aclk),
        .m_axis_oarg_91_aresetn(m_axis_oarg_91_aresetn),
        .m_axis_oarg_91_tlast(m_axis_oarg_91_tlast),
        .m_axis_oarg_91_tvalid(m_axis_oarg_91_tvalid),
        .m_axis_oarg_91_tkeep(m_axis_oarg_91_tkeep),
        .m_axis_oarg_91_tstrb(m_axis_oarg_91_tstrb),
        .m_axis_oarg_91_tdata(m_axis_oarg_91_tdata),
        .m_axis_oarg_91_tready(m_axis_oarg_91_tready),
        .ap_axis_oarg_91_tlast(ap_axis_oarg_91_tlast),
        .ap_axis_oarg_91_tvalid(ap_axis_oarg_91_tvalid),
        .ap_axis_oarg_91_tkeep(ap_axis_oarg_91_tkeep),
        .ap_axis_oarg_91_tstrb(ap_axis_oarg_91_tstrb),
        .ap_axis_oarg_91_tdata(ap_axis_oarg_91_tdata),
        .ap_axis_oarg_91_tready(ap_axis_oarg_91_tready),
        .m_axis_oarg_92_aclk(m_axis_oarg_92_aclk),
        .m_axis_oarg_92_aresetn(m_axis_oarg_92_aresetn),
        .m_axis_oarg_92_tlast(m_axis_oarg_92_tlast),
        .m_axis_oarg_92_tvalid(m_axis_oarg_92_tvalid),
        .m_axis_oarg_92_tkeep(m_axis_oarg_92_tkeep),
        .m_axis_oarg_92_tstrb(m_axis_oarg_92_tstrb),
        .m_axis_oarg_92_tdata(m_axis_oarg_92_tdata),
        .m_axis_oarg_92_tready(m_axis_oarg_92_tready),
        .ap_axis_oarg_92_tlast(ap_axis_oarg_92_tlast),
        .ap_axis_oarg_92_tvalid(ap_axis_oarg_92_tvalid),
        .ap_axis_oarg_92_tkeep(ap_axis_oarg_92_tkeep),
        .ap_axis_oarg_92_tstrb(ap_axis_oarg_92_tstrb),
        .ap_axis_oarg_92_tdata(ap_axis_oarg_92_tdata),
        .ap_axis_oarg_92_tready(ap_axis_oarg_92_tready),
        .m_axis_oarg_93_aclk(m_axis_oarg_93_aclk),
        .m_axis_oarg_93_aresetn(m_axis_oarg_93_aresetn),
        .m_axis_oarg_93_tlast(m_axis_oarg_93_tlast),
        .m_axis_oarg_93_tvalid(m_axis_oarg_93_tvalid),
        .m_axis_oarg_93_tkeep(m_axis_oarg_93_tkeep),
        .m_axis_oarg_93_tstrb(m_axis_oarg_93_tstrb),
        .m_axis_oarg_93_tdata(m_axis_oarg_93_tdata),
        .m_axis_oarg_93_tready(m_axis_oarg_93_tready),
        .ap_axis_oarg_93_tlast(ap_axis_oarg_93_tlast),
        .ap_axis_oarg_93_tvalid(ap_axis_oarg_93_tvalid),
        .ap_axis_oarg_93_tkeep(ap_axis_oarg_93_tkeep),
        .ap_axis_oarg_93_tstrb(ap_axis_oarg_93_tstrb),
        .ap_axis_oarg_93_tdata(ap_axis_oarg_93_tdata),
        .ap_axis_oarg_93_tready(ap_axis_oarg_93_tready),
        .m_axis_oarg_94_aclk(m_axis_oarg_94_aclk),
        .m_axis_oarg_94_aresetn(m_axis_oarg_94_aresetn),
        .m_axis_oarg_94_tlast(m_axis_oarg_94_tlast),
        .m_axis_oarg_94_tvalid(m_axis_oarg_94_tvalid),
        .m_axis_oarg_94_tkeep(m_axis_oarg_94_tkeep),
        .m_axis_oarg_94_tstrb(m_axis_oarg_94_tstrb),
        .m_axis_oarg_94_tdata(m_axis_oarg_94_tdata),
        .m_axis_oarg_94_tready(m_axis_oarg_94_tready),
        .ap_axis_oarg_94_tlast(ap_axis_oarg_94_tlast),
        .ap_axis_oarg_94_tvalid(ap_axis_oarg_94_tvalid),
        .ap_axis_oarg_94_tkeep(ap_axis_oarg_94_tkeep),
        .ap_axis_oarg_94_tstrb(ap_axis_oarg_94_tstrb),
        .ap_axis_oarg_94_tdata(ap_axis_oarg_94_tdata),
        .ap_axis_oarg_94_tready(ap_axis_oarg_94_tready),
        .m_axis_oarg_95_aclk(m_axis_oarg_95_aclk),
        .m_axis_oarg_95_aresetn(m_axis_oarg_95_aresetn),
        .m_axis_oarg_95_tlast(m_axis_oarg_95_tlast),
        .m_axis_oarg_95_tvalid(m_axis_oarg_95_tvalid),
        .m_axis_oarg_95_tkeep(m_axis_oarg_95_tkeep),
        .m_axis_oarg_95_tstrb(m_axis_oarg_95_tstrb),
        .m_axis_oarg_95_tdata(m_axis_oarg_95_tdata),
        .m_axis_oarg_95_tready(m_axis_oarg_95_tready),
        .ap_axis_oarg_95_tlast(ap_axis_oarg_95_tlast),
        .ap_axis_oarg_95_tvalid(ap_axis_oarg_95_tvalid),
        .ap_axis_oarg_95_tkeep(ap_axis_oarg_95_tkeep),
        .ap_axis_oarg_95_tstrb(ap_axis_oarg_95_tstrb),
        .ap_axis_oarg_95_tdata(ap_axis_oarg_95_tdata),
        .ap_axis_oarg_95_tready(ap_axis_oarg_95_tready),
        .m_axis_oarg_96_aclk(m_axis_oarg_96_aclk),
        .m_axis_oarg_96_aresetn(m_axis_oarg_96_aresetn),
        .m_axis_oarg_96_tlast(m_axis_oarg_96_tlast),
        .m_axis_oarg_96_tvalid(m_axis_oarg_96_tvalid),
        .m_axis_oarg_96_tkeep(m_axis_oarg_96_tkeep),
        .m_axis_oarg_96_tstrb(m_axis_oarg_96_tstrb),
        .m_axis_oarg_96_tdata(m_axis_oarg_96_tdata),
        .m_axis_oarg_96_tready(m_axis_oarg_96_tready),
        .ap_axis_oarg_96_tlast(ap_axis_oarg_96_tlast),
        .ap_axis_oarg_96_tvalid(ap_axis_oarg_96_tvalid),
        .ap_axis_oarg_96_tkeep(ap_axis_oarg_96_tkeep),
        .ap_axis_oarg_96_tstrb(ap_axis_oarg_96_tstrb),
        .ap_axis_oarg_96_tdata(ap_axis_oarg_96_tdata),
        .ap_axis_oarg_96_tready(ap_axis_oarg_96_tready),
        .m_axis_oarg_97_aclk(m_axis_oarg_97_aclk),
        .m_axis_oarg_97_aresetn(m_axis_oarg_97_aresetn),
        .m_axis_oarg_97_tlast(m_axis_oarg_97_tlast),
        .m_axis_oarg_97_tvalid(m_axis_oarg_97_tvalid),
        .m_axis_oarg_97_tkeep(m_axis_oarg_97_tkeep),
        .m_axis_oarg_97_tstrb(m_axis_oarg_97_tstrb),
        .m_axis_oarg_97_tdata(m_axis_oarg_97_tdata),
        .m_axis_oarg_97_tready(m_axis_oarg_97_tready),
        .ap_axis_oarg_97_tlast(ap_axis_oarg_97_tlast),
        .ap_axis_oarg_97_tvalid(ap_axis_oarg_97_tvalid),
        .ap_axis_oarg_97_tkeep(ap_axis_oarg_97_tkeep),
        .ap_axis_oarg_97_tstrb(ap_axis_oarg_97_tstrb),
        .ap_axis_oarg_97_tdata(ap_axis_oarg_97_tdata),
        .ap_axis_oarg_97_tready(ap_axis_oarg_97_tready),
        .m_axis_oarg_98_aclk(m_axis_oarg_98_aclk),
        .m_axis_oarg_98_aresetn(m_axis_oarg_98_aresetn),
        .m_axis_oarg_98_tlast(m_axis_oarg_98_tlast),
        .m_axis_oarg_98_tvalid(m_axis_oarg_98_tvalid),
        .m_axis_oarg_98_tkeep(m_axis_oarg_98_tkeep),
        .m_axis_oarg_98_tstrb(m_axis_oarg_98_tstrb),
        .m_axis_oarg_98_tdata(m_axis_oarg_98_tdata),
        .m_axis_oarg_98_tready(m_axis_oarg_98_tready),
        .ap_axis_oarg_98_tlast(ap_axis_oarg_98_tlast),
        .ap_axis_oarg_98_tvalid(ap_axis_oarg_98_tvalid),
        .ap_axis_oarg_98_tkeep(ap_axis_oarg_98_tkeep),
        .ap_axis_oarg_98_tstrb(ap_axis_oarg_98_tstrb),
        .ap_axis_oarg_98_tdata(ap_axis_oarg_98_tdata),
        .ap_axis_oarg_98_tready(ap_axis_oarg_98_tready),
        .m_axis_oarg_99_aclk(m_axis_oarg_99_aclk),
        .m_axis_oarg_99_aresetn(m_axis_oarg_99_aresetn),
        .m_axis_oarg_99_tlast(m_axis_oarg_99_tlast),
        .m_axis_oarg_99_tvalid(m_axis_oarg_99_tvalid),
        .m_axis_oarg_99_tkeep(m_axis_oarg_99_tkeep),
        .m_axis_oarg_99_tstrb(m_axis_oarg_99_tstrb),
        .m_axis_oarg_99_tdata(m_axis_oarg_99_tdata),
        .m_axis_oarg_99_tready(m_axis_oarg_99_tready),
        .ap_axis_oarg_99_tlast(ap_axis_oarg_99_tlast),
        .ap_axis_oarg_99_tvalid(ap_axis_oarg_99_tvalid),
        .ap_axis_oarg_99_tkeep(ap_axis_oarg_99_tkeep),
        .ap_axis_oarg_99_tstrb(ap_axis_oarg_99_tstrb),
        .ap_axis_oarg_99_tdata(ap_axis_oarg_99_tdata),
        .ap_axis_oarg_99_tready(ap_axis_oarg_99_tready),
        .m_axis_oarg_100_aclk(m_axis_oarg_100_aclk),
        .m_axis_oarg_100_aresetn(m_axis_oarg_100_aresetn),
        .m_axis_oarg_100_tlast(m_axis_oarg_100_tlast),
        .m_axis_oarg_100_tvalid(m_axis_oarg_100_tvalid),
        .m_axis_oarg_100_tkeep(m_axis_oarg_100_tkeep),
        .m_axis_oarg_100_tstrb(m_axis_oarg_100_tstrb),
        .m_axis_oarg_100_tdata(m_axis_oarg_100_tdata),
        .m_axis_oarg_100_tready(m_axis_oarg_100_tready),
        .ap_axis_oarg_100_tlast(ap_axis_oarg_100_tlast),
        .ap_axis_oarg_100_tvalid(ap_axis_oarg_100_tvalid),
        .ap_axis_oarg_100_tkeep(ap_axis_oarg_100_tkeep),
        .ap_axis_oarg_100_tstrb(ap_axis_oarg_100_tstrb),
        .ap_axis_oarg_100_tdata(ap_axis_oarg_100_tdata),
        .ap_axis_oarg_100_tready(ap_axis_oarg_100_tready),
        .m_axis_oarg_101_aclk(m_axis_oarg_101_aclk),
        .m_axis_oarg_101_aresetn(m_axis_oarg_101_aresetn),
        .m_axis_oarg_101_tlast(m_axis_oarg_101_tlast),
        .m_axis_oarg_101_tvalid(m_axis_oarg_101_tvalid),
        .m_axis_oarg_101_tkeep(m_axis_oarg_101_tkeep),
        .m_axis_oarg_101_tstrb(m_axis_oarg_101_tstrb),
        .m_axis_oarg_101_tdata(m_axis_oarg_101_tdata),
        .m_axis_oarg_101_tready(m_axis_oarg_101_tready),
        .ap_axis_oarg_101_tlast(ap_axis_oarg_101_tlast),
        .ap_axis_oarg_101_tvalid(ap_axis_oarg_101_tvalid),
        .ap_axis_oarg_101_tkeep(ap_axis_oarg_101_tkeep),
        .ap_axis_oarg_101_tstrb(ap_axis_oarg_101_tstrb),
        .ap_axis_oarg_101_tdata(ap_axis_oarg_101_tdata),
        .ap_axis_oarg_101_tready(ap_axis_oarg_101_tready),
        .m_axis_oarg_102_aclk(m_axis_oarg_102_aclk),
        .m_axis_oarg_102_aresetn(m_axis_oarg_102_aresetn),
        .m_axis_oarg_102_tlast(m_axis_oarg_102_tlast),
        .m_axis_oarg_102_tvalid(m_axis_oarg_102_tvalid),
        .m_axis_oarg_102_tkeep(m_axis_oarg_102_tkeep),
        .m_axis_oarg_102_tstrb(m_axis_oarg_102_tstrb),
        .m_axis_oarg_102_tdata(m_axis_oarg_102_tdata),
        .m_axis_oarg_102_tready(m_axis_oarg_102_tready),
        .ap_axis_oarg_102_tlast(ap_axis_oarg_102_tlast),
        .ap_axis_oarg_102_tvalid(ap_axis_oarg_102_tvalid),
        .ap_axis_oarg_102_tkeep(ap_axis_oarg_102_tkeep),
        .ap_axis_oarg_102_tstrb(ap_axis_oarg_102_tstrb),
        .ap_axis_oarg_102_tdata(ap_axis_oarg_102_tdata),
        .ap_axis_oarg_102_tready(ap_axis_oarg_102_tready),
        .m_axis_oarg_103_aclk(m_axis_oarg_103_aclk),
        .m_axis_oarg_103_aresetn(m_axis_oarg_103_aresetn),
        .m_axis_oarg_103_tlast(m_axis_oarg_103_tlast),
        .m_axis_oarg_103_tvalid(m_axis_oarg_103_tvalid),
        .m_axis_oarg_103_tkeep(m_axis_oarg_103_tkeep),
        .m_axis_oarg_103_tstrb(m_axis_oarg_103_tstrb),
        .m_axis_oarg_103_tdata(m_axis_oarg_103_tdata),
        .m_axis_oarg_103_tready(m_axis_oarg_103_tready),
        .ap_axis_oarg_103_tlast(ap_axis_oarg_103_tlast),
        .ap_axis_oarg_103_tvalid(ap_axis_oarg_103_tvalid),
        .ap_axis_oarg_103_tkeep(ap_axis_oarg_103_tkeep),
        .ap_axis_oarg_103_tstrb(ap_axis_oarg_103_tstrb),
        .ap_axis_oarg_103_tdata(ap_axis_oarg_103_tdata),
        .ap_axis_oarg_103_tready(ap_axis_oarg_103_tready),
        .m_axis_oarg_104_aclk(m_axis_oarg_104_aclk),
        .m_axis_oarg_104_aresetn(m_axis_oarg_104_aresetn),
        .m_axis_oarg_104_tlast(m_axis_oarg_104_tlast),
        .m_axis_oarg_104_tvalid(m_axis_oarg_104_tvalid),
        .m_axis_oarg_104_tkeep(m_axis_oarg_104_tkeep),
        .m_axis_oarg_104_tstrb(m_axis_oarg_104_tstrb),
        .m_axis_oarg_104_tdata(m_axis_oarg_104_tdata),
        .m_axis_oarg_104_tready(m_axis_oarg_104_tready),
        .ap_axis_oarg_104_tlast(ap_axis_oarg_104_tlast),
        .ap_axis_oarg_104_tvalid(ap_axis_oarg_104_tvalid),
        .ap_axis_oarg_104_tkeep(ap_axis_oarg_104_tkeep),
        .ap_axis_oarg_104_tstrb(ap_axis_oarg_104_tstrb),
        .ap_axis_oarg_104_tdata(ap_axis_oarg_104_tdata),
        .ap_axis_oarg_104_tready(ap_axis_oarg_104_tready),
        .m_axis_oarg_105_aclk(m_axis_oarg_105_aclk),
        .m_axis_oarg_105_aresetn(m_axis_oarg_105_aresetn),
        .m_axis_oarg_105_tlast(m_axis_oarg_105_tlast),
        .m_axis_oarg_105_tvalid(m_axis_oarg_105_tvalid),
        .m_axis_oarg_105_tkeep(m_axis_oarg_105_tkeep),
        .m_axis_oarg_105_tstrb(m_axis_oarg_105_tstrb),
        .m_axis_oarg_105_tdata(m_axis_oarg_105_tdata),
        .m_axis_oarg_105_tready(m_axis_oarg_105_tready),
        .ap_axis_oarg_105_tlast(ap_axis_oarg_105_tlast),
        .ap_axis_oarg_105_tvalid(ap_axis_oarg_105_tvalid),
        .ap_axis_oarg_105_tkeep(ap_axis_oarg_105_tkeep),
        .ap_axis_oarg_105_tstrb(ap_axis_oarg_105_tstrb),
        .ap_axis_oarg_105_tdata(ap_axis_oarg_105_tdata),
        .ap_axis_oarg_105_tready(ap_axis_oarg_105_tready),
        .m_axis_oarg_106_aclk(m_axis_oarg_106_aclk),
        .m_axis_oarg_106_aresetn(m_axis_oarg_106_aresetn),
        .m_axis_oarg_106_tlast(m_axis_oarg_106_tlast),
        .m_axis_oarg_106_tvalid(m_axis_oarg_106_tvalid),
        .m_axis_oarg_106_tkeep(m_axis_oarg_106_tkeep),
        .m_axis_oarg_106_tstrb(m_axis_oarg_106_tstrb),
        .m_axis_oarg_106_tdata(m_axis_oarg_106_tdata),
        .m_axis_oarg_106_tready(m_axis_oarg_106_tready),
        .ap_axis_oarg_106_tlast(ap_axis_oarg_106_tlast),
        .ap_axis_oarg_106_tvalid(ap_axis_oarg_106_tvalid),
        .ap_axis_oarg_106_tkeep(ap_axis_oarg_106_tkeep),
        .ap_axis_oarg_106_tstrb(ap_axis_oarg_106_tstrb),
        .ap_axis_oarg_106_tdata(ap_axis_oarg_106_tdata),
        .ap_axis_oarg_106_tready(ap_axis_oarg_106_tready),
        .m_axis_oarg_107_aclk(m_axis_oarg_107_aclk),
        .m_axis_oarg_107_aresetn(m_axis_oarg_107_aresetn),
        .m_axis_oarg_107_tlast(m_axis_oarg_107_tlast),
        .m_axis_oarg_107_tvalid(m_axis_oarg_107_tvalid),
        .m_axis_oarg_107_tkeep(m_axis_oarg_107_tkeep),
        .m_axis_oarg_107_tstrb(m_axis_oarg_107_tstrb),
        .m_axis_oarg_107_tdata(m_axis_oarg_107_tdata),
        .m_axis_oarg_107_tready(m_axis_oarg_107_tready),
        .ap_axis_oarg_107_tlast(ap_axis_oarg_107_tlast),
        .ap_axis_oarg_107_tvalid(ap_axis_oarg_107_tvalid),
        .ap_axis_oarg_107_tkeep(ap_axis_oarg_107_tkeep),
        .ap_axis_oarg_107_tstrb(ap_axis_oarg_107_tstrb),
        .ap_axis_oarg_107_tdata(ap_axis_oarg_107_tdata),
        .ap_axis_oarg_107_tready(ap_axis_oarg_107_tready),
        .m_axis_oarg_108_aclk(m_axis_oarg_108_aclk),
        .m_axis_oarg_108_aresetn(m_axis_oarg_108_aresetn),
        .m_axis_oarg_108_tlast(m_axis_oarg_108_tlast),
        .m_axis_oarg_108_tvalid(m_axis_oarg_108_tvalid),
        .m_axis_oarg_108_tkeep(m_axis_oarg_108_tkeep),
        .m_axis_oarg_108_tstrb(m_axis_oarg_108_tstrb),
        .m_axis_oarg_108_tdata(m_axis_oarg_108_tdata),
        .m_axis_oarg_108_tready(m_axis_oarg_108_tready),
        .ap_axis_oarg_108_tlast(ap_axis_oarg_108_tlast),
        .ap_axis_oarg_108_tvalid(ap_axis_oarg_108_tvalid),
        .ap_axis_oarg_108_tkeep(ap_axis_oarg_108_tkeep),
        .ap_axis_oarg_108_tstrb(ap_axis_oarg_108_tstrb),
        .ap_axis_oarg_108_tdata(ap_axis_oarg_108_tdata),
        .ap_axis_oarg_108_tready(ap_axis_oarg_108_tready),
        .m_axis_oarg_109_aclk(m_axis_oarg_109_aclk),
        .m_axis_oarg_109_aresetn(m_axis_oarg_109_aresetn),
        .m_axis_oarg_109_tlast(m_axis_oarg_109_tlast),
        .m_axis_oarg_109_tvalid(m_axis_oarg_109_tvalid),
        .m_axis_oarg_109_tkeep(m_axis_oarg_109_tkeep),
        .m_axis_oarg_109_tstrb(m_axis_oarg_109_tstrb),
        .m_axis_oarg_109_tdata(m_axis_oarg_109_tdata),
        .m_axis_oarg_109_tready(m_axis_oarg_109_tready),
        .ap_axis_oarg_109_tlast(ap_axis_oarg_109_tlast),
        .ap_axis_oarg_109_tvalid(ap_axis_oarg_109_tvalid),
        .ap_axis_oarg_109_tkeep(ap_axis_oarg_109_tkeep),
        .ap_axis_oarg_109_tstrb(ap_axis_oarg_109_tstrb),
        .ap_axis_oarg_109_tdata(ap_axis_oarg_109_tdata),
        .ap_axis_oarg_109_tready(ap_axis_oarg_109_tready),
        .m_axis_oarg_110_aclk(m_axis_oarg_110_aclk),
        .m_axis_oarg_110_aresetn(m_axis_oarg_110_aresetn),
        .m_axis_oarg_110_tlast(m_axis_oarg_110_tlast),
        .m_axis_oarg_110_tvalid(m_axis_oarg_110_tvalid),
        .m_axis_oarg_110_tkeep(m_axis_oarg_110_tkeep),
        .m_axis_oarg_110_tstrb(m_axis_oarg_110_tstrb),
        .m_axis_oarg_110_tdata(m_axis_oarg_110_tdata),
        .m_axis_oarg_110_tready(m_axis_oarg_110_tready),
        .ap_axis_oarg_110_tlast(ap_axis_oarg_110_tlast),
        .ap_axis_oarg_110_tvalid(ap_axis_oarg_110_tvalid),
        .ap_axis_oarg_110_tkeep(ap_axis_oarg_110_tkeep),
        .ap_axis_oarg_110_tstrb(ap_axis_oarg_110_tstrb),
        .ap_axis_oarg_110_tdata(ap_axis_oarg_110_tdata),
        .ap_axis_oarg_110_tready(ap_axis_oarg_110_tready),
        .m_axis_oarg_111_aclk(m_axis_oarg_111_aclk),
        .m_axis_oarg_111_aresetn(m_axis_oarg_111_aresetn),
        .m_axis_oarg_111_tlast(m_axis_oarg_111_tlast),
        .m_axis_oarg_111_tvalid(m_axis_oarg_111_tvalid),
        .m_axis_oarg_111_tkeep(m_axis_oarg_111_tkeep),
        .m_axis_oarg_111_tstrb(m_axis_oarg_111_tstrb),
        .m_axis_oarg_111_tdata(m_axis_oarg_111_tdata),
        .m_axis_oarg_111_tready(m_axis_oarg_111_tready),
        .ap_axis_oarg_111_tlast(ap_axis_oarg_111_tlast),
        .ap_axis_oarg_111_tvalid(ap_axis_oarg_111_tvalid),
        .ap_axis_oarg_111_tkeep(ap_axis_oarg_111_tkeep),
        .ap_axis_oarg_111_tstrb(ap_axis_oarg_111_tstrb),
        .ap_axis_oarg_111_tdata(ap_axis_oarg_111_tdata),
        .ap_axis_oarg_111_tready(ap_axis_oarg_111_tready),
        .m_axis_oarg_112_aclk(m_axis_oarg_112_aclk),
        .m_axis_oarg_112_aresetn(m_axis_oarg_112_aresetn),
        .m_axis_oarg_112_tlast(m_axis_oarg_112_tlast),
        .m_axis_oarg_112_tvalid(m_axis_oarg_112_tvalid),
        .m_axis_oarg_112_tkeep(m_axis_oarg_112_tkeep),
        .m_axis_oarg_112_tstrb(m_axis_oarg_112_tstrb),
        .m_axis_oarg_112_tdata(m_axis_oarg_112_tdata),
        .m_axis_oarg_112_tready(m_axis_oarg_112_tready),
        .ap_axis_oarg_112_tlast(ap_axis_oarg_112_tlast),
        .ap_axis_oarg_112_tvalid(ap_axis_oarg_112_tvalid),
        .ap_axis_oarg_112_tkeep(ap_axis_oarg_112_tkeep),
        .ap_axis_oarg_112_tstrb(ap_axis_oarg_112_tstrb),
        .ap_axis_oarg_112_tdata(ap_axis_oarg_112_tdata),
        .ap_axis_oarg_112_tready(ap_axis_oarg_112_tready),
        .m_axis_oarg_113_aclk(m_axis_oarg_113_aclk),
        .m_axis_oarg_113_aresetn(m_axis_oarg_113_aresetn),
        .m_axis_oarg_113_tlast(m_axis_oarg_113_tlast),
        .m_axis_oarg_113_tvalid(m_axis_oarg_113_tvalid),
        .m_axis_oarg_113_tkeep(m_axis_oarg_113_tkeep),
        .m_axis_oarg_113_tstrb(m_axis_oarg_113_tstrb),
        .m_axis_oarg_113_tdata(m_axis_oarg_113_tdata),
        .m_axis_oarg_113_tready(m_axis_oarg_113_tready),
        .ap_axis_oarg_113_tlast(ap_axis_oarg_113_tlast),
        .ap_axis_oarg_113_tvalid(ap_axis_oarg_113_tvalid),
        .ap_axis_oarg_113_tkeep(ap_axis_oarg_113_tkeep),
        .ap_axis_oarg_113_tstrb(ap_axis_oarg_113_tstrb),
        .ap_axis_oarg_113_tdata(ap_axis_oarg_113_tdata),
        .ap_axis_oarg_113_tready(ap_axis_oarg_113_tready),
        .m_axis_oarg_114_aclk(m_axis_oarg_114_aclk),
        .m_axis_oarg_114_aresetn(m_axis_oarg_114_aresetn),
        .m_axis_oarg_114_tlast(m_axis_oarg_114_tlast),
        .m_axis_oarg_114_tvalid(m_axis_oarg_114_tvalid),
        .m_axis_oarg_114_tkeep(m_axis_oarg_114_tkeep),
        .m_axis_oarg_114_tstrb(m_axis_oarg_114_tstrb),
        .m_axis_oarg_114_tdata(m_axis_oarg_114_tdata),
        .m_axis_oarg_114_tready(m_axis_oarg_114_tready),
        .ap_axis_oarg_114_tlast(ap_axis_oarg_114_tlast),
        .ap_axis_oarg_114_tvalid(ap_axis_oarg_114_tvalid),
        .ap_axis_oarg_114_tkeep(ap_axis_oarg_114_tkeep),
        .ap_axis_oarg_114_tstrb(ap_axis_oarg_114_tstrb),
        .ap_axis_oarg_114_tdata(ap_axis_oarg_114_tdata),
        .ap_axis_oarg_114_tready(ap_axis_oarg_114_tready),
        .m_axis_oarg_115_aclk(m_axis_oarg_115_aclk),
        .m_axis_oarg_115_aresetn(m_axis_oarg_115_aresetn),
        .m_axis_oarg_115_tlast(m_axis_oarg_115_tlast),
        .m_axis_oarg_115_tvalid(m_axis_oarg_115_tvalid),
        .m_axis_oarg_115_tkeep(m_axis_oarg_115_tkeep),
        .m_axis_oarg_115_tstrb(m_axis_oarg_115_tstrb),
        .m_axis_oarg_115_tdata(m_axis_oarg_115_tdata),
        .m_axis_oarg_115_tready(m_axis_oarg_115_tready),
        .ap_axis_oarg_115_tlast(ap_axis_oarg_115_tlast),
        .ap_axis_oarg_115_tvalid(ap_axis_oarg_115_tvalid),
        .ap_axis_oarg_115_tkeep(ap_axis_oarg_115_tkeep),
        .ap_axis_oarg_115_tstrb(ap_axis_oarg_115_tstrb),
        .ap_axis_oarg_115_tdata(ap_axis_oarg_115_tdata),
        .ap_axis_oarg_115_tready(ap_axis_oarg_115_tready),
        .m_axis_oarg_116_aclk(m_axis_oarg_116_aclk),
        .m_axis_oarg_116_aresetn(m_axis_oarg_116_aresetn),
        .m_axis_oarg_116_tlast(m_axis_oarg_116_tlast),
        .m_axis_oarg_116_tvalid(m_axis_oarg_116_tvalid),
        .m_axis_oarg_116_tkeep(m_axis_oarg_116_tkeep),
        .m_axis_oarg_116_tstrb(m_axis_oarg_116_tstrb),
        .m_axis_oarg_116_tdata(m_axis_oarg_116_tdata),
        .m_axis_oarg_116_tready(m_axis_oarg_116_tready),
        .ap_axis_oarg_116_tlast(ap_axis_oarg_116_tlast),
        .ap_axis_oarg_116_tvalid(ap_axis_oarg_116_tvalid),
        .ap_axis_oarg_116_tkeep(ap_axis_oarg_116_tkeep),
        .ap_axis_oarg_116_tstrb(ap_axis_oarg_116_tstrb),
        .ap_axis_oarg_116_tdata(ap_axis_oarg_116_tdata),
        .ap_axis_oarg_116_tready(ap_axis_oarg_116_tready),
        .m_axis_oarg_117_aclk(m_axis_oarg_117_aclk),
        .m_axis_oarg_117_aresetn(m_axis_oarg_117_aresetn),
        .m_axis_oarg_117_tlast(m_axis_oarg_117_tlast),
        .m_axis_oarg_117_tvalid(m_axis_oarg_117_tvalid),
        .m_axis_oarg_117_tkeep(m_axis_oarg_117_tkeep),
        .m_axis_oarg_117_tstrb(m_axis_oarg_117_tstrb),
        .m_axis_oarg_117_tdata(m_axis_oarg_117_tdata),
        .m_axis_oarg_117_tready(m_axis_oarg_117_tready),
        .ap_axis_oarg_117_tlast(ap_axis_oarg_117_tlast),
        .ap_axis_oarg_117_tvalid(ap_axis_oarg_117_tvalid),
        .ap_axis_oarg_117_tkeep(ap_axis_oarg_117_tkeep),
        .ap_axis_oarg_117_tstrb(ap_axis_oarg_117_tstrb),
        .ap_axis_oarg_117_tdata(ap_axis_oarg_117_tdata),
        .ap_axis_oarg_117_tready(ap_axis_oarg_117_tready),
        .m_axis_oarg_118_aclk(m_axis_oarg_118_aclk),
        .m_axis_oarg_118_aresetn(m_axis_oarg_118_aresetn),
        .m_axis_oarg_118_tlast(m_axis_oarg_118_tlast),
        .m_axis_oarg_118_tvalid(m_axis_oarg_118_tvalid),
        .m_axis_oarg_118_tkeep(m_axis_oarg_118_tkeep),
        .m_axis_oarg_118_tstrb(m_axis_oarg_118_tstrb),
        .m_axis_oarg_118_tdata(m_axis_oarg_118_tdata),
        .m_axis_oarg_118_tready(m_axis_oarg_118_tready),
        .ap_axis_oarg_118_tlast(ap_axis_oarg_118_tlast),
        .ap_axis_oarg_118_tvalid(ap_axis_oarg_118_tvalid),
        .ap_axis_oarg_118_tkeep(ap_axis_oarg_118_tkeep),
        .ap_axis_oarg_118_tstrb(ap_axis_oarg_118_tstrb),
        .ap_axis_oarg_118_tdata(ap_axis_oarg_118_tdata),
        .ap_axis_oarg_118_tready(ap_axis_oarg_118_tready),
        .m_axis_oarg_119_aclk(m_axis_oarg_119_aclk),
        .m_axis_oarg_119_aresetn(m_axis_oarg_119_aresetn),
        .m_axis_oarg_119_tlast(m_axis_oarg_119_tlast),
        .m_axis_oarg_119_tvalid(m_axis_oarg_119_tvalid),
        .m_axis_oarg_119_tkeep(m_axis_oarg_119_tkeep),
        .m_axis_oarg_119_tstrb(m_axis_oarg_119_tstrb),
        .m_axis_oarg_119_tdata(m_axis_oarg_119_tdata),
        .m_axis_oarg_119_tready(m_axis_oarg_119_tready),
        .ap_axis_oarg_119_tlast(ap_axis_oarg_119_tlast),
        .ap_axis_oarg_119_tvalid(ap_axis_oarg_119_tvalid),
        .ap_axis_oarg_119_tkeep(ap_axis_oarg_119_tkeep),
        .ap_axis_oarg_119_tstrb(ap_axis_oarg_119_tstrb),
        .ap_axis_oarg_119_tdata(ap_axis_oarg_119_tdata),
        .ap_axis_oarg_119_tready(ap_axis_oarg_119_tready),
        .m_axis_oarg_120_aclk(m_axis_oarg_120_aclk),
        .m_axis_oarg_120_aresetn(m_axis_oarg_120_aresetn),
        .m_axis_oarg_120_tlast(m_axis_oarg_120_tlast),
        .m_axis_oarg_120_tvalid(m_axis_oarg_120_tvalid),
        .m_axis_oarg_120_tkeep(m_axis_oarg_120_tkeep),
        .m_axis_oarg_120_tstrb(m_axis_oarg_120_tstrb),
        .m_axis_oarg_120_tdata(m_axis_oarg_120_tdata),
        .m_axis_oarg_120_tready(m_axis_oarg_120_tready),
        .ap_axis_oarg_120_tlast(ap_axis_oarg_120_tlast),
        .ap_axis_oarg_120_tvalid(ap_axis_oarg_120_tvalid),
        .ap_axis_oarg_120_tkeep(ap_axis_oarg_120_tkeep),
        .ap_axis_oarg_120_tstrb(ap_axis_oarg_120_tstrb),
        .ap_axis_oarg_120_tdata(ap_axis_oarg_120_tdata),
        .ap_axis_oarg_120_tready(ap_axis_oarg_120_tready),
        .m_axis_oarg_121_aclk(m_axis_oarg_121_aclk),
        .m_axis_oarg_121_aresetn(m_axis_oarg_121_aresetn),
        .m_axis_oarg_121_tlast(m_axis_oarg_121_tlast),
        .m_axis_oarg_121_tvalid(m_axis_oarg_121_tvalid),
        .m_axis_oarg_121_tkeep(m_axis_oarg_121_tkeep),
        .m_axis_oarg_121_tstrb(m_axis_oarg_121_tstrb),
        .m_axis_oarg_121_tdata(m_axis_oarg_121_tdata),
        .m_axis_oarg_121_tready(m_axis_oarg_121_tready),
        .ap_axis_oarg_121_tlast(ap_axis_oarg_121_tlast),
        .ap_axis_oarg_121_tvalid(ap_axis_oarg_121_tvalid),
        .ap_axis_oarg_121_tkeep(ap_axis_oarg_121_tkeep),
        .ap_axis_oarg_121_tstrb(ap_axis_oarg_121_tstrb),
        .ap_axis_oarg_121_tdata(ap_axis_oarg_121_tdata),
        .ap_axis_oarg_121_tready(ap_axis_oarg_121_tready),
        .m_axis_oarg_122_aclk(m_axis_oarg_122_aclk),
        .m_axis_oarg_122_aresetn(m_axis_oarg_122_aresetn),
        .m_axis_oarg_122_tlast(m_axis_oarg_122_tlast),
        .m_axis_oarg_122_tvalid(m_axis_oarg_122_tvalid),
        .m_axis_oarg_122_tkeep(m_axis_oarg_122_tkeep),
        .m_axis_oarg_122_tstrb(m_axis_oarg_122_tstrb),
        .m_axis_oarg_122_tdata(m_axis_oarg_122_tdata),
        .m_axis_oarg_122_tready(m_axis_oarg_122_tready),
        .ap_axis_oarg_122_tlast(ap_axis_oarg_122_tlast),
        .ap_axis_oarg_122_tvalid(ap_axis_oarg_122_tvalid),
        .ap_axis_oarg_122_tkeep(ap_axis_oarg_122_tkeep),
        .ap_axis_oarg_122_tstrb(ap_axis_oarg_122_tstrb),
        .ap_axis_oarg_122_tdata(ap_axis_oarg_122_tdata),
        .ap_axis_oarg_122_tready(ap_axis_oarg_122_tready),
        .m_axis_oarg_123_aclk(m_axis_oarg_123_aclk),
        .m_axis_oarg_123_aresetn(m_axis_oarg_123_aresetn),
        .m_axis_oarg_123_tlast(m_axis_oarg_123_tlast),
        .m_axis_oarg_123_tvalid(m_axis_oarg_123_tvalid),
        .m_axis_oarg_123_tkeep(m_axis_oarg_123_tkeep),
        .m_axis_oarg_123_tstrb(m_axis_oarg_123_tstrb),
        .m_axis_oarg_123_tdata(m_axis_oarg_123_tdata),
        .m_axis_oarg_123_tready(m_axis_oarg_123_tready),
        .ap_axis_oarg_123_tlast(ap_axis_oarg_123_tlast),
        .ap_axis_oarg_123_tvalid(ap_axis_oarg_123_tvalid),
        .ap_axis_oarg_123_tkeep(ap_axis_oarg_123_tkeep),
        .ap_axis_oarg_123_tstrb(ap_axis_oarg_123_tstrb),
        .ap_axis_oarg_123_tdata(ap_axis_oarg_123_tdata),
        .ap_axis_oarg_123_tready(ap_axis_oarg_123_tready),
        .m_axis_oarg_124_aclk(m_axis_oarg_124_aclk),
        .m_axis_oarg_124_aresetn(m_axis_oarg_124_aresetn),
        .m_axis_oarg_124_tlast(m_axis_oarg_124_tlast),
        .m_axis_oarg_124_tvalid(m_axis_oarg_124_tvalid),
        .m_axis_oarg_124_tkeep(m_axis_oarg_124_tkeep),
        .m_axis_oarg_124_tstrb(m_axis_oarg_124_tstrb),
        .m_axis_oarg_124_tdata(m_axis_oarg_124_tdata),
        .m_axis_oarg_124_tready(m_axis_oarg_124_tready),
        .ap_axis_oarg_124_tlast(ap_axis_oarg_124_tlast),
        .ap_axis_oarg_124_tvalid(ap_axis_oarg_124_tvalid),
        .ap_axis_oarg_124_tkeep(ap_axis_oarg_124_tkeep),
        .ap_axis_oarg_124_tstrb(ap_axis_oarg_124_tstrb),
        .ap_axis_oarg_124_tdata(ap_axis_oarg_124_tdata),
        .ap_axis_oarg_124_tready(ap_axis_oarg_124_tready),
        .m_axis_oarg_125_aclk(m_axis_oarg_125_aclk),
        .m_axis_oarg_125_aresetn(m_axis_oarg_125_aresetn),
        .m_axis_oarg_125_tlast(m_axis_oarg_125_tlast),
        .m_axis_oarg_125_tvalid(m_axis_oarg_125_tvalid),
        .m_axis_oarg_125_tkeep(m_axis_oarg_125_tkeep),
        .m_axis_oarg_125_tstrb(m_axis_oarg_125_tstrb),
        .m_axis_oarg_125_tdata(m_axis_oarg_125_tdata),
        .m_axis_oarg_125_tready(m_axis_oarg_125_tready),
        .ap_axis_oarg_125_tlast(ap_axis_oarg_125_tlast),
        .ap_axis_oarg_125_tvalid(ap_axis_oarg_125_tvalid),
        .ap_axis_oarg_125_tkeep(ap_axis_oarg_125_tkeep),
        .ap_axis_oarg_125_tstrb(ap_axis_oarg_125_tstrb),
        .ap_axis_oarg_125_tdata(ap_axis_oarg_125_tdata),
        .ap_axis_oarg_125_tready(ap_axis_oarg_125_tready),
        .m_axis_oarg_126_aclk(m_axis_oarg_126_aclk),
        .m_axis_oarg_126_aresetn(m_axis_oarg_126_aresetn),
        .m_axis_oarg_126_tlast(m_axis_oarg_126_tlast),
        .m_axis_oarg_126_tvalid(m_axis_oarg_126_tvalid),
        .m_axis_oarg_126_tkeep(m_axis_oarg_126_tkeep),
        .m_axis_oarg_126_tstrb(m_axis_oarg_126_tstrb),
        .m_axis_oarg_126_tdata(m_axis_oarg_126_tdata),
        .m_axis_oarg_126_tready(m_axis_oarg_126_tready),
        .ap_axis_oarg_126_tlast(ap_axis_oarg_126_tlast),
        .ap_axis_oarg_126_tvalid(ap_axis_oarg_126_tvalid),
        .ap_axis_oarg_126_tkeep(ap_axis_oarg_126_tkeep),
        .ap_axis_oarg_126_tstrb(ap_axis_oarg_126_tstrb),
        .ap_axis_oarg_126_tdata(ap_axis_oarg_126_tdata),
        .ap_axis_oarg_126_tready(ap_axis_oarg_126_tready),
        .m_axis_oarg_127_aclk(m_axis_oarg_127_aclk),
        .m_axis_oarg_127_aresetn(m_axis_oarg_127_aresetn),
        .m_axis_oarg_127_tlast(m_axis_oarg_127_tlast),
        .m_axis_oarg_127_tvalid(m_axis_oarg_127_tvalid),
        .m_axis_oarg_127_tkeep(m_axis_oarg_127_tkeep),
        .m_axis_oarg_127_tstrb(m_axis_oarg_127_tstrb),
        .m_axis_oarg_127_tdata(m_axis_oarg_127_tdata),
        .m_axis_oarg_127_tready(m_axis_oarg_127_tready),
        .ap_axis_oarg_127_tlast(ap_axis_oarg_127_tlast),
        .ap_axis_oarg_127_tvalid(ap_axis_oarg_127_tvalid),
        .ap_axis_oarg_127_tkeep(ap_axis_oarg_127_tkeep),
        .ap_axis_oarg_127_tstrb(ap_axis_oarg_127_tstrb),
        .ap_axis_oarg_127_tdata(ap_axis_oarg_127_tdata),
        .ap_axis_oarg_127_tready(ap_axis_oarg_127_tready)
    );
    
    aximm_args #(
        .C_NUM_AXIMMs(C_NUM_AXIMMs),
        .M_AXIMM_ADDR_WIDTH(M_AXIMM_ADDR_WIDTH),
        .M_AXIMM_0_ARUSER_WIDTH(M_AXIMM_0_ARUSER_WIDTH),
        .M_AXIMM_1_ARUSER_WIDTH(M_AXIMM_1_ARUSER_WIDTH),
        .M_AXIMM_2_ARUSER_WIDTH(M_AXIMM_2_ARUSER_WIDTH),
        .M_AXIMM_3_ARUSER_WIDTH(M_AXIMM_3_ARUSER_WIDTH),
        .M_AXIMM_4_ARUSER_WIDTH(M_AXIMM_4_ARUSER_WIDTH),
        .M_AXIMM_5_ARUSER_WIDTH(M_AXIMM_5_ARUSER_WIDTH),
        .M_AXIMM_6_ARUSER_WIDTH(M_AXIMM_6_ARUSER_WIDTH),
        .M_AXIMM_7_ARUSER_WIDTH(M_AXIMM_7_ARUSER_WIDTH),
        .M_AXIMM_8_ARUSER_WIDTH(M_AXIMM_8_ARUSER_WIDTH),
        .M_AXIMM_9_ARUSER_WIDTH(M_AXIMM_9_ARUSER_WIDTH),
        .M_AXIMM_10_ARUSER_WIDTH(M_AXIMM_10_ARUSER_WIDTH),
        .M_AXIMM_11_ARUSER_WIDTH(M_AXIMM_11_ARUSER_WIDTH),
        .M_AXIMM_12_ARUSER_WIDTH(M_AXIMM_12_ARUSER_WIDTH),
        .M_AXIMM_13_ARUSER_WIDTH(M_AXIMM_13_ARUSER_WIDTH),
        .M_AXIMM_14_ARUSER_WIDTH(M_AXIMM_14_ARUSER_WIDTH),
        .M_AXIMM_15_ARUSER_WIDTH(M_AXIMM_15_ARUSER_WIDTH),
        .M_AXIMM_16_ARUSER_WIDTH(M_AXIMM_16_ARUSER_WIDTH),
        .M_AXIMM_17_ARUSER_WIDTH(M_AXIMM_17_ARUSER_WIDTH),
        .M_AXIMM_18_ARUSER_WIDTH(M_AXIMM_18_ARUSER_WIDTH),
        .M_AXIMM_19_ARUSER_WIDTH(M_AXIMM_19_ARUSER_WIDTH),
        .M_AXIMM_20_ARUSER_WIDTH(M_AXIMM_20_ARUSER_WIDTH),
        .M_AXIMM_21_ARUSER_WIDTH(M_AXIMM_21_ARUSER_WIDTH),
        .M_AXIMM_22_ARUSER_WIDTH(M_AXIMM_22_ARUSER_WIDTH),
        .M_AXIMM_23_ARUSER_WIDTH(M_AXIMM_23_ARUSER_WIDTH),
        .M_AXIMM_24_ARUSER_WIDTH(M_AXIMM_24_ARUSER_WIDTH),
        .M_AXIMM_25_ARUSER_WIDTH(M_AXIMM_25_ARUSER_WIDTH),
        .M_AXIMM_26_ARUSER_WIDTH(M_AXIMM_26_ARUSER_WIDTH),
        .M_AXIMM_27_ARUSER_WIDTH(M_AXIMM_27_ARUSER_WIDTH),
        .M_AXIMM_28_ARUSER_WIDTH(M_AXIMM_28_ARUSER_WIDTH),
        .M_AXIMM_29_ARUSER_WIDTH(M_AXIMM_29_ARUSER_WIDTH),
        .M_AXIMM_30_ARUSER_WIDTH(M_AXIMM_30_ARUSER_WIDTH),
        .M_AXIMM_31_ARUSER_WIDTH(M_AXIMM_31_ARUSER_WIDTH),
        .M_AXIMM_32_ARUSER_WIDTH(M_AXIMM_32_ARUSER_WIDTH),
        .M_AXIMM_33_ARUSER_WIDTH(M_AXIMM_33_ARUSER_WIDTH),
        .M_AXIMM_34_ARUSER_WIDTH(M_AXIMM_34_ARUSER_WIDTH),
        .M_AXIMM_35_ARUSER_WIDTH(M_AXIMM_35_ARUSER_WIDTH),
        .M_AXIMM_36_ARUSER_WIDTH(M_AXIMM_36_ARUSER_WIDTH),
        .M_AXIMM_37_ARUSER_WIDTH(M_AXIMM_37_ARUSER_WIDTH),
        .M_AXIMM_38_ARUSER_WIDTH(M_AXIMM_38_ARUSER_WIDTH),
        .M_AXIMM_39_ARUSER_WIDTH(M_AXIMM_39_ARUSER_WIDTH),
        .M_AXIMM_40_ARUSER_WIDTH(M_AXIMM_40_ARUSER_WIDTH),
        .M_AXIMM_41_ARUSER_WIDTH(M_AXIMM_41_ARUSER_WIDTH),
        .M_AXIMM_42_ARUSER_WIDTH(M_AXIMM_42_ARUSER_WIDTH),
        .M_AXIMM_43_ARUSER_WIDTH(M_AXIMM_43_ARUSER_WIDTH),
        .M_AXIMM_44_ARUSER_WIDTH(M_AXIMM_44_ARUSER_WIDTH),
        .M_AXIMM_45_ARUSER_WIDTH(M_AXIMM_45_ARUSER_WIDTH),
        .M_AXIMM_46_ARUSER_WIDTH(M_AXIMM_46_ARUSER_WIDTH),
        .M_AXIMM_47_ARUSER_WIDTH(M_AXIMM_47_ARUSER_WIDTH),
        .M_AXIMM_48_ARUSER_WIDTH(M_AXIMM_48_ARUSER_WIDTH),
        .M_AXIMM_49_ARUSER_WIDTH(M_AXIMM_49_ARUSER_WIDTH),
        .M_AXIMM_50_ARUSER_WIDTH(M_AXIMM_50_ARUSER_WIDTH),
        .M_AXIMM_51_ARUSER_WIDTH(M_AXIMM_51_ARUSER_WIDTH),
        .M_AXIMM_52_ARUSER_WIDTH(M_AXIMM_52_ARUSER_WIDTH),
        .M_AXIMM_53_ARUSER_WIDTH(M_AXIMM_53_ARUSER_WIDTH),
        .M_AXIMM_54_ARUSER_WIDTH(M_AXIMM_54_ARUSER_WIDTH),
        .M_AXIMM_55_ARUSER_WIDTH(M_AXIMM_55_ARUSER_WIDTH),
        .M_AXIMM_56_ARUSER_WIDTH(M_AXIMM_56_ARUSER_WIDTH),
        .M_AXIMM_57_ARUSER_WIDTH(M_AXIMM_57_ARUSER_WIDTH),
        .M_AXIMM_58_ARUSER_WIDTH(M_AXIMM_58_ARUSER_WIDTH),
        .M_AXIMM_59_ARUSER_WIDTH(M_AXIMM_59_ARUSER_WIDTH),
        .M_AXIMM_60_ARUSER_WIDTH(M_AXIMM_60_ARUSER_WIDTH),
        .M_AXIMM_61_ARUSER_WIDTH(M_AXIMM_61_ARUSER_WIDTH),
        .M_AXIMM_62_ARUSER_WIDTH(M_AXIMM_62_ARUSER_WIDTH),
        .M_AXIMM_63_ARUSER_WIDTH(M_AXIMM_63_ARUSER_WIDTH),
        .M_AXIMM_64_ARUSER_WIDTH(M_AXIMM_64_ARUSER_WIDTH),
        .M_AXIMM_65_ARUSER_WIDTH(M_AXIMM_65_ARUSER_WIDTH),
        .M_AXIMM_66_ARUSER_WIDTH(M_AXIMM_66_ARUSER_WIDTH),
        .M_AXIMM_67_ARUSER_WIDTH(M_AXIMM_67_ARUSER_WIDTH),
        .M_AXIMM_68_ARUSER_WIDTH(M_AXIMM_68_ARUSER_WIDTH),
        .M_AXIMM_69_ARUSER_WIDTH(M_AXIMM_69_ARUSER_WIDTH),
        .M_AXIMM_70_ARUSER_WIDTH(M_AXIMM_70_ARUSER_WIDTH),
        .M_AXIMM_71_ARUSER_WIDTH(M_AXIMM_71_ARUSER_WIDTH),
        .M_AXIMM_72_ARUSER_WIDTH(M_AXIMM_72_ARUSER_WIDTH),
        .M_AXIMM_73_ARUSER_WIDTH(M_AXIMM_73_ARUSER_WIDTH),
        .M_AXIMM_74_ARUSER_WIDTH(M_AXIMM_74_ARUSER_WIDTH),
        .M_AXIMM_75_ARUSER_WIDTH(M_AXIMM_75_ARUSER_WIDTH),
        .M_AXIMM_76_ARUSER_WIDTH(M_AXIMM_76_ARUSER_WIDTH),
        .M_AXIMM_77_ARUSER_WIDTH(M_AXIMM_77_ARUSER_WIDTH),
        .M_AXIMM_78_ARUSER_WIDTH(M_AXIMM_78_ARUSER_WIDTH),
        .M_AXIMM_79_ARUSER_WIDTH(M_AXIMM_79_ARUSER_WIDTH),
        .M_AXIMM_80_ARUSER_WIDTH(M_AXIMM_80_ARUSER_WIDTH),
        .M_AXIMM_81_ARUSER_WIDTH(M_AXIMM_81_ARUSER_WIDTH),
        .M_AXIMM_82_ARUSER_WIDTH(M_AXIMM_82_ARUSER_WIDTH),
        .M_AXIMM_83_ARUSER_WIDTH(M_AXIMM_83_ARUSER_WIDTH),
        .M_AXIMM_84_ARUSER_WIDTH(M_AXIMM_84_ARUSER_WIDTH),
        .M_AXIMM_85_ARUSER_WIDTH(M_AXIMM_85_ARUSER_WIDTH),
        .M_AXIMM_86_ARUSER_WIDTH(M_AXIMM_86_ARUSER_WIDTH),
        .M_AXIMM_87_ARUSER_WIDTH(M_AXIMM_87_ARUSER_WIDTH),
        .M_AXIMM_88_ARUSER_WIDTH(M_AXIMM_88_ARUSER_WIDTH),
        .M_AXIMM_89_ARUSER_WIDTH(M_AXIMM_89_ARUSER_WIDTH),
        .M_AXIMM_90_ARUSER_WIDTH(M_AXIMM_90_ARUSER_WIDTH),
        .M_AXIMM_91_ARUSER_WIDTH(M_AXIMM_91_ARUSER_WIDTH),
        .M_AXIMM_92_ARUSER_WIDTH(M_AXIMM_92_ARUSER_WIDTH),
        .M_AXIMM_93_ARUSER_WIDTH(M_AXIMM_93_ARUSER_WIDTH),
        .M_AXIMM_94_ARUSER_WIDTH(M_AXIMM_94_ARUSER_WIDTH),
        .M_AXIMM_95_ARUSER_WIDTH(M_AXIMM_95_ARUSER_WIDTH),
        .M_AXIMM_96_ARUSER_WIDTH(M_AXIMM_96_ARUSER_WIDTH),
        .M_AXIMM_97_ARUSER_WIDTH(M_AXIMM_97_ARUSER_WIDTH),
        .M_AXIMM_98_ARUSER_WIDTH(M_AXIMM_98_ARUSER_WIDTH),
        .M_AXIMM_99_ARUSER_WIDTH(M_AXIMM_99_ARUSER_WIDTH),
        .M_AXIMM_100_ARUSER_WIDTH(M_AXIMM_100_ARUSER_WIDTH),
        .M_AXIMM_101_ARUSER_WIDTH(M_AXIMM_101_ARUSER_WIDTH),
        .M_AXIMM_102_ARUSER_WIDTH(M_AXIMM_102_ARUSER_WIDTH),
        .M_AXIMM_103_ARUSER_WIDTH(M_AXIMM_103_ARUSER_WIDTH),
        .M_AXIMM_104_ARUSER_WIDTH(M_AXIMM_104_ARUSER_WIDTH),
        .M_AXIMM_105_ARUSER_WIDTH(M_AXIMM_105_ARUSER_WIDTH),
        .M_AXIMM_106_ARUSER_WIDTH(M_AXIMM_106_ARUSER_WIDTH),
        .M_AXIMM_107_ARUSER_WIDTH(M_AXIMM_107_ARUSER_WIDTH),
        .M_AXIMM_108_ARUSER_WIDTH(M_AXIMM_108_ARUSER_WIDTH),
        .M_AXIMM_109_ARUSER_WIDTH(M_AXIMM_109_ARUSER_WIDTH),
        .M_AXIMM_110_ARUSER_WIDTH(M_AXIMM_110_ARUSER_WIDTH),
        .M_AXIMM_111_ARUSER_WIDTH(M_AXIMM_111_ARUSER_WIDTH),
        .M_AXIMM_112_ARUSER_WIDTH(M_AXIMM_112_ARUSER_WIDTH),
        .M_AXIMM_113_ARUSER_WIDTH(M_AXIMM_113_ARUSER_WIDTH),
        .M_AXIMM_114_ARUSER_WIDTH(M_AXIMM_114_ARUSER_WIDTH),
        .M_AXIMM_115_ARUSER_WIDTH(M_AXIMM_115_ARUSER_WIDTH),
        .M_AXIMM_116_ARUSER_WIDTH(M_AXIMM_116_ARUSER_WIDTH),
        .M_AXIMM_117_ARUSER_WIDTH(M_AXIMM_117_ARUSER_WIDTH),
        .M_AXIMM_118_ARUSER_WIDTH(M_AXIMM_118_ARUSER_WIDTH),
        .M_AXIMM_119_ARUSER_WIDTH(M_AXIMM_119_ARUSER_WIDTH),
        .M_AXIMM_120_ARUSER_WIDTH(M_AXIMM_120_ARUSER_WIDTH),
        .M_AXIMM_121_ARUSER_WIDTH(M_AXIMM_121_ARUSER_WIDTH),
        .M_AXIMM_122_ARUSER_WIDTH(M_AXIMM_122_ARUSER_WIDTH),
        .M_AXIMM_123_ARUSER_WIDTH(M_AXIMM_123_ARUSER_WIDTH),
        .M_AXIMM_124_ARUSER_WIDTH(M_AXIMM_124_ARUSER_WIDTH),
        .M_AXIMM_125_ARUSER_WIDTH(M_AXIMM_125_ARUSER_WIDTH),
        .M_AXIMM_126_ARUSER_WIDTH(M_AXIMM_126_ARUSER_WIDTH),
        .M_AXIMM_127_ARUSER_WIDTH(M_AXIMM_127_ARUSER_WIDTH),
        .M_AXIMM_0_AWUSER_WIDTH(M_AXIMM_0_AWUSER_WIDTH),
        .M_AXIMM_1_AWUSER_WIDTH(M_AXIMM_1_AWUSER_WIDTH),
        .M_AXIMM_2_AWUSER_WIDTH(M_AXIMM_2_AWUSER_WIDTH),
        .M_AXIMM_3_AWUSER_WIDTH(M_AXIMM_3_AWUSER_WIDTH),
        .M_AXIMM_4_AWUSER_WIDTH(M_AXIMM_4_AWUSER_WIDTH),
        .M_AXIMM_5_AWUSER_WIDTH(M_AXIMM_5_AWUSER_WIDTH),
        .M_AXIMM_6_AWUSER_WIDTH(M_AXIMM_6_AWUSER_WIDTH),
        .M_AXIMM_7_AWUSER_WIDTH(M_AXIMM_7_AWUSER_WIDTH),
        .M_AXIMM_8_AWUSER_WIDTH(M_AXIMM_8_AWUSER_WIDTH),
        .M_AXIMM_9_AWUSER_WIDTH(M_AXIMM_9_AWUSER_WIDTH),
        .M_AXIMM_10_AWUSER_WIDTH(M_AXIMM_10_AWUSER_WIDTH),
        .M_AXIMM_11_AWUSER_WIDTH(M_AXIMM_11_AWUSER_WIDTH),
        .M_AXIMM_12_AWUSER_WIDTH(M_AXIMM_12_AWUSER_WIDTH),
        .M_AXIMM_13_AWUSER_WIDTH(M_AXIMM_13_AWUSER_WIDTH),
        .M_AXIMM_14_AWUSER_WIDTH(M_AXIMM_14_AWUSER_WIDTH),
        .M_AXIMM_15_AWUSER_WIDTH(M_AXIMM_15_AWUSER_WIDTH),
        .M_AXIMM_16_AWUSER_WIDTH(M_AXIMM_16_AWUSER_WIDTH),
        .M_AXIMM_17_AWUSER_WIDTH(M_AXIMM_17_AWUSER_WIDTH),
        .M_AXIMM_18_AWUSER_WIDTH(M_AXIMM_18_AWUSER_WIDTH),
        .M_AXIMM_19_AWUSER_WIDTH(M_AXIMM_19_AWUSER_WIDTH),
        .M_AXIMM_20_AWUSER_WIDTH(M_AXIMM_20_AWUSER_WIDTH),
        .M_AXIMM_21_AWUSER_WIDTH(M_AXIMM_21_AWUSER_WIDTH),
        .M_AXIMM_22_AWUSER_WIDTH(M_AXIMM_22_AWUSER_WIDTH),
        .M_AXIMM_23_AWUSER_WIDTH(M_AXIMM_23_AWUSER_WIDTH),
        .M_AXIMM_24_AWUSER_WIDTH(M_AXIMM_24_AWUSER_WIDTH),
        .M_AXIMM_25_AWUSER_WIDTH(M_AXIMM_25_AWUSER_WIDTH),
        .M_AXIMM_26_AWUSER_WIDTH(M_AXIMM_26_AWUSER_WIDTH),
        .M_AXIMM_27_AWUSER_WIDTH(M_AXIMM_27_AWUSER_WIDTH),
        .M_AXIMM_28_AWUSER_WIDTH(M_AXIMM_28_AWUSER_WIDTH),
        .M_AXIMM_29_AWUSER_WIDTH(M_AXIMM_29_AWUSER_WIDTH),
        .M_AXIMM_30_AWUSER_WIDTH(M_AXIMM_30_AWUSER_WIDTH),
        .M_AXIMM_31_AWUSER_WIDTH(M_AXIMM_31_AWUSER_WIDTH),
        .M_AXIMM_32_AWUSER_WIDTH(M_AXIMM_32_AWUSER_WIDTH),
        .M_AXIMM_33_AWUSER_WIDTH(M_AXIMM_33_AWUSER_WIDTH),
        .M_AXIMM_34_AWUSER_WIDTH(M_AXIMM_34_AWUSER_WIDTH),
        .M_AXIMM_35_AWUSER_WIDTH(M_AXIMM_35_AWUSER_WIDTH),
        .M_AXIMM_36_AWUSER_WIDTH(M_AXIMM_36_AWUSER_WIDTH),
        .M_AXIMM_37_AWUSER_WIDTH(M_AXIMM_37_AWUSER_WIDTH),
        .M_AXIMM_38_AWUSER_WIDTH(M_AXIMM_38_AWUSER_WIDTH),
        .M_AXIMM_39_AWUSER_WIDTH(M_AXIMM_39_AWUSER_WIDTH),
        .M_AXIMM_40_AWUSER_WIDTH(M_AXIMM_40_AWUSER_WIDTH),
        .M_AXIMM_41_AWUSER_WIDTH(M_AXIMM_41_AWUSER_WIDTH),
        .M_AXIMM_42_AWUSER_WIDTH(M_AXIMM_42_AWUSER_WIDTH),
        .M_AXIMM_43_AWUSER_WIDTH(M_AXIMM_43_AWUSER_WIDTH),
        .M_AXIMM_44_AWUSER_WIDTH(M_AXIMM_44_AWUSER_WIDTH),
        .M_AXIMM_45_AWUSER_WIDTH(M_AXIMM_45_AWUSER_WIDTH),
        .M_AXIMM_46_AWUSER_WIDTH(M_AXIMM_46_AWUSER_WIDTH),
        .M_AXIMM_47_AWUSER_WIDTH(M_AXIMM_47_AWUSER_WIDTH),
        .M_AXIMM_48_AWUSER_WIDTH(M_AXIMM_48_AWUSER_WIDTH),
        .M_AXIMM_49_AWUSER_WIDTH(M_AXIMM_49_AWUSER_WIDTH),
        .M_AXIMM_50_AWUSER_WIDTH(M_AXIMM_50_AWUSER_WIDTH),
        .M_AXIMM_51_AWUSER_WIDTH(M_AXIMM_51_AWUSER_WIDTH),
        .M_AXIMM_52_AWUSER_WIDTH(M_AXIMM_52_AWUSER_WIDTH),
        .M_AXIMM_53_AWUSER_WIDTH(M_AXIMM_53_AWUSER_WIDTH),
        .M_AXIMM_54_AWUSER_WIDTH(M_AXIMM_54_AWUSER_WIDTH),
        .M_AXIMM_55_AWUSER_WIDTH(M_AXIMM_55_AWUSER_WIDTH),
        .M_AXIMM_56_AWUSER_WIDTH(M_AXIMM_56_AWUSER_WIDTH),
        .M_AXIMM_57_AWUSER_WIDTH(M_AXIMM_57_AWUSER_WIDTH),
        .M_AXIMM_58_AWUSER_WIDTH(M_AXIMM_58_AWUSER_WIDTH),
        .M_AXIMM_59_AWUSER_WIDTH(M_AXIMM_59_AWUSER_WIDTH),
        .M_AXIMM_60_AWUSER_WIDTH(M_AXIMM_60_AWUSER_WIDTH),
        .M_AXIMM_61_AWUSER_WIDTH(M_AXIMM_61_AWUSER_WIDTH),
        .M_AXIMM_62_AWUSER_WIDTH(M_AXIMM_62_AWUSER_WIDTH),
        .M_AXIMM_63_AWUSER_WIDTH(M_AXIMM_63_AWUSER_WIDTH),
        .M_AXIMM_64_AWUSER_WIDTH(M_AXIMM_64_AWUSER_WIDTH),
        .M_AXIMM_65_AWUSER_WIDTH(M_AXIMM_65_AWUSER_WIDTH),
        .M_AXIMM_66_AWUSER_WIDTH(M_AXIMM_66_AWUSER_WIDTH),
        .M_AXIMM_67_AWUSER_WIDTH(M_AXIMM_67_AWUSER_WIDTH),
        .M_AXIMM_68_AWUSER_WIDTH(M_AXIMM_68_AWUSER_WIDTH),
        .M_AXIMM_69_AWUSER_WIDTH(M_AXIMM_69_AWUSER_WIDTH),
        .M_AXIMM_70_AWUSER_WIDTH(M_AXIMM_70_AWUSER_WIDTH),
        .M_AXIMM_71_AWUSER_WIDTH(M_AXIMM_71_AWUSER_WIDTH),
        .M_AXIMM_72_AWUSER_WIDTH(M_AXIMM_72_AWUSER_WIDTH),
        .M_AXIMM_73_AWUSER_WIDTH(M_AXIMM_73_AWUSER_WIDTH),
        .M_AXIMM_74_AWUSER_WIDTH(M_AXIMM_74_AWUSER_WIDTH),
        .M_AXIMM_75_AWUSER_WIDTH(M_AXIMM_75_AWUSER_WIDTH),
        .M_AXIMM_76_AWUSER_WIDTH(M_AXIMM_76_AWUSER_WIDTH),
        .M_AXIMM_77_AWUSER_WIDTH(M_AXIMM_77_AWUSER_WIDTH),
        .M_AXIMM_78_AWUSER_WIDTH(M_AXIMM_78_AWUSER_WIDTH),
        .M_AXIMM_79_AWUSER_WIDTH(M_AXIMM_79_AWUSER_WIDTH),
        .M_AXIMM_80_AWUSER_WIDTH(M_AXIMM_80_AWUSER_WIDTH),
        .M_AXIMM_81_AWUSER_WIDTH(M_AXIMM_81_AWUSER_WIDTH),
        .M_AXIMM_82_AWUSER_WIDTH(M_AXIMM_82_AWUSER_WIDTH),
        .M_AXIMM_83_AWUSER_WIDTH(M_AXIMM_83_AWUSER_WIDTH),
        .M_AXIMM_84_AWUSER_WIDTH(M_AXIMM_84_AWUSER_WIDTH),
        .M_AXIMM_85_AWUSER_WIDTH(M_AXIMM_85_AWUSER_WIDTH),
        .M_AXIMM_86_AWUSER_WIDTH(M_AXIMM_86_AWUSER_WIDTH),
        .M_AXIMM_87_AWUSER_WIDTH(M_AXIMM_87_AWUSER_WIDTH),
        .M_AXIMM_88_AWUSER_WIDTH(M_AXIMM_88_AWUSER_WIDTH),
        .M_AXIMM_89_AWUSER_WIDTH(M_AXIMM_89_AWUSER_WIDTH),
        .M_AXIMM_90_AWUSER_WIDTH(M_AXIMM_90_AWUSER_WIDTH),
        .M_AXIMM_91_AWUSER_WIDTH(M_AXIMM_91_AWUSER_WIDTH),
        .M_AXIMM_92_AWUSER_WIDTH(M_AXIMM_92_AWUSER_WIDTH),
        .M_AXIMM_93_AWUSER_WIDTH(M_AXIMM_93_AWUSER_WIDTH),
        .M_AXIMM_94_AWUSER_WIDTH(M_AXIMM_94_AWUSER_WIDTH),
        .M_AXIMM_95_AWUSER_WIDTH(M_AXIMM_95_AWUSER_WIDTH),
        .M_AXIMM_96_AWUSER_WIDTH(M_AXIMM_96_AWUSER_WIDTH),
        .M_AXIMM_97_AWUSER_WIDTH(M_AXIMM_97_AWUSER_WIDTH),
        .M_AXIMM_98_AWUSER_WIDTH(M_AXIMM_98_AWUSER_WIDTH),
        .M_AXIMM_99_AWUSER_WIDTH(M_AXIMM_99_AWUSER_WIDTH),
        .M_AXIMM_100_AWUSER_WIDTH(M_AXIMM_100_AWUSER_WIDTH),
        .M_AXIMM_101_AWUSER_WIDTH(M_AXIMM_101_AWUSER_WIDTH),
        .M_AXIMM_102_AWUSER_WIDTH(M_AXIMM_102_AWUSER_WIDTH),
        .M_AXIMM_103_AWUSER_WIDTH(M_AXIMM_103_AWUSER_WIDTH),
        .M_AXIMM_104_AWUSER_WIDTH(M_AXIMM_104_AWUSER_WIDTH),
        .M_AXIMM_105_AWUSER_WIDTH(M_AXIMM_105_AWUSER_WIDTH),
        .M_AXIMM_106_AWUSER_WIDTH(M_AXIMM_106_AWUSER_WIDTH),
        .M_AXIMM_107_AWUSER_WIDTH(M_AXIMM_107_AWUSER_WIDTH),
        .M_AXIMM_108_AWUSER_WIDTH(M_AXIMM_108_AWUSER_WIDTH),
        .M_AXIMM_109_AWUSER_WIDTH(M_AXIMM_109_AWUSER_WIDTH),
        .M_AXIMM_110_AWUSER_WIDTH(M_AXIMM_110_AWUSER_WIDTH),
        .M_AXIMM_111_AWUSER_WIDTH(M_AXIMM_111_AWUSER_WIDTH),
        .M_AXIMM_112_AWUSER_WIDTH(M_AXIMM_112_AWUSER_WIDTH),
        .M_AXIMM_113_AWUSER_WIDTH(M_AXIMM_113_AWUSER_WIDTH),
        .M_AXIMM_114_AWUSER_WIDTH(M_AXIMM_114_AWUSER_WIDTH),
        .M_AXIMM_115_AWUSER_WIDTH(M_AXIMM_115_AWUSER_WIDTH),
        .M_AXIMM_116_AWUSER_WIDTH(M_AXIMM_116_AWUSER_WIDTH),
        .M_AXIMM_117_AWUSER_WIDTH(M_AXIMM_117_AWUSER_WIDTH),
        .M_AXIMM_118_AWUSER_WIDTH(M_AXIMM_118_AWUSER_WIDTH),
        .M_AXIMM_119_AWUSER_WIDTH(M_AXIMM_119_AWUSER_WIDTH),
        .M_AXIMM_120_AWUSER_WIDTH(M_AXIMM_120_AWUSER_WIDTH),
        .M_AXIMM_121_AWUSER_WIDTH(M_AXIMM_121_AWUSER_WIDTH),
        .M_AXIMM_122_AWUSER_WIDTH(M_AXIMM_122_AWUSER_WIDTH),
        .M_AXIMM_123_AWUSER_WIDTH(M_AXIMM_123_AWUSER_WIDTH),
        .M_AXIMM_124_AWUSER_WIDTH(M_AXIMM_124_AWUSER_WIDTH),
        .M_AXIMM_125_AWUSER_WIDTH(M_AXIMM_125_AWUSER_WIDTH),
        .M_AXIMM_126_AWUSER_WIDTH(M_AXIMM_126_AWUSER_WIDTH),
        .M_AXIMM_127_AWUSER_WIDTH(M_AXIMM_127_AWUSER_WIDTH),
        .M_AXIMM_0_WUSER_WIDTH(M_AXIMM_0_WUSER_WIDTH),
        .M_AXIMM_1_WUSER_WIDTH(M_AXIMM_1_WUSER_WIDTH),
        .M_AXIMM_2_WUSER_WIDTH(M_AXIMM_2_WUSER_WIDTH),
        .M_AXIMM_3_WUSER_WIDTH(M_AXIMM_3_WUSER_WIDTH),
        .M_AXIMM_4_WUSER_WIDTH(M_AXIMM_4_WUSER_WIDTH),
        .M_AXIMM_5_WUSER_WIDTH(M_AXIMM_5_WUSER_WIDTH),
        .M_AXIMM_6_WUSER_WIDTH(M_AXIMM_6_WUSER_WIDTH),
        .M_AXIMM_7_WUSER_WIDTH(M_AXIMM_7_WUSER_WIDTH),
        .M_AXIMM_8_WUSER_WIDTH(M_AXIMM_8_WUSER_WIDTH),
        .M_AXIMM_9_WUSER_WIDTH(M_AXIMM_9_WUSER_WIDTH),
        .M_AXIMM_10_WUSER_WIDTH(M_AXIMM_10_WUSER_WIDTH),
        .M_AXIMM_11_WUSER_WIDTH(M_AXIMM_11_WUSER_WIDTH),
        .M_AXIMM_12_WUSER_WIDTH(M_AXIMM_12_WUSER_WIDTH),
        .M_AXIMM_13_WUSER_WIDTH(M_AXIMM_13_WUSER_WIDTH),
        .M_AXIMM_14_WUSER_WIDTH(M_AXIMM_14_WUSER_WIDTH),
        .M_AXIMM_15_WUSER_WIDTH(M_AXIMM_15_WUSER_WIDTH),
        .M_AXIMM_16_WUSER_WIDTH(M_AXIMM_16_WUSER_WIDTH),
        .M_AXIMM_17_WUSER_WIDTH(M_AXIMM_17_WUSER_WIDTH),
        .M_AXIMM_18_WUSER_WIDTH(M_AXIMM_18_WUSER_WIDTH),
        .M_AXIMM_19_WUSER_WIDTH(M_AXIMM_19_WUSER_WIDTH),
        .M_AXIMM_20_WUSER_WIDTH(M_AXIMM_20_WUSER_WIDTH),
        .M_AXIMM_21_WUSER_WIDTH(M_AXIMM_21_WUSER_WIDTH),
        .M_AXIMM_22_WUSER_WIDTH(M_AXIMM_22_WUSER_WIDTH),
        .M_AXIMM_23_WUSER_WIDTH(M_AXIMM_23_WUSER_WIDTH),
        .M_AXIMM_24_WUSER_WIDTH(M_AXIMM_24_WUSER_WIDTH),
        .M_AXIMM_25_WUSER_WIDTH(M_AXIMM_25_WUSER_WIDTH),
        .M_AXIMM_26_WUSER_WIDTH(M_AXIMM_26_WUSER_WIDTH),
        .M_AXIMM_27_WUSER_WIDTH(M_AXIMM_27_WUSER_WIDTH),
        .M_AXIMM_28_WUSER_WIDTH(M_AXIMM_28_WUSER_WIDTH),
        .M_AXIMM_29_WUSER_WIDTH(M_AXIMM_29_WUSER_WIDTH),
        .M_AXIMM_30_WUSER_WIDTH(M_AXIMM_30_WUSER_WIDTH),
        .M_AXIMM_31_WUSER_WIDTH(M_AXIMM_31_WUSER_WIDTH),
        .M_AXIMM_32_WUSER_WIDTH(M_AXIMM_32_WUSER_WIDTH),
        .M_AXIMM_33_WUSER_WIDTH(M_AXIMM_33_WUSER_WIDTH),
        .M_AXIMM_34_WUSER_WIDTH(M_AXIMM_34_WUSER_WIDTH),
        .M_AXIMM_35_WUSER_WIDTH(M_AXIMM_35_WUSER_WIDTH),
        .M_AXIMM_36_WUSER_WIDTH(M_AXIMM_36_WUSER_WIDTH),
        .M_AXIMM_37_WUSER_WIDTH(M_AXIMM_37_WUSER_WIDTH),
        .M_AXIMM_38_WUSER_WIDTH(M_AXIMM_38_WUSER_WIDTH),
        .M_AXIMM_39_WUSER_WIDTH(M_AXIMM_39_WUSER_WIDTH),
        .M_AXIMM_40_WUSER_WIDTH(M_AXIMM_40_WUSER_WIDTH),
        .M_AXIMM_41_WUSER_WIDTH(M_AXIMM_41_WUSER_WIDTH),
        .M_AXIMM_42_WUSER_WIDTH(M_AXIMM_42_WUSER_WIDTH),
        .M_AXIMM_43_WUSER_WIDTH(M_AXIMM_43_WUSER_WIDTH),
        .M_AXIMM_44_WUSER_WIDTH(M_AXIMM_44_WUSER_WIDTH),
        .M_AXIMM_45_WUSER_WIDTH(M_AXIMM_45_WUSER_WIDTH),
        .M_AXIMM_46_WUSER_WIDTH(M_AXIMM_46_WUSER_WIDTH),
        .M_AXIMM_47_WUSER_WIDTH(M_AXIMM_47_WUSER_WIDTH),
        .M_AXIMM_48_WUSER_WIDTH(M_AXIMM_48_WUSER_WIDTH),
        .M_AXIMM_49_WUSER_WIDTH(M_AXIMM_49_WUSER_WIDTH),
        .M_AXIMM_50_WUSER_WIDTH(M_AXIMM_50_WUSER_WIDTH),
        .M_AXIMM_51_WUSER_WIDTH(M_AXIMM_51_WUSER_WIDTH),
        .M_AXIMM_52_WUSER_WIDTH(M_AXIMM_52_WUSER_WIDTH),
        .M_AXIMM_53_WUSER_WIDTH(M_AXIMM_53_WUSER_WIDTH),
        .M_AXIMM_54_WUSER_WIDTH(M_AXIMM_54_WUSER_WIDTH),
        .M_AXIMM_55_WUSER_WIDTH(M_AXIMM_55_WUSER_WIDTH),
        .M_AXIMM_56_WUSER_WIDTH(M_AXIMM_56_WUSER_WIDTH),
        .M_AXIMM_57_WUSER_WIDTH(M_AXIMM_57_WUSER_WIDTH),
        .M_AXIMM_58_WUSER_WIDTH(M_AXIMM_58_WUSER_WIDTH),
        .M_AXIMM_59_WUSER_WIDTH(M_AXIMM_59_WUSER_WIDTH),
        .M_AXIMM_60_WUSER_WIDTH(M_AXIMM_60_WUSER_WIDTH),
        .M_AXIMM_61_WUSER_WIDTH(M_AXIMM_61_WUSER_WIDTH),
        .M_AXIMM_62_WUSER_WIDTH(M_AXIMM_62_WUSER_WIDTH),
        .M_AXIMM_63_WUSER_WIDTH(M_AXIMM_63_WUSER_WIDTH),
        .M_AXIMM_64_WUSER_WIDTH(M_AXIMM_64_WUSER_WIDTH),
        .M_AXIMM_65_WUSER_WIDTH(M_AXIMM_65_WUSER_WIDTH),
        .M_AXIMM_66_WUSER_WIDTH(M_AXIMM_66_WUSER_WIDTH),
        .M_AXIMM_67_WUSER_WIDTH(M_AXIMM_67_WUSER_WIDTH),
        .M_AXIMM_68_WUSER_WIDTH(M_AXIMM_68_WUSER_WIDTH),
        .M_AXIMM_69_WUSER_WIDTH(M_AXIMM_69_WUSER_WIDTH),
        .M_AXIMM_70_WUSER_WIDTH(M_AXIMM_70_WUSER_WIDTH),
        .M_AXIMM_71_WUSER_WIDTH(M_AXIMM_71_WUSER_WIDTH),
        .M_AXIMM_72_WUSER_WIDTH(M_AXIMM_72_WUSER_WIDTH),
        .M_AXIMM_73_WUSER_WIDTH(M_AXIMM_73_WUSER_WIDTH),
        .M_AXIMM_74_WUSER_WIDTH(M_AXIMM_74_WUSER_WIDTH),
        .M_AXIMM_75_WUSER_WIDTH(M_AXIMM_75_WUSER_WIDTH),
        .M_AXIMM_76_WUSER_WIDTH(M_AXIMM_76_WUSER_WIDTH),
        .M_AXIMM_77_WUSER_WIDTH(M_AXIMM_77_WUSER_WIDTH),
        .M_AXIMM_78_WUSER_WIDTH(M_AXIMM_78_WUSER_WIDTH),
        .M_AXIMM_79_WUSER_WIDTH(M_AXIMM_79_WUSER_WIDTH),
        .M_AXIMM_80_WUSER_WIDTH(M_AXIMM_80_WUSER_WIDTH),
        .M_AXIMM_81_WUSER_WIDTH(M_AXIMM_81_WUSER_WIDTH),
        .M_AXIMM_82_WUSER_WIDTH(M_AXIMM_82_WUSER_WIDTH),
        .M_AXIMM_83_WUSER_WIDTH(M_AXIMM_83_WUSER_WIDTH),
        .M_AXIMM_84_WUSER_WIDTH(M_AXIMM_84_WUSER_WIDTH),
        .M_AXIMM_85_WUSER_WIDTH(M_AXIMM_85_WUSER_WIDTH),
        .M_AXIMM_86_WUSER_WIDTH(M_AXIMM_86_WUSER_WIDTH),
        .M_AXIMM_87_WUSER_WIDTH(M_AXIMM_87_WUSER_WIDTH),
        .M_AXIMM_88_WUSER_WIDTH(M_AXIMM_88_WUSER_WIDTH),
        .M_AXIMM_89_WUSER_WIDTH(M_AXIMM_89_WUSER_WIDTH),
        .M_AXIMM_90_WUSER_WIDTH(M_AXIMM_90_WUSER_WIDTH),
        .M_AXIMM_91_WUSER_WIDTH(M_AXIMM_91_WUSER_WIDTH),
        .M_AXIMM_92_WUSER_WIDTH(M_AXIMM_92_WUSER_WIDTH),
        .M_AXIMM_93_WUSER_WIDTH(M_AXIMM_93_WUSER_WIDTH),
        .M_AXIMM_94_WUSER_WIDTH(M_AXIMM_94_WUSER_WIDTH),
        .M_AXIMM_95_WUSER_WIDTH(M_AXIMM_95_WUSER_WIDTH),
        .M_AXIMM_96_WUSER_WIDTH(M_AXIMM_96_WUSER_WIDTH),
        .M_AXIMM_97_WUSER_WIDTH(M_AXIMM_97_WUSER_WIDTH),
        .M_AXIMM_98_WUSER_WIDTH(M_AXIMM_98_WUSER_WIDTH),
        .M_AXIMM_99_WUSER_WIDTH(M_AXIMM_99_WUSER_WIDTH),
        .M_AXIMM_100_WUSER_WIDTH(M_AXIMM_100_WUSER_WIDTH),
        .M_AXIMM_101_WUSER_WIDTH(M_AXIMM_101_WUSER_WIDTH),
        .M_AXIMM_102_WUSER_WIDTH(M_AXIMM_102_WUSER_WIDTH),
        .M_AXIMM_103_WUSER_WIDTH(M_AXIMM_103_WUSER_WIDTH),
        .M_AXIMM_104_WUSER_WIDTH(M_AXIMM_104_WUSER_WIDTH),
        .M_AXIMM_105_WUSER_WIDTH(M_AXIMM_105_WUSER_WIDTH),
        .M_AXIMM_106_WUSER_WIDTH(M_AXIMM_106_WUSER_WIDTH),
        .M_AXIMM_107_WUSER_WIDTH(M_AXIMM_107_WUSER_WIDTH),
        .M_AXIMM_108_WUSER_WIDTH(M_AXIMM_108_WUSER_WIDTH),
        .M_AXIMM_109_WUSER_WIDTH(M_AXIMM_109_WUSER_WIDTH),
        .M_AXIMM_110_WUSER_WIDTH(M_AXIMM_110_WUSER_WIDTH),
        .M_AXIMM_111_WUSER_WIDTH(M_AXIMM_111_WUSER_WIDTH),
        .M_AXIMM_112_WUSER_WIDTH(M_AXIMM_112_WUSER_WIDTH),
        .M_AXIMM_113_WUSER_WIDTH(M_AXIMM_113_WUSER_WIDTH),
        .M_AXIMM_114_WUSER_WIDTH(M_AXIMM_114_WUSER_WIDTH),
        .M_AXIMM_115_WUSER_WIDTH(M_AXIMM_115_WUSER_WIDTH),
        .M_AXIMM_116_WUSER_WIDTH(M_AXIMM_116_WUSER_WIDTH),
        .M_AXIMM_117_WUSER_WIDTH(M_AXIMM_117_WUSER_WIDTH),
        .M_AXIMM_118_WUSER_WIDTH(M_AXIMM_118_WUSER_WIDTH),
        .M_AXIMM_119_WUSER_WIDTH(M_AXIMM_119_WUSER_WIDTH),
        .M_AXIMM_120_WUSER_WIDTH(M_AXIMM_120_WUSER_WIDTH),
        .M_AXIMM_121_WUSER_WIDTH(M_AXIMM_121_WUSER_WIDTH),
        .M_AXIMM_122_WUSER_WIDTH(M_AXIMM_122_WUSER_WIDTH),
        .M_AXIMM_123_WUSER_WIDTH(M_AXIMM_123_WUSER_WIDTH),
        .M_AXIMM_124_WUSER_WIDTH(M_AXIMM_124_WUSER_WIDTH),
        .M_AXIMM_125_WUSER_WIDTH(M_AXIMM_125_WUSER_WIDTH),
        .M_AXIMM_126_WUSER_WIDTH(M_AXIMM_126_WUSER_WIDTH),
        .M_AXIMM_127_WUSER_WIDTH(M_AXIMM_127_WUSER_WIDTH),
        .M_AXIMM_0_BUSER_WIDTH(M_AXIMM_0_BUSER_WIDTH),
        .M_AXIMM_1_BUSER_WIDTH(M_AXIMM_1_BUSER_WIDTH),
        .M_AXIMM_2_BUSER_WIDTH(M_AXIMM_2_BUSER_WIDTH),
        .M_AXIMM_3_BUSER_WIDTH(M_AXIMM_3_BUSER_WIDTH),
        .M_AXIMM_4_BUSER_WIDTH(M_AXIMM_4_BUSER_WIDTH),
        .M_AXIMM_5_BUSER_WIDTH(M_AXIMM_5_BUSER_WIDTH),
        .M_AXIMM_6_BUSER_WIDTH(M_AXIMM_6_BUSER_WIDTH),
        .M_AXIMM_7_BUSER_WIDTH(M_AXIMM_7_BUSER_WIDTH),
        .M_AXIMM_8_BUSER_WIDTH(M_AXIMM_8_BUSER_WIDTH),
        .M_AXIMM_9_BUSER_WIDTH(M_AXIMM_9_BUSER_WIDTH),
        .M_AXIMM_10_BUSER_WIDTH(M_AXIMM_10_BUSER_WIDTH),
        .M_AXIMM_11_BUSER_WIDTH(M_AXIMM_11_BUSER_WIDTH),
        .M_AXIMM_12_BUSER_WIDTH(M_AXIMM_12_BUSER_WIDTH),
        .M_AXIMM_13_BUSER_WIDTH(M_AXIMM_13_BUSER_WIDTH),
        .M_AXIMM_14_BUSER_WIDTH(M_AXIMM_14_BUSER_WIDTH),
        .M_AXIMM_15_BUSER_WIDTH(M_AXIMM_15_BUSER_WIDTH),
        .M_AXIMM_16_BUSER_WIDTH(M_AXIMM_16_BUSER_WIDTH),
        .M_AXIMM_17_BUSER_WIDTH(M_AXIMM_17_BUSER_WIDTH),
        .M_AXIMM_18_BUSER_WIDTH(M_AXIMM_18_BUSER_WIDTH),
        .M_AXIMM_19_BUSER_WIDTH(M_AXIMM_19_BUSER_WIDTH),
        .M_AXIMM_20_BUSER_WIDTH(M_AXIMM_20_BUSER_WIDTH),
        .M_AXIMM_21_BUSER_WIDTH(M_AXIMM_21_BUSER_WIDTH),
        .M_AXIMM_22_BUSER_WIDTH(M_AXIMM_22_BUSER_WIDTH),
        .M_AXIMM_23_BUSER_WIDTH(M_AXIMM_23_BUSER_WIDTH),
        .M_AXIMM_24_BUSER_WIDTH(M_AXIMM_24_BUSER_WIDTH),
        .M_AXIMM_25_BUSER_WIDTH(M_AXIMM_25_BUSER_WIDTH),
        .M_AXIMM_26_BUSER_WIDTH(M_AXIMM_26_BUSER_WIDTH),
        .M_AXIMM_27_BUSER_WIDTH(M_AXIMM_27_BUSER_WIDTH),
        .M_AXIMM_28_BUSER_WIDTH(M_AXIMM_28_BUSER_WIDTH),
        .M_AXIMM_29_BUSER_WIDTH(M_AXIMM_29_BUSER_WIDTH),
        .M_AXIMM_30_BUSER_WIDTH(M_AXIMM_30_BUSER_WIDTH),
        .M_AXIMM_31_BUSER_WIDTH(M_AXIMM_31_BUSER_WIDTH),
        .M_AXIMM_32_BUSER_WIDTH(M_AXIMM_32_BUSER_WIDTH),
        .M_AXIMM_33_BUSER_WIDTH(M_AXIMM_33_BUSER_WIDTH),
        .M_AXIMM_34_BUSER_WIDTH(M_AXIMM_34_BUSER_WIDTH),
        .M_AXIMM_35_BUSER_WIDTH(M_AXIMM_35_BUSER_WIDTH),
        .M_AXIMM_36_BUSER_WIDTH(M_AXIMM_36_BUSER_WIDTH),
        .M_AXIMM_37_BUSER_WIDTH(M_AXIMM_37_BUSER_WIDTH),
        .M_AXIMM_38_BUSER_WIDTH(M_AXIMM_38_BUSER_WIDTH),
        .M_AXIMM_39_BUSER_WIDTH(M_AXIMM_39_BUSER_WIDTH),
        .M_AXIMM_40_BUSER_WIDTH(M_AXIMM_40_BUSER_WIDTH),
        .M_AXIMM_41_BUSER_WIDTH(M_AXIMM_41_BUSER_WIDTH),
        .M_AXIMM_42_BUSER_WIDTH(M_AXIMM_42_BUSER_WIDTH),
        .M_AXIMM_43_BUSER_WIDTH(M_AXIMM_43_BUSER_WIDTH),
        .M_AXIMM_44_BUSER_WIDTH(M_AXIMM_44_BUSER_WIDTH),
        .M_AXIMM_45_BUSER_WIDTH(M_AXIMM_45_BUSER_WIDTH),
        .M_AXIMM_46_BUSER_WIDTH(M_AXIMM_46_BUSER_WIDTH),
        .M_AXIMM_47_BUSER_WIDTH(M_AXIMM_47_BUSER_WIDTH),
        .M_AXIMM_48_BUSER_WIDTH(M_AXIMM_48_BUSER_WIDTH),
        .M_AXIMM_49_BUSER_WIDTH(M_AXIMM_49_BUSER_WIDTH),
        .M_AXIMM_50_BUSER_WIDTH(M_AXIMM_50_BUSER_WIDTH),
        .M_AXIMM_51_BUSER_WIDTH(M_AXIMM_51_BUSER_WIDTH),
        .M_AXIMM_52_BUSER_WIDTH(M_AXIMM_52_BUSER_WIDTH),
        .M_AXIMM_53_BUSER_WIDTH(M_AXIMM_53_BUSER_WIDTH),
        .M_AXIMM_54_BUSER_WIDTH(M_AXIMM_54_BUSER_WIDTH),
        .M_AXIMM_55_BUSER_WIDTH(M_AXIMM_55_BUSER_WIDTH),
        .M_AXIMM_56_BUSER_WIDTH(M_AXIMM_56_BUSER_WIDTH),
        .M_AXIMM_57_BUSER_WIDTH(M_AXIMM_57_BUSER_WIDTH),
        .M_AXIMM_58_BUSER_WIDTH(M_AXIMM_58_BUSER_WIDTH),
        .M_AXIMM_59_BUSER_WIDTH(M_AXIMM_59_BUSER_WIDTH),
        .M_AXIMM_60_BUSER_WIDTH(M_AXIMM_60_BUSER_WIDTH),
        .M_AXIMM_61_BUSER_WIDTH(M_AXIMM_61_BUSER_WIDTH),
        .M_AXIMM_62_BUSER_WIDTH(M_AXIMM_62_BUSER_WIDTH),
        .M_AXIMM_63_BUSER_WIDTH(M_AXIMM_63_BUSER_WIDTH),
        .M_AXIMM_64_BUSER_WIDTH(M_AXIMM_64_BUSER_WIDTH),
        .M_AXIMM_65_BUSER_WIDTH(M_AXIMM_65_BUSER_WIDTH),
        .M_AXIMM_66_BUSER_WIDTH(M_AXIMM_66_BUSER_WIDTH),
        .M_AXIMM_67_BUSER_WIDTH(M_AXIMM_67_BUSER_WIDTH),
        .M_AXIMM_68_BUSER_WIDTH(M_AXIMM_68_BUSER_WIDTH),
        .M_AXIMM_69_BUSER_WIDTH(M_AXIMM_69_BUSER_WIDTH),
        .M_AXIMM_70_BUSER_WIDTH(M_AXIMM_70_BUSER_WIDTH),
        .M_AXIMM_71_BUSER_WIDTH(M_AXIMM_71_BUSER_WIDTH),
        .M_AXIMM_72_BUSER_WIDTH(M_AXIMM_72_BUSER_WIDTH),
        .M_AXIMM_73_BUSER_WIDTH(M_AXIMM_73_BUSER_WIDTH),
        .M_AXIMM_74_BUSER_WIDTH(M_AXIMM_74_BUSER_WIDTH),
        .M_AXIMM_75_BUSER_WIDTH(M_AXIMM_75_BUSER_WIDTH),
        .M_AXIMM_76_BUSER_WIDTH(M_AXIMM_76_BUSER_WIDTH),
        .M_AXIMM_77_BUSER_WIDTH(M_AXIMM_77_BUSER_WIDTH),
        .M_AXIMM_78_BUSER_WIDTH(M_AXIMM_78_BUSER_WIDTH),
        .M_AXIMM_79_BUSER_WIDTH(M_AXIMM_79_BUSER_WIDTH),
        .M_AXIMM_80_BUSER_WIDTH(M_AXIMM_80_BUSER_WIDTH),
        .M_AXIMM_81_BUSER_WIDTH(M_AXIMM_81_BUSER_WIDTH),
        .M_AXIMM_82_BUSER_WIDTH(M_AXIMM_82_BUSER_WIDTH),
        .M_AXIMM_83_BUSER_WIDTH(M_AXIMM_83_BUSER_WIDTH),
        .M_AXIMM_84_BUSER_WIDTH(M_AXIMM_84_BUSER_WIDTH),
        .M_AXIMM_85_BUSER_WIDTH(M_AXIMM_85_BUSER_WIDTH),
        .M_AXIMM_86_BUSER_WIDTH(M_AXIMM_86_BUSER_WIDTH),
        .M_AXIMM_87_BUSER_WIDTH(M_AXIMM_87_BUSER_WIDTH),
        .M_AXIMM_88_BUSER_WIDTH(M_AXIMM_88_BUSER_WIDTH),
        .M_AXIMM_89_BUSER_WIDTH(M_AXIMM_89_BUSER_WIDTH),
        .M_AXIMM_90_BUSER_WIDTH(M_AXIMM_90_BUSER_WIDTH),
        .M_AXIMM_91_BUSER_WIDTH(M_AXIMM_91_BUSER_WIDTH),
        .M_AXIMM_92_BUSER_WIDTH(M_AXIMM_92_BUSER_WIDTH),
        .M_AXIMM_93_BUSER_WIDTH(M_AXIMM_93_BUSER_WIDTH),
        .M_AXIMM_94_BUSER_WIDTH(M_AXIMM_94_BUSER_WIDTH),
        .M_AXIMM_95_BUSER_WIDTH(M_AXIMM_95_BUSER_WIDTH),
        .M_AXIMM_96_BUSER_WIDTH(M_AXIMM_96_BUSER_WIDTH),
        .M_AXIMM_97_BUSER_WIDTH(M_AXIMM_97_BUSER_WIDTH),
        .M_AXIMM_98_BUSER_WIDTH(M_AXIMM_98_BUSER_WIDTH),
        .M_AXIMM_99_BUSER_WIDTH(M_AXIMM_99_BUSER_WIDTH),
        .M_AXIMM_100_BUSER_WIDTH(M_AXIMM_100_BUSER_WIDTH),
        .M_AXIMM_101_BUSER_WIDTH(M_AXIMM_101_BUSER_WIDTH),
        .M_AXIMM_102_BUSER_WIDTH(M_AXIMM_102_BUSER_WIDTH),
        .M_AXIMM_103_BUSER_WIDTH(M_AXIMM_103_BUSER_WIDTH),
        .M_AXIMM_104_BUSER_WIDTH(M_AXIMM_104_BUSER_WIDTH),
        .M_AXIMM_105_BUSER_WIDTH(M_AXIMM_105_BUSER_WIDTH),
        .M_AXIMM_106_BUSER_WIDTH(M_AXIMM_106_BUSER_WIDTH),
        .M_AXIMM_107_BUSER_WIDTH(M_AXIMM_107_BUSER_WIDTH),
        .M_AXIMM_108_BUSER_WIDTH(M_AXIMM_108_BUSER_WIDTH),
        .M_AXIMM_109_BUSER_WIDTH(M_AXIMM_109_BUSER_WIDTH),
        .M_AXIMM_110_BUSER_WIDTH(M_AXIMM_110_BUSER_WIDTH),
        .M_AXIMM_111_BUSER_WIDTH(M_AXIMM_111_BUSER_WIDTH),
        .M_AXIMM_112_BUSER_WIDTH(M_AXIMM_112_BUSER_WIDTH),
        .M_AXIMM_113_BUSER_WIDTH(M_AXIMM_113_BUSER_WIDTH),
        .M_AXIMM_114_BUSER_WIDTH(M_AXIMM_114_BUSER_WIDTH),
        .M_AXIMM_115_BUSER_WIDTH(M_AXIMM_115_BUSER_WIDTH),
        .M_AXIMM_116_BUSER_WIDTH(M_AXIMM_116_BUSER_WIDTH),
        .M_AXIMM_117_BUSER_WIDTH(M_AXIMM_117_BUSER_WIDTH),
        .M_AXIMM_118_BUSER_WIDTH(M_AXIMM_118_BUSER_WIDTH),
        .M_AXIMM_119_BUSER_WIDTH(M_AXIMM_119_BUSER_WIDTH),
        .M_AXIMM_120_BUSER_WIDTH(M_AXIMM_120_BUSER_WIDTH),
        .M_AXIMM_121_BUSER_WIDTH(M_AXIMM_121_BUSER_WIDTH),
        .M_AXIMM_122_BUSER_WIDTH(M_AXIMM_122_BUSER_WIDTH),
        .M_AXIMM_123_BUSER_WIDTH(M_AXIMM_123_BUSER_WIDTH),
        .M_AXIMM_124_BUSER_WIDTH(M_AXIMM_124_BUSER_WIDTH),
        .M_AXIMM_125_BUSER_WIDTH(M_AXIMM_125_BUSER_WIDTH),
        .M_AXIMM_126_BUSER_WIDTH(M_AXIMM_126_BUSER_WIDTH),
        .M_AXIMM_127_BUSER_WIDTH(M_AXIMM_127_BUSER_WIDTH),
        .M_AXIMM_0_RUSER_WIDTH(M_AXIMM_0_RUSER_WIDTH),
        .M_AXIMM_1_RUSER_WIDTH(M_AXIMM_1_RUSER_WIDTH),
        .M_AXIMM_2_RUSER_WIDTH(M_AXIMM_2_RUSER_WIDTH),
        .M_AXIMM_3_RUSER_WIDTH(M_AXIMM_3_RUSER_WIDTH),
        .M_AXIMM_4_RUSER_WIDTH(M_AXIMM_4_RUSER_WIDTH),
        .M_AXIMM_5_RUSER_WIDTH(M_AXIMM_5_RUSER_WIDTH),
        .M_AXIMM_6_RUSER_WIDTH(M_AXIMM_6_RUSER_WIDTH),
        .M_AXIMM_7_RUSER_WIDTH(M_AXIMM_7_RUSER_WIDTH),
        .M_AXIMM_8_RUSER_WIDTH(M_AXIMM_8_RUSER_WIDTH),
        .M_AXIMM_9_RUSER_WIDTH(M_AXIMM_9_RUSER_WIDTH),
        .M_AXIMM_10_RUSER_WIDTH(M_AXIMM_10_RUSER_WIDTH),
        .M_AXIMM_11_RUSER_WIDTH(M_AXIMM_11_RUSER_WIDTH),
        .M_AXIMM_12_RUSER_WIDTH(M_AXIMM_12_RUSER_WIDTH),
        .M_AXIMM_13_RUSER_WIDTH(M_AXIMM_13_RUSER_WIDTH),
        .M_AXIMM_14_RUSER_WIDTH(M_AXIMM_14_RUSER_WIDTH),
        .M_AXIMM_15_RUSER_WIDTH(M_AXIMM_15_RUSER_WIDTH),
        .M_AXIMM_16_RUSER_WIDTH(M_AXIMM_16_RUSER_WIDTH),
        .M_AXIMM_17_RUSER_WIDTH(M_AXIMM_17_RUSER_WIDTH),
        .M_AXIMM_18_RUSER_WIDTH(M_AXIMM_18_RUSER_WIDTH),
        .M_AXIMM_19_RUSER_WIDTH(M_AXIMM_19_RUSER_WIDTH),
        .M_AXIMM_20_RUSER_WIDTH(M_AXIMM_20_RUSER_WIDTH),
        .M_AXIMM_21_RUSER_WIDTH(M_AXIMM_21_RUSER_WIDTH),
        .M_AXIMM_22_RUSER_WIDTH(M_AXIMM_22_RUSER_WIDTH),
        .M_AXIMM_23_RUSER_WIDTH(M_AXIMM_23_RUSER_WIDTH),
        .M_AXIMM_24_RUSER_WIDTH(M_AXIMM_24_RUSER_WIDTH),
        .M_AXIMM_25_RUSER_WIDTH(M_AXIMM_25_RUSER_WIDTH),
        .M_AXIMM_26_RUSER_WIDTH(M_AXIMM_26_RUSER_WIDTH),
        .M_AXIMM_27_RUSER_WIDTH(M_AXIMM_27_RUSER_WIDTH),
        .M_AXIMM_28_RUSER_WIDTH(M_AXIMM_28_RUSER_WIDTH),
        .M_AXIMM_29_RUSER_WIDTH(M_AXIMM_29_RUSER_WIDTH),
        .M_AXIMM_30_RUSER_WIDTH(M_AXIMM_30_RUSER_WIDTH),
        .M_AXIMM_31_RUSER_WIDTH(M_AXIMM_31_RUSER_WIDTH),
        .M_AXIMM_32_RUSER_WIDTH(M_AXIMM_32_RUSER_WIDTH),
        .M_AXIMM_33_RUSER_WIDTH(M_AXIMM_33_RUSER_WIDTH),
        .M_AXIMM_34_RUSER_WIDTH(M_AXIMM_34_RUSER_WIDTH),
        .M_AXIMM_35_RUSER_WIDTH(M_AXIMM_35_RUSER_WIDTH),
        .M_AXIMM_36_RUSER_WIDTH(M_AXIMM_36_RUSER_WIDTH),
        .M_AXIMM_37_RUSER_WIDTH(M_AXIMM_37_RUSER_WIDTH),
        .M_AXIMM_38_RUSER_WIDTH(M_AXIMM_38_RUSER_WIDTH),
        .M_AXIMM_39_RUSER_WIDTH(M_AXIMM_39_RUSER_WIDTH),
        .M_AXIMM_40_RUSER_WIDTH(M_AXIMM_40_RUSER_WIDTH),
        .M_AXIMM_41_RUSER_WIDTH(M_AXIMM_41_RUSER_WIDTH),
        .M_AXIMM_42_RUSER_WIDTH(M_AXIMM_42_RUSER_WIDTH),
        .M_AXIMM_43_RUSER_WIDTH(M_AXIMM_43_RUSER_WIDTH),
        .M_AXIMM_44_RUSER_WIDTH(M_AXIMM_44_RUSER_WIDTH),
        .M_AXIMM_45_RUSER_WIDTH(M_AXIMM_45_RUSER_WIDTH),
        .M_AXIMM_46_RUSER_WIDTH(M_AXIMM_46_RUSER_WIDTH),
        .M_AXIMM_47_RUSER_WIDTH(M_AXIMM_47_RUSER_WIDTH),
        .M_AXIMM_48_RUSER_WIDTH(M_AXIMM_48_RUSER_WIDTH),
        .M_AXIMM_49_RUSER_WIDTH(M_AXIMM_49_RUSER_WIDTH),
        .M_AXIMM_50_RUSER_WIDTH(M_AXIMM_50_RUSER_WIDTH),
        .M_AXIMM_51_RUSER_WIDTH(M_AXIMM_51_RUSER_WIDTH),
        .M_AXIMM_52_RUSER_WIDTH(M_AXIMM_52_RUSER_WIDTH),
        .M_AXIMM_53_RUSER_WIDTH(M_AXIMM_53_RUSER_WIDTH),
        .M_AXIMM_54_RUSER_WIDTH(M_AXIMM_54_RUSER_WIDTH),
        .M_AXIMM_55_RUSER_WIDTH(M_AXIMM_55_RUSER_WIDTH),
        .M_AXIMM_56_RUSER_WIDTH(M_AXIMM_56_RUSER_WIDTH),
        .M_AXIMM_57_RUSER_WIDTH(M_AXIMM_57_RUSER_WIDTH),
        .M_AXIMM_58_RUSER_WIDTH(M_AXIMM_58_RUSER_WIDTH),
        .M_AXIMM_59_RUSER_WIDTH(M_AXIMM_59_RUSER_WIDTH),
        .M_AXIMM_60_RUSER_WIDTH(M_AXIMM_60_RUSER_WIDTH),
        .M_AXIMM_61_RUSER_WIDTH(M_AXIMM_61_RUSER_WIDTH),
        .M_AXIMM_62_RUSER_WIDTH(M_AXIMM_62_RUSER_WIDTH),
        .M_AXIMM_63_RUSER_WIDTH(M_AXIMM_63_RUSER_WIDTH),
        .M_AXIMM_64_RUSER_WIDTH(M_AXIMM_64_RUSER_WIDTH),
        .M_AXIMM_65_RUSER_WIDTH(M_AXIMM_65_RUSER_WIDTH),
        .M_AXIMM_66_RUSER_WIDTH(M_AXIMM_66_RUSER_WIDTH),
        .M_AXIMM_67_RUSER_WIDTH(M_AXIMM_67_RUSER_WIDTH),
        .M_AXIMM_68_RUSER_WIDTH(M_AXIMM_68_RUSER_WIDTH),
        .M_AXIMM_69_RUSER_WIDTH(M_AXIMM_69_RUSER_WIDTH),
        .M_AXIMM_70_RUSER_WIDTH(M_AXIMM_70_RUSER_WIDTH),
        .M_AXIMM_71_RUSER_WIDTH(M_AXIMM_71_RUSER_WIDTH),
        .M_AXIMM_72_RUSER_WIDTH(M_AXIMM_72_RUSER_WIDTH),
        .M_AXIMM_73_RUSER_WIDTH(M_AXIMM_73_RUSER_WIDTH),
        .M_AXIMM_74_RUSER_WIDTH(M_AXIMM_74_RUSER_WIDTH),
        .M_AXIMM_75_RUSER_WIDTH(M_AXIMM_75_RUSER_WIDTH),
        .M_AXIMM_76_RUSER_WIDTH(M_AXIMM_76_RUSER_WIDTH),
        .M_AXIMM_77_RUSER_WIDTH(M_AXIMM_77_RUSER_WIDTH),
        .M_AXIMM_78_RUSER_WIDTH(M_AXIMM_78_RUSER_WIDTH),
        .M_AXIMM_79_RUSER_WIDTH(M_AXIMM_79_RUSER_WIDTH),
        .M_AXIMM_80_RUSER_WIDTH(M_AXIMM_80_RUSER_WIDTH),
        .M_AXIMM_81_RUSER_WIDTH(M_AXIMM_81_RUSER_WIDTH),
        .M_AXIMM_82_RUSER_WIDTH(M_AXIMM_82_RUSER_WIDTH),
        .M_AXIMM_83_RUSER_WIDTH(M_AXIMM_83_RUSER_WIDTH),
        .M_AXIMM_84_RUSER_WIDTH(M_AXIMM_84_RUSER_WIDTH),
        .M_AXIMM_85_RUSER_WIDTH(M_AXIMM_85_RUSER_WIDTH),
        .M_AXIMM_86_RUSER_WIDTH(M_AXIMM_86_RUSER_WIDTH),
        .M_AXIMM_87_RUSER_WIDTH(M_AXIMM_87_RUSER_WIDTH),
        .M_AXIMM_88_RUSER_WIDTH(M_AXIMM_88_RUSER_WIDTH),
        .M_AXIMM_89_RUSER_WIDTH(M_AXIMM_89_RUSER_WIDTH),
        .M_AXIMM_90_RUSER_WIDTH(M_AXIMM_90_RUSER_WIDTH),
        .M_AXIMM_91_RUSER_WIDTH(M_AXIMM_91_RUSER_WIDTH),
        .M_AXIMM_92_RUSER_WIDTH(M_AXIMM_92_RUSER_WIDTH),
        .M_AXIMM_93_RUSER_WIDTH(M_AXIMM_93_RUSER_WIDTH),
        .M_AXIMM_94_RUSER_WIDTH(M_AXIMM_94_RUSER_WIDTH),
        .M_AXIMM_95_RUSER_WIDTH(M_AXIMM_95_RUSER_WIDTH),
        .M_AXIMM_96_RUSER_WIDTH(M_AXIMM_96_RUSER_WIDTH),
        .M_AXIMM_97_RUSER_WIDTH(M_AXIMM_97_RUSER_WIDTH),
        .M_AXIMM_98_RUSER_WIDTH(M_AXIMM_98_RUSER_WIDTH),
        .M_AXIMM_99_RUSER_WIDTH(M_AXIMM_99_RUSER_WIDTH),
        .M_AXIMM_100_RUSER_WIDTH(M_AXIMM_100_RUSER_WIDTH),
        .M_AXIMM_101_RUSER_WIDTH(M_AXIMM_101_RUSER_WIDTH),
        .M_AXIMM_102_RUSER_WIDTH(M_AXIMM_102_RUSER_WIDTH),
        .M_AXIMM_103_RUSER_WIDTH(M_AXIMM_103_RUSER_WIDTH),
        .M_AXIMM_104_RUSER_WIDTH(M_AXIMM_104_RUSER_WIDTH),
        .M_AXIMM_105_RUSER_WIDTH(M_AXIMM_105_RUSER_WIDTH),
        .M_AXIMM_106_RUSER_WIDTH(M_AXIMM_106_RUSER_WIDTH),
        .M_AXIMM_107_RUSER_WIDTH(M_AXIMM_107_RUSER_WIDTH),
        .M_AXIMM_108_RUSER_WIDTH(M_AXIMM_108_RUSER_WIDTH),
        .M_AXIMM_109_RUSER_WIDTH(M_AXIMM_109_RUSER_WIDTH),
        .M_AXIMM_110_RUSER_WIDTH(M_AXIMM_110_RUSER_WIDTH),
        .M_AXIMM_111_RUSER_WIDTH(M_AXIMM_111_RUSER_WIDTH),
        .M_AXIMM_112_RUSER_WIDTH(M_AXIMM_112_RUSER_WIDTH),
        .M_AXIMM_113_RUSER_WIDTH(M_AXIMM_113_RUSER_WIDTH),
        .M_AXIMM_114_RUSER_WIDTH(M_AXIMM_114_RUSER_WIDTH),
        .M_AXIMM_115_RUSER_WIDTH(M_AXIMM_115_RUSER_WIDTH),
        .M_AXIMM_116_RUSER_WIDTH(M_AXIMM_116_RUSER_WIDTH),
        .M_AXIMM_117_RUSER_WIDTH(M_AXIMM_117_RUSER_WIDTH),
        .M_AXIMM_118_RUSER_WIDTH(M_AXIMM_118_RUSER_WIDTH),
        .M_AXIMM_119_RUSER_WIDTH(M_AXIMM_119_RUSER_WIDTH),
        .M_AXIMM_120_RUSER_WIDTH(M_AXIMM_120_RUSER_WIDTH),
        .M_AXIMM_121_RUSER_WIDTH(M_AXIMM_121_RUSER_WIDTH),
        .M_AXIMM_122_RUSER_WIDTH(M_AXIMM_122_RUSER_WIDTH),
        .M_AXIMM_123_RUSER_WIDTH(M_AXIMM_123_RUSER_WIDTH),
        .M_AXIMM_124_RUSER_WIDTH(M_AXIMM_124_RUSER_WIDTH),
        .M_AXIMM_125_RUSER_WIDTH(M_AXIMM_125_RUSER_WIDTH),
        .M_AXIMM_126_RUSER_WIDTH(M_AXIMM_126_RUSER_WIDTH),
        .M_AXIMM_127_RUSER_WIDTH(M_AXIMM_127_RUSER_WIDTH),
        .M_AXIMM_0_ARID_WIDTH(M_AXIMM_0_ARID_WIDTH),
        .M_AXIMM_1_ARID_WIDTH(M_AXIMM_1_ARID_WIDTH),
        .M_AXIMM_2_ARID_WIDTH(M_AXIMM_2_ARID_WIDTH),
        .M_AXIMM_3_ARID_WIDTH(M_AXIMM_3_ARID_WIDTH),
        .M_AXIMM_4_ARID_WIDTH(M_AXIMM_4_ARID_WIDTH),
        .M_AXIMM_5_ARID_WIDTH(M_AXIMM_5_ARID_WIDTH),
        .M_AXIMM_6_ARID_WIDTH(M_AXIMM_6_ARID_WIDTH),
        .M_AXIMM_7_ARID_WIDTH(M_AXIMM_7_ARID_WIDTH),
        .M_AXIMM_8_ARID_WIDTH(M_AXIMM_8_ARID_WIDTH),
        .M_AXIMM_9_ARID_WIDTH(M_AXIMM_9_ARID_WIDTH),
        .M_AXIMM_10_ARID_WIDTH(M_AXIMM_10_ARID_WIDTH),
        .M_AXIMM_11_ARID_WIDTH(M_AXIMM_11_ARID_WIDTH),
        .M_AXIMM_12_ARID_WIDTH(M_AXIMM_12_ARID_WIDTH),
        .M_AXIMM_13_ARID_WIDTH(M_AXIMM_13_ARID_WIDTH),
        .M_AXIMM_14_ARID_WIDTH(M_AXIMM_14_ARID_WIDTH),
        .M_AXIMM_15_ARID_WIDTH(M_AXIMM_15_ARID_WIDTH),
        .M_AXIMM_16_ARID_WIDTH(M_AXIMM_16_ARID_WIDTH),
        .M_AXIMM_17_ARID_WIDTH(M_AXIMM_17_ARID_WIDTH),
        .M_AXIMM_18_ARID_WIDTH(M_AXIMM_18_ARID_WIDTH),
        .M_AXIMM_19_ARID_WIDTH(M_AXIMM_19_ARID_WIDTH),
        .M_AXIMM_20_ARID_WIDTH(M_AXIMM_20_ARID_WIDTH),
        .M_AXIMM_21_ARID_WIDTH(M_AXIMM_21_ARID_WIDTH),
        .M_AXIMM_22_ARID_WIDTH(M_AXIMM_22_ARID_WIDTH),
        .M_AXIMM_23_ARID_WIDTH(M_AXIMM_23_ARID_WIDTH),
        .M_AXIMM_24_ARID_WIDTH(M_AXIMM_24_ARID_WIDTH),
        .M_AXIMM_25_ARID_WIDTH(M_AXIMM_25_ARID_WIDTH),
        .M_AXIMM_26_ARID_WIDTH(M_AXIMM_26_ARID_WIDTH),
        .M_AXIMM_27_ARID_WIDTH(M_AXIMM_27_ARID_WIDTH),
        .M_AXIMM_28_ARID_WIDTH(M_AXIMM_28_ARID_WIDTH),
        .M_AXIMM_29_ARID_WIDTH(M_AXIMM_29_ARID_WIDTH),
        .M_AXIMM_30_ARID_WIDTH(M_AXIMM_30_ARID_WIDTH),
        .M_AXIMM_31_ARID_WIDTH(M_AXIMM_31_ARID_WIDTH),
        .M_AXIMM_32_ARID_WIDTH(M_AXIMM_32_ARID_WIDTH),
        .M_AXIMM_33_ARID_WIDTH(M_AXIMM_33_ARID_WIDTH),
        .M_AXIMM_34_ARID_WIDTH(M_AXIMM_34_ARID_WIDTH),
        .M_AXIMM_35_ARID_WIDTH(M_AXIMM_35_ARID_WIDTH),
        .M_AXIMM_36_ARID_WIDTH(M_AXIMM_36_ARID_WIDTH),
        .M_AXIMM_37_ARID_WIDTH(M_AXIMM_37_ARID_WIDTH),
        .M_AXIMM_38_ARID_WIDTH(M_AXIMM_38_ARID_WIDTH),
        .M_AXIMM_39_ARID_WIDTH(M_AXIMM_39_ARID_WIDTH),
        .M_AXIMM_40_ARID_WIDTH(M_AXIMM_40_ARID_WIDTH),
        .M_AXIMM_41_ARID_WIDTH(M_AXIMM_41_ARID_WIDTH),
        .M_AXIMM_42_ARID_WIDTH(M_AXIMM_42_ARID_WIDTH),
        .M_AXIMM_43_ARID_WIDTH(M_AXIMM_43_ARID_WIDTH),
        .M_AXIMM_44_ARID_WIDTH(M_AXIMM_44_ARID_WIDTH),
        .M_AXIMM_45_ARID_WIDTH(M_AXIMM_45_ARID_WIDTH),
        .M_AXIMM_46_ARID_WIDTH(M_AXIMM_46_ARID_WIDTH),
        .M_AXIMM_47_ARID_WIDTH(M_AXIMM_47_ARID_WIDTH),
        .M_AXIMM_48_ARID_WIDTH(M_AXIMM_48_ARID_WIDTH),
        .M_AXIMM_49_ARID_WIDTH(M_AXIMM_49_ARID_WIDTH),
        .M_AXIMM_50_ARID_WIDTH(M_AXIMM_50_ARID_WIDTH),
        .M_AXIMM_51_ARID_WIDTH(M_AXIMM_51_ARID_WIDTH),
        .M_AXIMM_52_ARID_WIDTH(M_AXIMM_52_ARID_WIDTH),
        .M_AXIMM_53_ARID_WIDTH(M_AXIMM_53_ARID_WIDTH),
        .M_AXIMM_54_ARID_WIDTH(M_AXIMM_54_ARID_WIDTH),
        .M_AXIMM_55_ARID_WIDTH(M_AXIMM_55_ARID_WIDTH),
        .M_AXIMM_56_ARID_WIDTH(M_AXIMM_56_ARID_WIDTH),
        .M_AXIMM_57_ARID_WIDTH(M_AXIMM_57_ARID_WIDTH),
        .M_AXIMM_58_ARID_WIDTH(M_AXIMM_58_ARID_WIDTH),
        .M_AXIMM_59_ARID_WIDTH(M_AXIMM_59_ARID_WIDTH),
        .M_AXIMM_60_ARID_WIDTH(M_AXIMM_60_ARID_WIDTH),
        .M_AXIMM_61_ARID_WIDTH(M_AXIMM_61_ARID_WIDTH),
        .M_AXIMM_62_ARID_WIDTH(M_AXIMM_62_ARID_WIDTH),
        .M_AXIMM_63_ARID_WIDTH(M_AXIMM_63_ARID_WIDTH),
        .M_AXIMM_64_ARID_WIDTH(M_AXIMM_64_ARID_WIDTH),
        .M_AXIMM_65_ARID_WIDTH(M_AXIMM_65_ARID_WIDTH),
        .M_AXIMM_66_ARID_WIDTH(M_AXIMM_66_ARID_WIDTH),
        .M_AXIMM_67_ARID_WIDTH(M_AXIMM_67_ARID_WIDTH),
        .M_AXIMM_68_ARID_WIDTH(M_AXIMM_68_ARID_WIDTH),
        .M_AXIMM_69_ARID_WIDTH(M_AXIMM_69_ARID_WIDTH),
        .M_AXIMM_70_ARID_WIDTH(M_AXIMM_70_ARID_WIDTH),
        .M_AXIMM_71_ARID_WIDTH(M_AXIMM_71_ARID_WIDTH),
        .M_AXIMM_72_ARID_WIDTH(M_AXIMM_72_ARID_WIDTH),
        .M_AXIMM_73_ARID_WIDTH(M_AXIMM_73_ARID_WIDTH),
        .M_AXIMM_74_ARID_WIDTH(M_AXIMM_74_ARID_WIDTH),
        .M_AXIMM_75_ARID_WIDTH(M_AXIMM_75_ARID_WIDTH),
        .M_AXIMM_76_ARID_WIDTH(M_AXIMM_76_ARID_WIDTH),
        .M_AXIMM_77_ARID_WIDTH(M_AXIMM_77_ARID_WIDTH),
        .M_AXIMM_78_ARID_WIDTH(M_AXIMM_78_ARID_WIDTH),
        .M_AXIMM_79_ARID_WIDTH(M_AXIMM_79_ARID_WIDTH),
        .M_AXIMM_80_ARID_WIDTH(M_AXIMM_80_ARID_WIDTH),
        .M_AXIMM_81_ARID_WIDTH(M_AXIMM_81_ARID_WIDTH),
        .M_AXIMM_82_ARID_WIDTH(M_AXIMM_82_ARID_WIDTH),
        .M_AXIMM_83_ARID_WIDTH(M_AXIMM_83_ARID_WIDTH),
        .M_AXIMM_84_ARID_WIDTH(M_AXIMM_84_ARID_WIDTH),
        .M_AXIMM_85_ARID_WIDTH(M_AXIMM_85_ARID_WIDTH),
        .M_AXIMM_86_ARID_WIDTH(M_AXIMM_86_ARID_WIDTH),
        .M_AXIMM_87_ARID_WIDTH(M_AXIMM_87_ARID_WIDTH),
        .M_AXIMM_88_ARID_WIDTH(M_AXIMM_88_ARID_WIDTH),
        .M_AXIMM_89_ARID_WIDTH(M_AXIMM_89_ARID_WIDTH),
        .M_AXIMM_90_ARID_WIDTH(M_AXIMM_90_ARID_WIDTH),
        .M_AXIMM_91_ARID_WIDTH(M_AXIMM_91_ARID_WIDTH),
        .M_AXIMM_92_ARID_WIDTH(M_AXIMM_92_ARID_WIDTH),
        .M_AXIMM_93_ARID_WIDTH(M_AXIMM_93_ARID_WIDTH),
        .M_AXIMM_94_ARID_WIDTH(M_AXIMM_94_ARID_WIDTH),
        .M_AXIMM_95_ARID_WIDTH(M_AXIMM_95_ARID_WIDTH),
        .M_AXIMM_96_ARID_WIDTH(M_AXIMM_96_ARID_WIDTH),
        .M_AXIMM_97_ARID_WIDTH(M_AXIMM_97_ARID_WIDTH),
        .M_AXIMM_98_ARID_WIDTH(M_AXIMM_98_ARID_WIDTH),
        .M_AXIMM_99_ARID_WIDTH(M_AXIMM_99_ARID_WIDTH),
        .M_AXIMM_100_ARID_WIDTH(M_AXIMM_100_ARID_WIDTH),
        .M_AXIMM_101_ARID_WIDTH(M_AXIMM_101_ARID_WIDTH),
        .M_AXIMM_102_ARID_WIDTH(M_AXIMM_102_ARID_WIDTH),
        .M_AXIMM_103_ARID_WIDTH(M_AXIMM_103_ARID_WIDTH),
        .M_AXIMM_104_ARID_WIDTH(M_AXIMM_104_ARID_WIDTH),
        .M_AXIMM_105_ARID_WIDTH(M_AXIMM_105_ARID_WIDTH),
        .M_AXIMM_106_ARID_WIDTH(M_AXIMM_106_ARID_WIDTH),
        .M_AXIMM_107_ARID_WIDTH(M_AXIMM_107_ARID_WIDTH),
        .M_AXIMM_108_ARID_WIDTH(M_AXIMM_108_ARID_WIDTH),
        .M_AXIMM_109_ARID_WIDTH(M_AXIMM_109_ARID_WIDTH),
        .M_AXIMM_110_ARID_WIDTH(M_AXIMM_110_ARID_WIDTH),
        .M_AXIMM_111_ARID_WIDTH(M_AXIMM_111_ARID_WIDTH),
        .M_AXIMM_112_ARID_WIDTH(M_AXIMM_112_ARID_WIDTH),
        .M_AXIMM_113_ARID_WIDTH(M_AXIMM_113_ARID_WIDTH),
        .M_AXIMM_114_ARID_WIDTH(M_AXIMM_114_ARID_WIDTH),
        .M_AXIMM_115_ARID_WIDTH(M_AXIMM_115_ARID_WIDTH),
        .M_AXIMM_116_ARID_WIDTH(M_AXIMM_116_ARID_WIDTH),
        .M_AXIMM_117_ARID_WIDTH(M_AXIMM_117_ARID_WIDTH),
        .M_AXIMM_118_ARID_WIDTH(M_AXIMM_118_ARID_WIDTH),
        .M_AXIMM_119_ARID_WIDTH(M_AXIMM_119_ARID_WIDTH),
        .M_AXIMM_120_ARID_WIDTH(M_AXIMM_120_ARID_WIDTH),
        .M_AXIMM_121_ARID_WIDTH(M_AXIMM_121_ARID_WIDTH),
        .M_AXIMM_122_ARID_WIDTH(M_AXIMM_122_ARID_WIDTH),
        .M_AXIMM_123_ARID_WIDTH(M_AXIMM_123_ARID_WIDTH),
        .M_AXIMM_124_ARID_WIDTH(M_AXIMM_124_ARID_WIDTH),
        .M_AXIMM_125_ARID_WIDTH(M_AXIMM_125_ARID_WIDTH),
        .M_AXIMM_126_ARID_WIDTH(M_AXIMM_126_ARID_WIDTH),
        .M_AXIMM_127_ARID_WIDTH(M_AXIMM_127_ARID_WIDTH),
        .M_AXIMM_0_AWID_WIDTH(M_AXIMM_0_AWID_WIDTH),
        .M_AXIMM_1_AWID_WIDTH(M_AXIMM_1_AWID_WIDTH),
        .M_AXIMM_2_AWID_WIDTH(M_AXIMM_2_AWID_WIDTH),
        .M_AXIMM_3_AWID_WIDTH(M_AXIMM_3_AWID_WIDTH),
        .M_AXIMM_4_AWID_WIDTH(M_AXIMM_4_AWID_WIDTH),
        .M_AXIMM_5_AWID_WIDTH(M_AXIMM_5_AWID_WIDTH),
        .M_AXIMM_6_AWID_WIDTH(M_AXIMM_6_AWID_WIDTH),
        .M_AXIMM_7_AWID_WIDTH(M_AXIMM_7_AWID_WIDTH),
        .M_AXIMM_8_AWID_WIDTH(M_AXIMM_8_AWID_WIDTH),
        .M_AXIMM_9_AWID_WIDTH(M_AXIMM_9_AWID_WIDTH),
        .M_AXIMM_10_AWID_WIDTH(M_AXIMM_10_AWID_WIDTH),
        .M_AXIMM_11_AWID_WIDTH(M_AXIMM_11_AWID_WIDTH),
        .M_AXIMM_12_AWID_WIDTH(M_AXIMM_12_AWID_WIDTH),
        .M_AXIMM_13_AWID_WIDTH(M_AXIMM_13_AWID_WIDTH),
        .M_AXIMM_14_AWID_WIDTH(M_AXIMM_14_AWID_WIDTH),
        .M_AXIMM_15_AWID_WIDTH(M_AXIMM_15_AWID_WIDTH),
        .M_AXIMM_16_AWID_WIDTH(M_AXIMM_16_AWID_WIDTH),
        .M_AXIMM_17_AWID_WIDTH(M_AXIMM_17_AWID_WIDTH),
        .M_AXIMM_18_AWID_WIDTH(M_AXIMM_18_AWID_WIDTH),
        .M_AXIMM_19_AWID_WIDTH(M_AXIMM_19_AWID_WIDTH),
        .M_AXIMM_20_AWID_WIDTH(M_AXIMM_20_AWID_WIDTH),
        .M_AXIMM_21_AWID_WIDTH(M_AXIMM_21_AWID_WIDTH),
        .M_AXIMM_22_AWID_WIDTH(M_AXIMM_22_AWID_WIDTH),
        .M_AXIMM_23_AWID_WIDTH(M_AXIMM_23_AWID_WIDTH),
        .M_AXIMM_24_AWID_WIDTH(M_AXIMM_24_AWID_WIDTH),
        .M_AXIMM_25_AWID_WIDTH(M_AXIMM_25_AWID_WIDTH),
        .M_AXIMM_26_AWID_WIDTH(M_AXIMM_26_AWID_WIDTH),
        .M_AXIMM_27_AWID_WIDTH(M_AXIMM_27_AWID_WIDTH),
        .M_AXIMM_28_AWID_WIDTH(M_AXIMM_28_AWID_WIDTH),
        .M_AXIMM_29_AWID_WIDTH(M_AXIMM_29_AWID_WIDTH),
        .M_AXIMM_30_AWID_WIDTH(M_AXIMM_30_AWID_WIDTH),
        .M_AXIMM_31_AWID_WIDTH(M_AXIMM_31_AWID_WIDTH),
        .M_AXIMM_32_AWID_WIDTH(M_AXIMM_32_AWID_WIDTH),
        .M_AXIMM_33_AWID_WIDTH(M_AXIMM_33_AWID_WIDTH),
        .M_AXIMM_34_AWID_WIDTH(M_AXIMM_34_AWID_WIDTH),
        .M_AXIMM_35_AWID_WIDTH(M_AXIMM_35_AWID_WIDTH),
        .M_AXIMM_36_AWID_WIDTH(M_AXIMM_36_AWID_WIDTH),
        .M_AXIMM_37_AWID_WIDTH(M_AXIMM_37_AWID_WIDTH),
        .M_AXIMM_38_AWID_WIDTH(M_AXIMM_38_AWID_WIDTH),
        .M_AXIMM_39_AWID_WIDTH(M_AXIMM_39_AWID_WIDTH),
        .M_AXIMM_40_AWID_WIDTH(M_AXIMM_40_AWID_WIDTH),
        .M_AXIMM_41_AWID_WIDTH(M_AXIMM_41_AWID_WIDTH),
        .M_AXIMM_42_AWID_WIDTH(M_AXIMM_42_AWID_WIDTH),
        .M_AXIMM_43_AWID_WIDTH(M_AXIMM_43_AWID_WIDTH),
        .M_AXIMM_44_AWID_WIDTH(M_AXIMM_44_AWID_WIDTH),
        .M_AXIMM_45_AWID_WIDTH(M_AXIMM_45_AWID_WIDTH),
        .M_AXIMM_46_AWID_WIDTH(M_AXIMM_46_AWID_WIDTH),
        .M_AXIMM_47_AWID_WIDTH(M_AXIMM_47_AWID_WIDTH),
        .M_AXIMM_48_AWID_WIDTH(M_AXIMM_48_AWID_WIDTH),
        .M_AXIMM_49_AWID_WIDTH(M_AXIMM_49_AWID_WIDTH),
        .M_AXIMM_50_AWID_WIDTH(M_AXIMM_50_AWID_WIDTH),
        .M_AXIMM_51_AWID_WIDTH(M_AXIMM_51_AWID_WIDTH),
        .M_AXIMM_52_AWID_WIDTH(M_AXIMM_52_AWID_WIDTH),
        .M_AXIMM_53_AWID_WIDTH(M_AXIMM_53_AWID_WIDTH),
        .M_AXIMM_54_AWID_WIDTH(M_AXIMM_54_AWID_WIDTH),
        .M_AXIMM_55_AWID_WIDTH(M_AXIMM_55_AWID_WIDTH),
        .M_AXIMM_56_AWID_WIDTH(M_AXIMM_56_AWID_WIDTH),
        .M_AXIMM_57_AWID_WIDTH(M_AXIMM_57_AWID_WIDTH),
        .M_AXIMM_58_AWID_WIDTH(M_AXIMM_58_AWID_WIDTH),
        .M_AXIMM_59_AWID_WIDTH(M_AXIMM_59_AWID_WIDTH),
        .M_AXIMM_60_AWID_WIDTH(M_AXIMM_60_AWID_WIDTH),
        .M_AXIMM_61_AWID_WIDTH(M_AXIMM_61_AWID_WIDTH),
        .M_AXIMM_62_AWID_WIDTH(M_AXIMM_62_AWID_WIDTH),
        .M_AXIMM_63_AWID_WIDTH(M_AXIMM_63_AWID_WIDTH),
        .M_AXIMM_64_AWID_WIDTH(M_AXIMM_64_AWID_WIDTH),
        .M_AXIMM_65_AWID_WIDTH(M_AXIMM_65_AWID_WIDTH),
        .M_AXIMM_66_AWID_WIDTH(M_AXIMM_66_AWID_WIDTH),
        .M_AXIMM_67_AWID_WIDTH(M_AXIMM_67_AWID_WIDTH),
        .M_AXIMM_68_AWID_WIDTH(M_AXIMM_68_AWID_WIDTH),
        .M_AXIMM_69_AWID_WIDTH(M_AXIMM_69_AWID_WIDTH),
        .M_AXIMM_70_AWID_WIDTH(M_AXIMM_70_AWID_WIDTH),
        .M_AXIMM_71_AWID_WIDTH(M_AXIMM_71_AWID_WIDTH),
        .M_AXIMM_72_AWID_WIDTH(M_AXIMM_72_AWID_WIDTH),
        .M_AXIMM_73_AWID_WIDTH(M_AXIMM_73_AWID_WIDTH),
        .M_AXIMM_74_AWID_WIDTH(M_AXIMM_74_AWID_WIDTH),
        .M_AXIMM_75_AWID_WIDTH(M_AXIMM_75_AWID_WIDTH),
        .M_AXIMM_76_AWID_WIDTH(M_AXIMM_76_AWID_WIDTH),
        .M_AXIMM_77_AWID_WIDTH(M_AXIMM_77_AWID_WIDTH),
        .M_AXIMM_78_AWID_WIDTH(M_AXIMM_78_AWID_WIDTH),
        .M_AXIMM_79_AWID_WIDTH(M_AXIMM_79_AWID_WIDTH),
        .M_AXIMM_80_AWID_WIDTH(M_AXIMM_80_AWID_WIDTH),
        .M_AXIMM_81_AWID_WIDTH(M_AXIMM_81_AWID_WIDTH),
        .M_AXIMM_82_AWID_WIDTH(M_AXIMM_82_AWID_WIDTH),
        .M_AXIMM_83_AWID_WIDTH(M_AXIMM_83_AWID_WIDTH),
        .M_AXIMM_84_AWID_WIDTH(M_AXIMM_84_AWID_WIDTH),
        .M_AXIMM_85_AWID_WIDTH(M_AXIMM_85_AWID_WIDTH),
        .M_AXIMM_86_AWID_WIDTH(M_AXIMM_86_AWID_WIDTH),
        .M_AXIMM_87_AWID_WIDTH(M_AXIMM_87_AWID_WIDTH),
        .M_AXIMM_88_AWID_WIDTH(M_AXIMM_88_AWID_WIDTH),
        .M_AXIMM_89_AWID_WIDTH(M_AXIMM_89_AWID_WIDTH),
        .M_AXIMM_90_AWID_WIDTH(M_AXIMM_90_AWID_WIDTH),
        .M_AXIMM_91_AWID_WIDTH(M_AXIMM_91_AWID_WIDTH),
        .M_AXIMM_92_AWID_WIDTH(M_AXIMM_92_AWID_WIDTH),
        .M_AXIMM_93_AWID_WIDTH(M_AXIMM_93_AWID_WIDTH),
        .M_AXIMM_94_AWID_WIDTH(M_AXIMM_94_AWID_WIDTH),
        .M_AXIMM_95_AWID_WIDTH(M_AXIMM_95_AWID_WIDTH),
        .M_AXIMM_96_AWID_WIDTH(M_AXIMM_96_AWID_WIDTH),
        .M_AXIMM_97_AWID_WIDTH(M_AXIMM_97_AWID_WIDTH),
        .M_AXIMM_98_AWID_WIDTH(M_AXIMM_98_AWID_WIDTH),
        .M_AXIMM_99_AWID_WIDTH(M_AXIMM_99_AWID_WIDTH),
        .M_AXIMM_100_AWID_WIDTH(M_AXIMM_100_AWID_WIDTH),
        .M_AXIMM_101_AWID_WIDTH(M_AXIMM_101_AWID_WIDTH),
        .M_AXIMM_102_AWID_WIDTH(M_AXIMM_102_AWID_WIDTH),
        .M_AXIMM_103_AWID_WIDTH(M_AXIMM_103_AWID_WIDTH),
        .M_AXIMM_104_AWID_WIDTH(M_AXIMM_104_AWID_WIDTH),
        .M_AXIMM_105_AWID_WIDTH(M_AXIMM_105_AWID_WIDTH),
        .M_AXIMM_106_AWID_WIDTH(M_AXIMM_106_AWID_WIDTH),
        .M_AXIMM_107_AWID_WIDTH(M_AXIMM_107_AWID_WIDTH),
        .M_AXIMM_108_AWID_WIDTH(M_AXIMM_108_AWID_WIDTH),
        .M_AXIMM_109_AWID_WIDTH(M_AXIMM_109_AWID_WIDTH),
        .M_AXIMM_110_AWID_WIDTH(M_AXIMM_110_AWID_WIDTH),
        .M_AXIMM_111_AWID_WIDTH(M_AXIMM_111_AWID_WIDTH),
        .M_AXIMM_112_AWID_WIDTH(M_AXIMM_112_AWID_WIDTH),
        .M_AXIMM_113_AWID_WIDTH(M_AXIMM_113_AWID_WIDTH),
        .M_AXIMM_114_AWID_WIDTH(M_AXIMM_114_AWID_WIDTH),
        .M_AXIMM_115_AWID_WIDTH(M_AXIMM_115_AWID_WIDTH),
        .M_AXIMM_116_AWID_WIDTH(M_AXIMM_116_AWID_WIDTH),
        .M_AXIMM_117_AWID_WIDTH(M_AXIMM_117_AWID_WIDTH),
        .M_AXIMM_118_AWID_WIDTH(M_AXIMM_118_AWID_WIDTH),
        .M_AXIMM_119_AWID_WIDTH(M_AXIMM_119_AWID_WIDTH),
        .M_AXIMM_120_AWID_WIDTH(M_AXIMM_120_AWID_WIDTH),
        .M_AXIMM_121_AWID_WIDTH(M_AXIMM_121_AWID_WIDTH),
        .M_AXIMM_122_AWID_WIDTH(M_AXIMM_122_AWID_WIDTH),
        .M_AXIMM_123_AWID_WIDTH(M_AXIMM_123_AWID_WIDTH),
        .M_AXIMM_124_AWID_WIDTH(M_AXIMM_124_AWID_WIDTH),
        .M_AXIMM_125_AWID_WIDTH(M_AXIMM_125_AWID_WIDTH),
        .M_AXIMM_126_AWID_WIDTH(M_AXIMM_126_AWID_WIDTH),
        .M_AXIMM_127_AWID_WIDTH(M_AXIMM_127_AWID_WIDTH),
        .M_AXIMM_0_WID_WIDTH(M_AXIMM_0_WID_WIDTH),
        .M_AXIMM_1_WID_WIDTH(M_AXIMM_1_WID_WIDTH),
        .M_AXIMM_2_WID_WIDTH(M_AXIMM_2_WID_WIDTH),
        .M_AXIMM_3_WID_WIDTH(M_AXIMM_3_WID_WIDTH),
        .M_AXIMM_4_WID_WIDTH(M_AXIMM_4_WID_WIDTH),
        .M_AXIMM_5_WID_WIDTH(M_AXIMM_5_WID_WIDTH),
        .M_AXIMM_6_WID_WIDTH(M_AXIMM_6_WID_WIDTH),
        .M_AXIMM_7_WID_WIDTH(M_AXIMM_7_WID_WIDTH),
        .M_AXIMM_8_WID_WIDTH(M_AXIMM_8_WID_WIDTH),
        .M_AXIMM_9_WID_WIDTH(M_AXIMM_9_WID_WIDTH),
        .M_AXIMM_10_WID_WIDTH(M_AXIMM_10_WID_WIDTH),
        .M_AXIMM_11_WID_WIDTH(M_AXIMM_11_WID_WIDTH),
        .M_AXIMM_12_WID_WIDTH(M_AXIMM_12_WID_WIDTH),
        .M_AXIMM_13_WID_WIDTH(M_AXIMM_13_WID_WIDTH),
        .M_AXIMM_14_WID_WIDTH(M_AXIMM_14_WID_WIDTH),
        .M_AXIMM_15_WID_WIDTH(M_AXIMM_15_WID_WIDTH),
        .M_AXIMM_16_WID_WIDTH(M_AXIMM_16_WID_WIDTH),
        .M_AXIMM_17_WID_WIDTH(M_AXIMM_17_WID_WIDTH),
        .M_AXIMM_18_WID_WIDTH(M_AXIMM_18_WID_WIDTH),
        .M_AXIMM_19_WID_WIDTH(M_AXIMM_19_WID_WIDTH),
        .M_AXIMM_20_WID_WIDTH(M_AXIMM_20_WID_WIDTH),
        .M_AXIMM_21_WID_WIDTH(M_AXIMM_21_WID_WIDTH),
        .M_AXIMM_22_WID_WIDTH(M_AXIMM_22_WID_WIDTH),
        .M_AXIMM_23_WID_WIDTH(M_AXIMM_23_WID_WIDTH),
        .M_AXIMM_24_WID_WIDTH(M_AXIMM_24_WID_WIDTH),
        .M_AXIMM_25_WID_WIDTH(M_AXIMM_25_WID_WIDTH),
        .M_AXIMM_26_WID_WIDTH(M_AXIMM_26_WID_WIDTH),
        .M_AXIMM_27_WID_WIDTH(M_AXIMM_27_WID_WIDTH),
        .M_AXIMM_28_WID_WIDTH(M_AXIMM_28_WID_WIDTH),
        .M_AXIMM_29_WID_WIDTH(M_AXIMM_29_WID_WIDTH),
        .M_AXIMM_30_WID_WIDTH(M_AXIMM_30_WID_WIDTH),
        .M_AXIMM_31_WID_WIDTH(M_AXIMM_31_WID_WIDTH),
        .M_AXIMM_32_WID_WIDTH(M_AXIMM_32_WID_WIDTH),
        .M_AXIMM_33_WID_WIDTH(M_AXIMM_33_WID_WIDTH),
        .M_AXIMM_34_WID_WIDTH(M_AXIMM_34_WID_WIDTH),
        .M_AXIMM_35_WID_WIDTH(M_AXIMM_35_WID_WIDTH),
        .M_AXIMM_36_WID_WIDTH(M_AXIMM_36_WID_WIDTH),
        .M_AXIMM_37_WID_WIDTH(M_AXIMM_37_WID_WIDTH),
        .M_AXIMM_38_WID_WIDTH(M_AXIMM_38_WID_WIDTH),
        .M_AXIMM_39_WID_WIDTH(M_AXIMM_39_WID_WIDTH),
        .M_AXIMM_40_WID_WIDTH(M_AXIMM_40_WID_WIDTH),
        .M_AXIMM_41_WID_WIDTH(M_AXIMM_41_WID_WIDTH),
        .M_AXIMM_42_WID_WIDTH(M_AXIMM_42_WID_WIDTH),
        .M_AXIMM_43_WID_WIDTH(M_AXIMM_43_WID_WIDTH),
        .M_AXIMM_44_WID_WIDTH(M_AXIMM_44_WID_WIDTH),
        .M_AXIMM_45_WID_WIDTH(M_AXIMM_45_WID_WIDTH),
        .M_AXIMM_46_WID_WIDTH(M_AXIMM_46_WID_WIDTH),
        .M_AXIMM_47_WID_WIDTH(M_AXIMM_47_WID_WIDTH),
        .M_AXIMM_48_WID_WIDTH(M_AXIMM_48_WID_WIDTH),
        .M_AXIMM_49_WID_WIDTH(M_AXIMM_49_WID_WIDTH),
        .M_AXIMM_50_WID_WIDTH(M_AXIMM_50_WID_WIDTH),
        .M_AXIMM_51_WID_WIDTH(M_AXIMM_51_WID_WIDTH),
        .M_AXIMM_52_WID_WIDTH(M_AXIMM_52_WID_WIDTH),
        .M_AXIMM_53_WID_WIDTH(M_AXIMM_53_WID_WIDTH),
        .M_AXIMM_54_WID_WIDTH(M_AXIMM_54_WID_WIDTH),
        .M_AXIMM_55_WID_WIDTH(M_AXIMM_55_WID_WIDTH),
        .M_AXIMM_56_WID_WIDTH(M_AXIMM_56_WID_WIDTH),
        .M_AXIMM_57_WID_WIDTH(M_AXIMM_57_WID_WIDTH),
        .M_AXIMM_58_WID_WIDTH(M_AXIMM_58_WID_WIDTH),
        .M_AXIMM_59_WID_WIDTH(M_AXIMM_59_WID_WIDTH),
        .M_AXIMM_60_WID_WIDTH(M_AXIMM_60_WID_WIDTH),
        .M_AXIMM_61_WID_WIDTH(M_AXIMM_61_WID_WIDTH),
        .M_AXIMM_62_WID_WIDTH(M_AXIMM_62_WID_WIDTH),
        .M_AXIMM_63_WID_WIDTH(M_AXIMM_63_WID_WIDTH),
        .M_AXIMM_64_WID_WIDTH(M_AXIMM_64_WID_WIDTH),
        .M_AXIMM_65_WID_WIDTH(M_AXIMM_65_WID_WIDTH),
        .M_AXIMM_66_WID_WIDTH(M_AXIMM_66_WID_WIDTH),
        .M_AXIMM_67_WID_WIDTH(M_AXIMM_67_WID_WIDTH),
        .M_AXIMM_68_WID_WIDTH(M_AXIMM_68_WID_WIDTH),
        .M_AXIMM_69_WID_WIDTH(M_AXIMM_69_WID_WIDTH),
        .M_AXIMM_70_WID_WIDTH(M_AXIMM_70_WID_WIDTH),
        .M_AXIMM_71_WID_WIDTH(M_AXIMM_71_WID_WIDTH),
        .M_AXIMM_72_WID_WIDTH(M_AXIMM_72_WID_WIDTH),
        .M_AXIMM_73_WID_WIDTH(M_AXIMM_73_WID_WIDTH),
        .M_AXIMM_74_WID_WIDTH(M_AXIMM_74_WID_WIDTH),
        .M_AXIMM_75_WID_WIDTH(M_AXIMM_75_WID_WIDTH),
        .M_AXIMM_76_WID_WIDTH(M_AXIMM_76_WID_WIDTH),
        .M_AXIMM_77_WID_WIDTH(M_AXIMM_77_WID_WIDTH),
        .M_AXIMM_78_WID_WIDTH(M_AXIMM_78_WID_WIDTH),
        .M_AXIMM_79_WID_WIDTH(M_AXIMM_79_WID_WIDTH),
        .M_AXIMM_80_WID_WIDTH(M_AXIMM_80_WID_WIDTH),
        .M_AXIMM_81_WID_WIDTH(M_AXIMM_81_WID_WIDTH),
        .M_AXIMM_82_WID_WIDTH(M_AXIMM_82_WID_WIDTH),
        .M_AXIMM_83_WID_WIDTH(M_AXIMM_83_WID_WIDTH),
        .M_AXIMM_84_WID_WIDTH(M_AXIMM_84_WID_WIDTH),
        .M_AXIMM_85_WID_WIDTH(M_AXIMM_85_WID_WIDTH),
        .M_AXIMM_86_WID_WIDTH(M_AXIMM_86_WID_WIDTH),
        .M_AXIMM_87_WID_WIDTH(M_AXIMM_87_WID_WIDTH),
        .M_AXIMM_88_WID_WIDTH(M_AXIMM_88_WID_WIDTH),
        .M_AXIMM_89_WID_WIDTH(M_AXIMM_89_WID_WIDTH),
        .M_AXIMM_90_WID_WIDTH(M_AXIMM_90_WID_WIDTH),
        .M_AXIMM_91_WID_WIDTH(M_AXIMM_91_WID_WIDTH),
        .M_AXIMM_92_WID_WIDTH(M_AXIMM_92_WID_WIDTH),
        .M_AXIMM_93_WID_WIDTH(M_AXIMM_93_WID_WIDTH),
        .M_AXIMM_94_WID_WIDTH(M_AXIMM_94_WID_WIDTH),
        .M_AXIMM_95_WID_WIDTH(M_AXIMM_95_WID_WIDTH),
        .M_AXIMM_96_WID_WIDTH(M_AXIMM_96_WID_WIDTH),
        .M_AXIMM_97_WID_WIDTH(M_AXIMM_97_WID_WIDTH),
        .M_AXIMM_98_WID_WIDTH(M_AXIMM_98_WID_WIDTH),
        .M_AXIMM_99_WID_WIDTH(M_AXIMM_99_WID_WIDTH),
        .M_AXIMM_100_WID_WIDTH(M_AXIMM_100_WID_WIDTH),
        .M_AXIMM_101_WID_WIDTH(M_AXIMM_101_WID_WIDTH),
        .M_AXIMM_102_WID_WIDTH(M_AXIMM_102_WID_WIDTH),
        .M_AXIMM_103_WID_WIDTH(M_AXIMM_103_WID_WIDTH),
        .M_AXIMM_104_WID_WIDTH(M_AXIMM_104_WID_WIDTH),
        .M_AXIMM_105_WID_WIDTH(M_AXIMM_105_WID_WIDTH),
        .M_AXIMM_106_WID_WIDTH(M_AXIMM_106_WID_WIDTH),
        .M_AXIMM_107_WID_WIDTH(M_AXIMM_107_WID_WIDTH),
        .M_AXIMM_108_WID_WIDTH(M_AXIMM_108_WID_WIDTH),
        .M_AXIMM_109_WID_WIDTH(M_AXIMM_109_WID_WIDTH),
        .M_AXIMM_110_WID_WIDTH(M_AXIMM_110_WID_WIDTH),
        .M_AXIMM_111_WID_WIDTH(M_AXIMM_111_WID_WIDTH),
        .M_AXIMM_112_WID_WIDTH(M_AXIMM_112_WID_WIDTH),
        .M_AXIMM_113_WID_WIDTH(M_AXIMM_113_WID_WIDTH),
        .M_AXIMM_114_WID_WIDTH(M_AXIMM_114_WID_WIDTH),
        .M_AXIMM_115_WID_WIDTH(M_AXIMM_115_WID_WIDTH),
        .M_AXIMM_116_WID_WIDTH(M_AXIMM_116_WID_WIDTH),
        .M_AXIMM_117_WID_WIDTH(M_AXIMM_117_WID_WIDTH),
        .M_AXIMM_118_WID_WIDTH(M_AXIMM_118_WID_WIDTH),
        .M_AXIMM_119_WID_WIDTH(M_AXIMM_119_WID_WIDTH),
        .M_AXIMM_120_WID_WIDTH(M_AXIMM_120_WID_WIDTH),
        .M_AXIMM_121_WID_WIDTH(M_AXIMM_121_WID_WIDTH),
        .M_AXIMM_122_WID_WIDTH(M_AXIMM_122_WID_WIDTH),
        .M_AXIMM_123_WID_WIDTH(M_AXIMM_123_WID_WIDTH),
        .M_AXIMM_124_WID_WIDTH(M_AXIMM_124_WID_WIDTH),
        .M_AXIMM_125_WID_WIDTH(M_AXIMM_125_WID_WIDTH),
        .M_AXIMM_126_WID_WIDTH(M_AXIMM_126_WID_WIDTH),
        .M_AXIMM_127_WID_WIDTH(M_AXIMM_127_WID_WIDTH),
        .M_AXIMM_0_BID_WIDTH(M_AXIMM_0_BID_WIDTH),
        .M_AXIMM_1_BID_WIDTH(M_AXIMM_1_BID_WIDTH),
        .M_AXIMM_2_BID_WIDTH(M_AXIMM_2_BID_WIDTH),
        .M_AXIMM_3_BID_WIDTH(M_AXIMM_3_BID_WIDTH),
        .M_AXIMM_4_BID_WIDTH(M_AXIMM_4_BID_WIDTH),
        .M_AXIMM_5_BID_WIDTH(M_AXIMM_5_BID_WIDTH),
        .M_AXIMM_6_BID_WIDTH(M_AXIMM_6_BID_WIDTH),
        .M_AXIMM_7_BID_WIDTH(M_AXIMM_7_BID_WIDTH),
        .M_AXIMM_8_BID_WIDTH(M_AXIMM_8_BID_WIDTH),
        .M_AXIMM_9_BID_WIDTH(M_AXIMM_9_BID_WIDTH),
        .M_AXIMM_10_BID_WIDTH(M_AXIMM_10_BID_WIDTH),
        .M_AXIMM_11_BID_WIDTH(M_AXIMM_11_BID_WIDTH),
        .M_AXIMM_12_BID_WIDTH(M_AXIMM_12_BID_WIDTH),
        .M_AXIMM_13_BID_WIDTH(M_AXIMM_13_BID_WIDTH),
        .M_AXIMM_14_BID_WIDTH(M_AXIMM_14_BID_WIDTH),
        .M_AXIMM_15_BID_WIDTH(M_AXIMM_15_BID_WIDTH),
        .M_AXIMM_16_BID_WIDTH(M_AXIMM_16_BID_WIDTH),
        .M_AXIMM_17_BID_WIDTH(M_AXIMM_17_BID_WIDTH),
        .M_AXIMM_18_BID_WIDTH(M_AXIMM_18_BID_WIDTH),
        .M_AXIMM_19_BID_WIDTH(M_AXIMM_19_BID_WIDTH),
        .M_AXIMM_20_BID_WIDTH(M_AXIMM_20_BID_WIDTH),
        .M_AXIMM_21_BID_WIDTH(M_AXIMM_21_BID_WIDTH),
        .M_AXIMM_22_BID_WIDTH(M_AXIMM_22_BID_WIDTH),
        .M_AXIMM_23_BID_WIDTH(M_AXIMM_23_BID_WIDTH),
        .M_AXIMM_24_BID_WIDTH(M_AXIMM_24_BID_WIDTH),
        .M_AXIMM_25_BID_WIDTH(M_AXIMM_25_BID_WIDTH),
        .M_AXIMM_26_BID_WIDTH(M_AXIMM_26_BID_WIDTH),
        .M_AXIMM_27_BID_WIDTH(M_AXIMM_27_BID_WIDTH),
        .M_AXIMM_28_BID_WIDTH(M_AXIMM_28_BID_WIDTH),
        .M_AXIMM_29_BID_WIDTH(M_AXIMM_29_BID_WIDTH),
        .M_AXIMM_30_BID_WIDTH(M_AXIMM_30_BID_WIDTH),
        .M_AXIMM_31_BID_WIDTH(M_AXIMM_31_BID_WIDTH),
        .M_AXIMM_32_BID_WIDTH(M_AXIMM_32_BID_WIDTH),
        .M_AXIMM_33_BID_WIDTH(M_AXIMM_33_BID_WIDTH),
        .M_AXIMM_34_BID_WIDTH(M_AXIMM_34_BID_WIDTH),
        .M_AXIMM_35_BID_WIDTH(M_AXIMM_35_BID_WIDTH),
        .M_AXIMM_36_BID_WIDTH(M_AXIMM_36_BID_WIDTH),
        .M_AXIMM_37_BID_WIDTH(M_AXIMM_37_BID_WIDTH),
        .M_AXIMM_38_BID_WIDTH(M_AXIMM_38_BID_WIDTH),
        .M_AXIMM_39_BID_WIDTH(M_AXIMM_39_BID_WIDTH),
        .M_AXIMM_40_BID_WIDTH(M_AXIMM_40_BID_WIDTH),
        .M_AXIMM_41_BID_WIDTH(M_AXIMM_41_BID_WIDTH),
        .M_AXIMM_42_BID_WIDTH(M_AXIMM_42_BID_WIDTH),
        .M_AXIMM_43_BID_WIDTH(M_AXIMM_43_BID_WIDTH),
        .M_AXIMM_44_BID_WIDTH(M_AXIMM_44_BID_WIDTH),
        .M_AXIMM_45_BID_WIDTH(M_AXIMM_45_BID_WIDTH),
        .M_AXIMM_46_BID_WIDTH(M_AXIMM_46_BID_WIDTH),
        .M_AXIMM_47_BID_WIDTH(M_AXIMM_47_BID_WIDTH),
        .M_AXIMM_48_BID_WIDTH(M_AXIMM_48_BID_WIDTH),
        .M_AXIMM_49_BID_WIDTH(M_AXIMM_49_BID_WIDTH),
        .M_AXIMM_50_BID_WIDTH(M_AXIMM_50_BID_WIDTH),
        .M_AXIMM_51_BID_WIDTH(M_AXIMM_51_BID_WIDTH),
        .M_AXIMM_52_BID_WIDTH(M_AXIMM_52_BID_WIDTH),
        .M_AXIMM_53_BID_WIDTH(M_AXIMM_53_BID_WIDTH),
        .M_AXIMM_54_BID_WIDTH(M_AXIMM_54_BID_WIDTH),
        .M_AXIMM_55_BID_WIDTH(M_AXIMM_55_BID_WIDTH),
        .M_AXIMM_56_BID_WIDTH(M_AXIMM_56_BID_WIDTH),
        .M_AXIMM_57_BID_WIDTH(M_AXIMM_57_BID_WIDTH),
        .M_AXIMM_58_BID_WIDTH(M_AXIMM_58_BID_WIDTH),
        .M_AXIMM_59_BID_WIDTH(M_AXIMM_59_BID_WIDTH),
        .M_AXIMM_60_BID_WIDTH(M_AXIMM_60_BID_WIDTH),
        .M_AXIMM_61_BID_WIDTH(M_AXIMM_61_BID_WIDTH),
        .M_AXIMM_62_BID_WIDTH(M_AXIMM_62_BID_WIDTH),
        .M_AXIMM_63_BID_WIDTH(M_AXIMM_63_BID_WIDTH),
        .M_AXIMM_64_BID_WIDTH(M_AXIMM_64_BID_WIDTH),
        .M_AXIMM_65_BID_WIDTH(M_AXIMM_65_BID_WIDTH),
        .M_AXIMM_66_BID_WIDTH(M_AXIMM_66_BID_WIDTH),
        .M_AXIMM_67_BID_WIDTH(M_AXIMM_67_BID_WIDTH),
        .M_AXIMM_68_BID_WIDTH(M_AXIMM_68_BID_WIDTH),
        .M_AXIMM_69_BID_WIDTH(M_AXIMM_69_BID_WIDTH),
        .M_AXIMM_70_BID_WIDTH(M_AXIMM_70_BID_WIDTH),
        .M_AXIMM_71_BID_WIDTH(M_AXIMM_71_BID_WIDTH),
        .M_AXIMM_72_BID_WIDTH(M_AXIMM_72_BID_WIDTH),
        .M_AXIMM_73_BID_WIDTH(M_AXIMM_73_BID_WIDTH),
        .M_AXIMM_74_BID_WIDTH(M_AXIMM_74_BID_WIDTH),
        .M_AXIMM_75_BID_WIDTH(M_AXIMM_75_BID_WIDTH),
        .M_AXIMM_76_BID_WIDTH(M_AXIMM_76_BID_WIDTH),
        .M_AXIMM_77_BID_WIDTH(M_AXIMM_77_BID_WIDTH),
        .M_AXIMM_78_BID_WIDTH(M_AXIMM_78_BID_WIDTH),
        .M_AXIMM_79_BID_WIDTH(M_AXIMM_79_BID_WIDTH),
        .M_AXIMM_80_BID_WIDTH(M_AXIMM_80_BID_WIDTH),
        .M_AXIMM_81_BID_WIDTH(M_AXIMM_81_BID_WIDTH),
        .M_AXIMM_82_BID_WIDTH(M_AXIMM_82_BID_WIDTH),
        .M_AXIMM_83_BID_WIDTH(M_AXIMM_83_BID_WIDTH),
        .M_AXIMM_84_BID_WIDTH(M_AXIMM_84_BID_WIDTH),
        .M_AXIMM_85_BID_WIDTH(M_AXIMM_85_BID_WIDTH),
        .M_AXIMM_86_BID_WIDTH(M_AXIMM_86_BID_WIDTH),
        .M_AXIMM_87_BID_WIDTH(M_AXIMM_87_BID_WIDTH),
        .M_AXIMM_88_BID_WIDTH(M_AXIMM_88_BID_WIDTH),
        .M_AXIMM_89_BID_WIDTH(M_AXIMM_89_BID_WIDTH),
        .M_AXIMM_90_BID_WIDTH(M_AXIMM_90_BID_WIDTH),
        .M_AXIMM_91_BID_WIDTH(M_AXIMM_91_BID_WIDTH),
        .M_AXIMM_92_BID_WIDTH(M_AXIMM_92_BID_WIDTH),
        .M_AXIMM_93_BID_WIDTH(M_AXIMM_93_BID_WIDTH),
        .M_AXIMM_94_BID_WIDTH(M_AXIMM_94_BID_WIDTH),
        .M_AXIMM_95_BID_WIDTH(M_AXIMM_95_BID_WIDTH),
        .M_AXIMM_96_BID_WIDTH(M_AXIMM_96_BID_WIDTH),
        .M_AXIMM_97_BID_WIDTH(M_AXIMM_97_BID_WIDTH),
        .M_AXIMM_98_BID_WIDTH(M_AXIMM_98_BID_WIDTH),
        .M_AXIMM_99_BID_WIDTH(M_AXIMM_99_BID_WIDTH),
        .M_AXIMM_100_BID_WIDTH(M_AXIMM_100_BID_WIDTH),
        .M_AXIMM_101_BID_WIDTH(M_AXIMM_101_BID_WIDTH),
        .M_AXIMM_102_BID_WIDTH(M_AXIMM_102_BID_WIDTH),
        .M_AXIMM_103_BID_WIDTH(M_AXIMM_103_BID_WIDTH),
        .M_AXIMM_104_BID_WIDTH(M_AXIMM_104_BID_WIDTH),
        .M_AXIMM_105_BID_WIDTH(M_AXIMM_105_BID_WIDTH),
        .M_AXIMM_106_BID_WIDTH(M_AXIMM_106_BID_WIDTH),
        .M_AXIMM_107_BID_WIDTH(M_AXIMM_107_BID_WIDTH),
        .M_AXIMM_108_BID_WIDTH(M_AXIMM_108_BID_WIDTH),
        .M_AXIMM_109_BID_WIDTH(M_AXIMM_109_BID_WIDTH),
        .M_AXIMM_110_BID_WIDTH(M_AXIMM_110_BID_WIDTH),
        .M_AXIMM_111_BID_WIDTH(M_AXIMM_111_BID_WIDTH),
        .M_AXIMM_112_BID_WIDTH(M_AXIMM_112_BID_WIDTH),
        .M_AXIMM_113_BID_WIDTH(M_AXIMM_113_BID_WIDTH),
        .M_AXIMM_114_BID_WIDTH(M_AXIMM_114_BID_WIDTH),
        .M_AXIMM_115_BID_WIDTH(M_AXIMM_115_BID_WIDTH),
        .M_AXIMM_116_BID_WIDTH(M_AXIMM_116_BID_WIDTH),
        .M_AXIMM_117_BID_WIDTH(M_AXIMM_117_BID_WIDTH),
        .M_AXIMM_118_BID_WIDTH(M_AXIMM_118_BID_WIDTH),
        .M_AXIMM_119_BID_WIDTH(M_AXIMM_119_BID_WIDTH),
        .M_AXIMM_120_BID_WIDTH(M_AXIMM_120_BID_WIDTH),
        .M_AXIMM_121_BID_WIDTH(M_AXIMM_121_BID_WIDTH),
        .M_AXIMM_122_BID_WIDTH(M_AXIMM_122_BID_WIDTH),
        .M_AXIMM_123_BID_WIDTH(M_AXIMM_123_BID_WIDTH),
        .M_AXIMM_124_BID_WIDTH(M_AXIMM_124_BID_WIDTH),
        .M_AXIMM_125_BID_WIDTH(M_AXIMM_125_BID_WIDTH),
        .M_AXIMM_126_BID_WIDTH(M_AXIMM_126_BID_WIDTH),
        .M_AXIMM_127_BID_WIDTH(M_AXIMM_127_BID_WIDTH),
        .M_AXIMM_0_RID_WIDTH(M_AXIMM_0_RID_WIDTH),
        .M_AXIMM_1_RID_WIDTH(M_AXIMM_1_RID_WIDTH),
        .M_AXIMM_2_RID_WIDTH(M_AXIMM_2_RID_WIDTH),
        .M_AXIMM_3_RID_WIDTH(M_AXIMM_3_RID_WIDTH),
        .M_AXIMM_4_RID_WIDTH(M_AXIMM_4_RID_WIDTH),
        .M_AXIMM_5_RID_WIDTH(M_AXIMM_5_RID_WIDTH),
        .M_AXIMM_6_RID_WIDTH(M_AXIMM_6_RID_WIDTH),
        .M_AXIMM_7_RID_WIDTH(M_AXIMM_7_RID_WIDTH),
        .M_AXIMM_8_RID_WIDTH(M_AXIMM_8_RID_WIDTH),
        .M_AXIMM_9_RID_WIDTH(M_AXIMM_9_RID_WIDTH),
        .M_AXIMM_10_RID_WIDTH(M_AXIMM_10_RID_WIDTH),
        .M_AXIMM_11_RID_WIDTH(M_AXIMM_11_RID_WIDTH),
        .M_AXIMM_12_RID_WIDTH(M_AXIMM_12_RID_WIDTH),
        .M_AXIMM_13_RID_WIDTH(M_AXIMM_13_RID_WIDTH),
        .M_AXIMM_14_RID_WIDTH(M_AXIMM_14_RID_WIDTH),
        .M_AXIMM_15_RID_WIDTH(M_AXIMM_15_RID_WIDTH),
        .M_AXIMM_16_RID_WIDTH(M_AXIMM_16_RID_WIDTH),
        .M_AXIMM_17_RID_WIDTH(M_AXIMM_17_RID_WIDTH),
        .M_AXIMM_18_RID_WIDTH(M_AXIMM_18_RID_WIDTH),
        .M_AXIMM_19_RID_WIDTH(M_AXIMM_19_RID_WIDTH),
        .M_AXIMM_20_RID_WIDTH(M_AXIMM_20_RID_WIDTH),
        .M_AXIMM_21_RID_WIDTH(M_AXIMM_21_RID_WIDTH),
        .M_AXIMM_22_RID_WIDTH(M_AXIMM_22_RID_WIDTH),
        .M_AXIMM_23_RID_WIDTH(M_AXIMM_23_RID_WIDTH),
        .M_AXIMM_24_RID_WIDTH(M_AXIMM_24_RID_WIDTH),
        .M_AXIMM_25_RID_WIDTH(M_AXIMM_25_RID_WIDTH),
        .M_AXIMM_26_RID_WIDTH(M_AXIMM_26_RID_WIDTH),
        .M_AXIMM_27_RID_WIDTH(M_AXIMM_27_RID_WIDTH),
        .M_AXIMM_28_RID_WIDTH(M_AXIMM_28_RID_WIDTH),
        .M_AXIMM_29_RID_WIDTH(M_AXIMM_29_RID_WIDTH),
        .M_AXIMM_30_RID_WIDTH(M_AXIMM_30_RID_WIDTH),
        .M_AXIMM_31_RID_WIDTH(M_AXIMM_31_RID_WIDTH),
        .M_AXIMM_32_RID_WIDTH(M_AXIMM_32_RID_WIDTH),
        .M_AXIMM_33_RID_WIDTH(M_AXIMM_33_RID_WIDTH),
        .M_AXIMM_34_RID_WIDTH(M_AXIMM_34_RID_WIDTH),
        .M_AXIMM_35_RID_WIDTH(M_AXIMM_35_RID_WIDTH),
        .M_AXIMM_36_RID_WIDTH(M_AXIMM_36_RID_WIDTH),
        .M_AXIMM_37_RID_WIDTH(M_AXIMM_37_RID_WIDTH),
        .M_AXIMM_38_RID_WIDTH(M_AXIMM_38_RID_WIDTH),
        .M_AXIMM_39_RID_WIDTH(M_AXIMM_39_RID_WIDTH),
        .M_AXIMM_40_RID_WIDTH(M_AXIMM_40_RID_WIDTH),
        .M_AXIMM_41_RID_WIDTH(M_AXIMM_41_RID_WIDTH),
        .M_AXIMM_42_RID_WIDTH(M_AXIMM_42_RID_WIDTH),
        .M_AXIMM_43_RID_WIDTH(M_AXIMM_43_RID_WIDTH),
        .M_AXIMM_44_RID_WIDTH(M_AXIMM_44_RID_WIDTH),
        .M_AXIMM_45_RID_WIDTH(M_AXIMM_45_RID_WIDTH),
        .M_AXIMM_46_RID_WIDTH(M_AXIMM_46_RID_WIDTH),
        .M_AXIMM_47_RID_WIDTH(M_AXIMM_47_RID_WIDTH),
        .M_AXIMM_48_RID_WIDTH(M_AXIMM_48_RID_WIDTH),
        .M_AXIMM_49_RID_WIDTH(M_AXIMM_49_RID_WIDTH),
        .M_AXIMM_50_RID_WIDTH(M_AXIMM_50_RID_WIDTH),
        .M_AXIMM_51_RID_WIDTH(M_AXIMM_51_RID_WIDTH),
        .M_AXIMM_52_RID_WIDTH(M_AXIMM_52_RID_WIDTH),
        .M_AXIMM_53_RID_WIDTH(M_AXIMM_53_RID_WIDTH),
        .M_AXIMM_54_RID_WIDTH(M_AXIMM_54_RID_WIDTH),
        .M_AXIMM_55_RID_WIDTH(M_AXIMM_55_RID_WIDTH),
        .M_AXIMM_56_RID_WIDTH(M_AXIMM_56_RID_WIDTH),
        .M_AXIMM_57_RID_WIDTH(M_AXIMM_57_RID_WIDTH),
        .M_AXIMM_58_RID_WIDTH(M_AXIMM_58_RID_WIDTH),
        .M_AXIMM_59_RID_WIDTH(M_AXIMM_59_RID_WIDTH),
        .M_AXIMM_60_RID_WIDTH(M_AXIMM_60_RID_WIDTH),
        .M_AXIMM_61_RID_WIDTH(M_AXIMM_61_RID_WIDTH),
        .M_AXIMM_62_RID_WIDTH(M_AXIMM_62_RID_WIDTH),
        .M_AXIMM_63_RID_WIDTH(M_AXIMM_63_RID_WIDTH),
        .M_AXIMM_64_RID_WIDTH(M_AXIMM_64_RID_WIDTH),
        .M_AXIMM_65_RID_WIDTH(M_AXIMM_65_RID_WIDTH),
        .M_AXIMM_66_RID_WIDTH(M_AXIMM_66_RID_WIDTH),
        .M_AXIMM_67_RID_WIDTH(M_AXIMM_67_RID_WIDTH),
        .M_AXIMM_68_RID_WIDTH(M_AXIMM_68_RID_WIDTH),
        .M_AXIMM_69_RID_WIDTH(M_AXIMM_69_RID_WIDTH),
        .M_AXIMM_70_RID_WIDTH(M_AXIMM_70_RID_WIDTH),
        .M_AXIMM_71_RID_WIDTH(M_AXIMM_71_RID_WIDTH),
        .M_AXIMM_72_RID_WIDTH(M_AXIMM_72_RID_WIDTH),
        .M_AXIMM_73_RID_WIDTH(M_AXIMM_73_RID_WIDTH),
        .M_AXIMM_74_RID_WIDTH(M_AXIMM_74_RID_WIDTH),
        .M_AXIMM_75_RID_WIDTH(M_AXIMM_75_RID_WIDTH),
        .M_AXIMM_76_RID_WIDTH(M_AXIMM_76_RID_WIDTH),
        .M_AXIMM_77_RID_WIDTH(M_AXIMM_77_RID_WIDTH),
        .M_AXIMM_78_RID_WIDTH(M_AXIMM_78_RID_WIDTH),
        .M_AXIMM_79_RID_WIDTH(M_AXIMM_79_RID_WIDTH),
        .M_AXIMM_80_RID_WIDTH(M_AXIMM_80_RID_WIDTH),
        .M_AXIMM_81_RID_WIDTH(M_AXIMM_81_RID_WIDTH),
        .M_AXIMM_82_RID_WIDTH(M_AXIMM_82_RID_WIDTH),
        .M_AXIMM_83_RID_WIDTH(M_AXIMM_83_RID_WIDTH),
        .M_AXIMM_84_RID_WIDTH(M_AXIMM_84_RID_WIDTH),
        .M_AXIMM_85_RID_WIDTH(M_AXIMM_85_RID_WIDTH),
        .M_AXIMM_86_RID_WIDTH(M_AXIMM_86_RID_WIDTH),
        .M_AXIMM_87_RID_WIDTH(M_AXIMM_87_RID_WIDTH),
        .M_AXIMM_88_RID_WIDTH(M_AXIMM_88_RID_WIDTH),
        .M_AXIMM_89_RID_WIDTH(M_AXIMM_89_RID_WIDTH),
        .M_AXIMM_90_RID_WIDTH(M_AXIMM_90_RID_WIDTH),
        .M_AXIMM_91_RID_WIDTH(M_AXIMM_91_RID_WIDTH),
        .M_AXIMM_92_RID_WIDTH(M_AXIMM_92_RID_WIDTH),
        .M_AXIMM_93_RID_WIDTH(M_AXIMM_93_RID_WIDTH),
        .M_AXIMM_94_RID_WIDTH(M_AXIMM_94_RID_WIDTH),
        .M_AXIMM_95_RID_WIDTH(M_AXIMM_95_RID_WIDTH),
        .M_AXIMM_96_RID_WIDTH(M_AXIMM_96_RID_WIDTH),
        .M_AXIMM_97_RID_WIDTH(M_AXIMM_97_RID_WIDTH),
        .M_AXIMM_98_RID_WIDTH(M_AXIMM_98_RID_WIDTH),
        .M_AXIMM_99_RID_WIDTH(M_AXIMM_99_RID_WIDTH),
        .M_AXIMM_100_RID_WIDTH(M_AXIMM_100_RID_WIDTH),
        .M_AXIMM_101_RID_WIDTH(M_AXIMM_101_RID_WIDTH),
        .M_AXIMM_102_RID_WIDTH(M_AXIMM_102_RID_WIDTH),
        .M_AXIMM_103_RID_WIDTH(M_AXIMM_103_RID_WIDTH),
        .M_AXIMM_104_RID_WIDTH(M_AXIMM_104_RID_WIDTH),
        .M_AXIMM_105_RID_WIDTH(M_AXIMM_105_RID_WIDTH),
        .M_AXIMM_106_RID_WIDTH(M_AXIMM_106_RID_WIDTH),
        .M_AXIMM_107_RID_WIDTH(M_AXIMM_107_RID_WIDTH),
        .M_AXIMM_108_RID_WIDTH(M_AXIMM_108_RID_WIDTH),
        .M_AXIMM_109_RID_WIDTH(M_AXIMM_109_RID_WIDTH),
        .M_AXIMM_110_RID_WIDTH(M_AXIMM_110_RID_WIDTH),
        .M_AXIMM_111_RID_WIDTH(M_AXIMM_111_RID_WIDTH),
        .M_AXIMM_112_RID_WIDTH(M_AXIMM_112_RID_WIDTH),
        .M_AXIMM_113_RID_WIDTH(M_AXIMM_113_RID_WIDTH),
        .M_AXIMM_114_RID_WIDTH(M_AXIMM_114_RID_WIDTH),
        .M_AXIMM_115_RID_WIDTH(M_AXIMM_115_RID_WIDTH),
        .M_AXIMM_116_RID_WIDTH(M_AXIMM_116_RID_WIDTH),
        .M_AXIMM_117_RID_WIDTH(M_AXIMM_117_RID_WIDTH),
        .M_AXIMM_118_RID_WIDTH(M_AXIMM_118_RID_WIDTH),
        .M_AXIMM_119_RID_WIDTH(M_AXIMM_119_RID_WIDTH),
        .M_AXIMM_120_RID_WIDTH(M_AXIMM_120_RID_WIDTH),
        .M_AXIMM_121_RID_WIDTH(M_AXIMM_121_RID_WIDTH),
        .M_AXIMM_122_RID_WIDTH(M_AXIMM_122_RID_WIDTH),
        .M_AXIMM_123_RID_WIDTH(M_AXIMM_123_RID_WIDTH),
        .M_AXIMM_124_RID_WIDTH(M_AXIMM_124_RID_WIDTH),
        .M_AXIMM_125_RID_WIDTH(M_AXIMM_125_RID_WIDTH),
        .M_AXIMM_126_RID_WIDTH(M_AXIMM_126_RID_WIDTH),
        .M_AXIMM_127_RID_WIDTH(M_AXIMM_127_RID_WIDTH),
        .M_AXIMM_0_DATA_WIDTH(M_AXIMM_0_DATA_WIDTH),
        .M_AXIMM_1_DATA_WIDTH(M_AXIMM_1_DATA_WIDTH),
        .M_AXIMM_2_DATA_WIDTH(M_AXIMM_2_DATA_WIDTH),
        .M_AXIMM_3_DATA_WIDTH(M_AXIMM_3_DATA_WIDTH),
        .M_AXIMM_4_DATA_WIDTH(M_AXIMM_4_DATA_WIDTH),
        .M_AXIMM_5_DATA_WIDTH(M_AXIMM_5_DATA_WIDTH),
        .M_AXIMM_6_DATA_WIDTH(M_AXIMM_6_DATA_WIDTH),
        .M_AXIMM_7_DATA_WIDTH(M_AXIMM_7_DATA_WIDTH),
        .M_AXIMM_8_DATA_WIDTH(M_AXIMM_8_DATA_WIDTH),
        .M_AXIMM_9_DATA_WIDTH(M_AXIMM_9_DATA_WIDTH),
        .M_AXIMM_10_DATA_WIDTH(M_AXIMM_10_DATA_WIDTH),
        .M_AXIMM_11_DATA_WIDTH(M_AXIMM_11_DATA_WIDTH),
        .M_AXIMM_12_DATA_WIDTH(M_AXIMM_12_DATA_WIDTH),
        .M_AXIMM_13_DATA_WIDTH(M_AXIMM_13_DATA_WIDTH),
        .M_AXIMM_14_DATA_WIDTH(M_AXIMM_14_DATA_WIDTH),
        .M_AXIMM_15_DATA_WIDTH(M_AXIMM_15_DATA_WIDTH),
        .M_AXIMM_16_DATA_WIDTH(M_AXIMM_16_DATA_WIDTH),
        .M_AXIMM_17_DATA_WIDTH(M_AXIMM_17_DATA_WIDTH),
        .M_AXIMM_18_DATA_WIDTH(M_AXIMM_18_DATA_WIDTH),
        .M_AXIMM_19_DATA_WIDTH(M_AXIMM_19_DATA_WIDTH),
        .M_AXIMM_20_DATA_WIDTH(M_AXIMM_20_DATA_WIDTH),
        .M_AXIMM_21_DATA_WIDTH(M_AXIMM_21_DATA_WIDTH),
        .M_AXIMM_22_DATA_WIDTH(M_AXIMM_22_DATA_WIDTH),
        .M_AXIMM_23_DATA_WIDTH(M_AXIMM_23_DATA_WIDTH),
        .M_AXIMM_24_DATA_WIDTH(M_AXIMM_24_DATA_WIDTH),
        .M_AXIMM_25_DATA_WIDTH(M_AXIMM_25_DATA_WIDTH),
        .M_AXIMM_26_DATA_WIDTH(M_AXIMM_26_DATA_WIDTH),
        .M_AXIMM_27_DATA_WIDTH(M_AXIMM_27_DATA_WIDTH),
        .M_AXIMM_28_DATA_WIDTH(M_AXIMM_28_DATA_WIDTH),
        .M_AXIMM_29_DATA_WIDTH(M_AXIMM_29_DATA_WIDTH),
        .M_AXIMM_30_DATA_WIDTH(M_AXIMM_30_DATA_WIDTH),
        .M_AXIMM_31_DATA_WIDTH(M_AXIMM_31_DATA_WIDTH),
        .M_AXIMM_32_DATA_WIDTH(M_AXIMM_32_DATA_WIDTH),
        .M_AXIMM_33_DATA_WIDTH(M_AXIMM_33_DATA_WIDTH),
        .M_AXIMM_34_DATA_WIDTH(M_AXIMM_34_DATA_WIDTH),
        .M_AXIMM_35_DATA_WIDTH(M_AXIMM_35_DATA_WIDTH),
        .M_AXIMM_36_DATA_WIDTH(M_AXIMM_36_DATA_WIDTH),
        .M_AXIMM_37_DATA_WIDTH(M_AXIMM_37_DATA_WIDTH),
        .M_AXIMM_38_DATA_WIDTH(M_AXIMM_38_DATA_WIDTH),
        .M_AXIMM_39_DATA_WIDTH(M_AXIMM_39_DATA_WIDTH),
        .M_AXIMM_40_DATA_WIDTH(M_AXIMM_40_DATA_WIDTH),
        .M_AXIMM_41_DATA_WIDTH(M_AXIMM_41_DATA_WIDTH),
        .M_AXIMM_42_DATA_WIDTH(M_AXIMM_42_DATA_WIDTH),
        .M_AXIMM_43_DATA_WIDTH(M_AXIMM_43_DATA_WIDTH),
        .M_AXIMM_44_DATA_WIDTH(M_AXIMM_44_DATA_WIDTH),
        .M_AXIMM_45_DATA_WIDTH(M_AXIMM_45_DATA_WIDTH),
        .M_AXIMM_46_DATA_WIDTH(M_AXIMM_46_DATA_WIDTH),
        .M_AXIMM_47_DATA_WIDTH(M_AXIMM_47_DATA_WIDTH),
        .M_AXIMM_48_DATA_WIDTH(M_AXIMM_48_DATA_WIDTH),
        .M_AXIMM_49_DATA_WIDTH(M_AXIMM_49_DATA_WIDTH),
        .M_AXIMM_50_DATA_WIDTH(M_AXIMM_50_DATA_WIDTH),
        .M_AXIMM_51_DATA_WIDTH(M_AXIMM_51_DATA_WIDTH),
        .M_AXIMM_52_DATA_WIDTH(M_AXIMM_52_DATA_WIDTH),
        .M_AXIMM_53_DATA_WIDTH(M_AXIMM_53_DATA_WIDTH),
        .M_AXIMM_54_DATA_WIDTH(M_AXIMM_54_DATA_WIDTH),
        .M_AXIMM_55_DATA_WIDTH(M_AXIMM_55_DATA_WIDTH),
        .M_AXIMM_56_DATA_WIDTH(M_AXIMM_56_DATA_WIDTH),
        .M_AXIMM_57_DATA_WIDTH(M_AXIMM_57_DATA_WIDTH),
        .M_AXIMM_58_DATA_WIDTH(M_AXIMM_58_DATA_WIDTH),
        .M_AXIMM_59_DATA_WIDTH(M_AXIMM_59_DATA_WIDTH),
        .M_AXIMM_60_DATA_WIDTH(M_AXIMM_60_DATA_WIDTH),
        .M_AXIMM_61_DATA_WIDTH(M_AXIMM_61_DATA_WIDTH),
        .M_AXIMM_62_DATA_WIDTH(M_AXIMM_62_DATA_WIDTH),
        .M_AXIMM_63_DATA_WIDTH(M_AXIMM_63_DATA_WIDTH),
        .M_AXIMM_64_DATA_WIDTH(M_AXIMM_64_DATA_WIDTH),
        .M_AXIMM_65_DATA_WIDTH(M_AXIMM_65_DATA_WIDTH),
        .M_AXIMM_66_DATA_WIDTH(M_AXIMM_66_DATA_WIDTH),
        .M_AXIMM_67_DATA_WIDTH(M_AXIMM_67_DATA_WIDTH),
        .M_AXIMM_68_DATA_WIDTH(M_AXIMM_68_DATA_WIDTH),
        .M_AXIMM_69_DATA_WIDTH(M_AXIMM_69_DATA_WIDTH),
        .M_AXIMM_70_DATA_WIDTH(M_AXIMM_70_DATA_WIDTH),
        .M_AXIMM_71_DATA_WIDTH(M_AXIMM_71_DATA_WIDTH),
        .M_AXIMM_72_DATA_WIDTH(M_AXIMM_72_DATA_WIDTH),
        .M_AXIMM_73_DATA_WIDTH(M_AXIMM_73_DATA_WIDTH),
        .M_AXIMM_74_DATA_WIDTH(M_AXIMM_74_DATA_WIDTH),
        .M_AXIMM_75_DATA_WIDTH(M_AXIMM_75_DATA_WIDTH),
        .M_AXIMM_76_DATA_WIDTH(M_AXIMM_76_DATA_WIDTH),
        .M_AXIMM_77_DATA_WIDTH(M_AXIMM_77_DATA_WIDTH),
        .M_AXIMM_78_DATA_WIDTH(M_AXIMM_78_DATA_WIDTH),
        .M_AXIMM_79_DATA_WIDTH(M_AXIMM_79_DATA_WIDTH),
        .M_AXIMM_80_DATA_WIDTH(M_AXIMM_80_DATA_WIDTH),
        .M_AXIMM_81_DATA_WIDTH(M_AXIMM_81_DATA_WIDTH),
        .M_AXIMM_82_DATA_WIDTH(M_AXIMM_82_DATA_WIDTH),
        .M_AXIMM_83_DATA_WIDTH(M_AXIMM_83_DATA_WIDTH),
        .M_AXIMM_84_DATA_WIDTH(M_AXIMM_84_DATA_WIDTH),
        .M_AXIMM_85_DATA_WIDTH(M_AXIMM_85_DATA_WIDTH),
        .M_AXIMM_86_DATA_WIDTH(M_AXIMM_86_DATA_WIDTH),
        .M_AXIMM_87_DATA_WIDTH(M_AXIMM_87_DATA_WIDTH),
        .M_AXIMM_88_DATA_WIDTH(M_AXIMM_88_DATA_WIDTH),
        .M_AXIMM_89_DATA_WIDTH(M_AXIMM_89_DATA_WIDTH),
        .M_AXIMM_90_DATA_WIDTH(M_AXIMM_90_DATA_WIDTH),
        .M_AXIMM_91_DATA_WIDTH(M_AXIMM_91_DATA_WIDTH),
        .M_AXIMM_92_DATA_WIDTH(M_AXIMM_92_DATA_WIDTH),
        .M_AXIMM_93_DATA_WIDTH(M_AXIMM_93_DATA_WIDTH),
        .M_AXIMM_94_DATA_WIDTH(M_AXIMM_94_DATA_WIDTH),
        .M_AXIMM_95_DATA_WIDTH(M_AXIMM_95_DATA_WIDTH),
        .M_AXIMM_96_DATA_WIDTH(M_AXIMM_96_DATA_WIDTH),
        .M_AXIMM_97_DATA_WIDTH(M_AXIMM_97_DATA_WIDTH),
        .M_AXIMM_98_DATA_WIDTH(M_AXIMM_98_DATA_WIDTH),
        .M_AXIMM_99_DATA_WIDTH(M_AXIMM_99_DATA_WIDTH),
        .M_AXIMM_100_DATA_WIDTH(M_AXIMM_100_DATA_WIDTH),
        .M_AXIMM_101_DATA_WIDTH(M_AXIMM_101_DATA_WIDTH),
        .M_AXIMM_102_DATA_WIDTH(M_AXIMM_102_DATA_WIDTH),
        .M_AXIMM_103_DATA_WIDTH(M_AXIMM_103_DATA_WIDTH),
        .M_AXIMM_104_DATA_WIDTH(M_AXIMM_104_DATA_WIDTH),
        .M_AXIMM_105_DATA_WIDTH(M_AXIMM_105_DATA_WIDTH),
        .M_AXIMM_106_DATA_WIDTH(M_AXIMM_106_DATA_WIDTH),
        .M_AXIMM_107_DATA_WIDTH(M_AXIMM_107_DATA_WIDTH),
        .M_AXIMM_108_DATA_WIDTH(M_AXIMM_108_DATA_WIDTH),
        .M_AXIMM_109_DATA_WIDTH(M_AXIMM_109_DATA_WIDTH),
        .M_AXIMM_110_DATA_WIDTH(M_AXIMM_110_DATA_WIDTH),
        .M_AXIMM_111_DATA_WIDTH(M_AXIMM_111_DATA_WIDTH),
        .M_AXIMM_112_DATA_WIDTH(M_AXIMM_112_DATA_WIDTH),
        .M_AXIMM_113_DATA_WIDTH(M_AXIMM_113_DATA_WIDTH),
        .M_AXIMM_114_DATA_WIDTH(M_AXIMM_114_DATA_WIDTH),
        .M_AXIMM_115_DATA_WIDTH(M_AXIMM_115_DATA_WIDTH),
        .M_AXIMM_116_DATA_WIDTH(M_AXIMM_116_DATA_WIDTH),
        .M_AXIMM_117_DATA_WIDTH(M_AXIMM_117_DATA_WIDTH),
        .M_AXIMM_118_DATA_WIDTH(M_AXIMM_118_DATA_WIDTH),
        .M_AXIMM_119_DATA_WIDTH(M_AXIMM_119_DATA_WIDTH),
        .M_AXIMM_120_DATA_WIDTH(M_AXIMM_120_DATA_WIDTH),
        .M_AXIMM_121_DATA_WIDTH(M_AXIMM_121_DATA_WIDTH),
        .M_AXIMM_122_DATA_WIDTH(M_AXIMM_122_DATA_WIDTH),
        .M_AXIMM_123_DATA_WIDTH(M_AXIMM_123_DATA_WIDTH),
        .M_AXIMM_124_DATA_WIDTH(M_AXIMM_124_DATA_WIDTH),
        .M_AXIMM_125_DATA_WIDTH(M_AXIMM_125_DATA_WIDTH),
        .M_AXIMM_126_DATA_WIDTH(M_AXIMM_126_DATA_WIDTH),
        .M_AXIMM_127_DATA_WIDTH(M_AXIMM_127_DATA_WIDTH)
    ) aximm_args_i (
        .acc_clk(acc_aclk),
        .dm_clk(s_axi_aclk),
        .aresetn(s_axi_aresetn),
        .AP_AXIMM_0_AWADDR(AP_AXIMM_0_AWADDR),
        .AP_AXIMM_0_AWLEN(AP_AXIMM_0_AWLEN),
        .AP_AXIMM_0_AWSIZE(AP_AXIMM_0_AWSIZE),
        .AP_AXIMM_0_AWBURST(AP_AXIMM_0_AWBURST),
        .AP_AXIMM_0_AWLOCK(AP_AXIMM_0_AWLOCK),
        .AP_AXIMM_0_AWCACHE(AP_AXIMM_0_AWCACHE),
        .AP_AXIMM_0_AWPROT(AP_AXIMM_0_AWPROT),
        .AP_AXIMM_0_AWREGION(AP_AXIMM_0_AWREGION),
        .AP_AXIMM_0_AWQOS(AP_AXIMM_0_AWQOS),
        .AP_AXIMM_0_AWVALID(AP_AXIMM_0_AWVALID),
        .AP_AXIMM_0_AWREADY(AP_AXIMM_0_AWREADY),
        .AP_AXIMM_0_WDATA(AP_AXIMM_0_WDATA),
        .AP_AXIMM_0_WSTRB(AP_AXIMM_0_WSTRB),
        .AP_AXIMM_0_WLAST(AP_AXIMM_0_WLAST),
        .AP_AXIMM_0_WVALID(AP_AXIMM_0_WVALID),
        .AP_AXIMM_0_WREADY(AP_AXIMM_0_WREADY),
        .AP_AXIMM_0_BRESP(AP_AXIMM_0_BRESP),
        .AP_AXIMM_0_BVALID(AP_AXIMM_0_BVALID),
        .AP_AXIMM_0_BREADY(AP_AXIMM_0_BREADY),
        .AP_AXIMM_0_ARADDR(AP_AXIMM_0_ARADDR),
        .AP_AXIMM_0_ARLEN(AP_AXIMM_0_ARLEN),
        .AP_AXIMM_0_ARSIZE(AP_AXIMM_0_ARSIZE),
        .AP_AXIMM_0_ARBURST(AP_AXIMM_0_ARBURST),
        .AP_AXIMM_0_ARLOCK(AP_AXIMM_0_ARLOCK),
        .AP_AXIMM_0_ARCACHE(AP_AXIMM_0_ARCACHE),
        .AP_AXIMM_0_ARPROT(AP_AXIMM_0_ARPROT),
        .AP_AXIMM_0_ARREGION(AP_AXIMM_0_ARREGION),
        .AP_AXIMM_0_ARQOS(AP_AXIMM_0_ARQOS),
        .AP_AXIMM_0_ARVALID(AP_AXIMM_0_ARVALID),
        .AP_AXIMM_0_ARREADY(AP_AXIMM_0_ARREADY),
        .AP_AXIMM_0_RDATA(AP_AXIMM_0_RDATA),
        .AP_AXIMM_0_RRESP(AP_AXIMM_0_RRESP),
        .AP_AXIMM_0_RLAST(AP_AXIMM_0_RLAST),
        .AP_AXIMM_0_RVALID(AP_AXIMM_0_RVALID),
        .AP_AXIMM_0_RREADY(AP_AXIMM_0_RREADY),
        .M_AXIMM_0_AWADDR(M_AXIMM_0_AWADDR),
        .M_AXIMM_0_AWLEN(M_AXIMM_0_AWLEN),
        .M_AXIMM_0_AWSIZE(M_AXIMM_0_AWSIZE),
        .M_AXIMM_0_AWBURST(M_AXIMM_0_AWBURST),
        .M_AXIMM_0_AWLOCK(M_AXIMM_0_AWLOCK),
        .M_AXIMM_0_AWCACHE(M_AXIMM_0_AWCACHE),
        .M_AXIMM_0_AWPROT(M_AXIMM_0_AWPROT),
        .M_AXIMM_0_AWREGION(M_AXIMM_0_AWREGION),
        .M_AXIMM_0_AWQOS(M_AXIMM_0_AWQOS),
        .M_AXIMM_0_AWVALID(M_AXIMM_0_AWVALID),
        .M_AXIMM_0_AWREADY(M_AXIMM_0_AWREADY),
        .M_AXIMM_0_WDATA(M_AXIMM_0_WDATA),
        .M_AXIMM_0_WSTRB(M_AXIMM_0_WSTRB),
        .M_AXIMM_0_WLAST(M_AXIMM_0_WLAST),
        .M_AXIMM_0_WVALID(M_AXIMM_0_WVALID),
        .M_AXIMM_0_WREADY(M_AXIMM_0_WREADY),
        .M_AXIMM_0_BRESP(M_AXIMM_0_BRESP),
        .M_AXIMM_0_BVALID(M_AXIMM_0_BVALID),
        .M_AXIMM_0_BREADY(M_AXIMM_0_BREADY),
        .M_AXIMM_0_ARADDR(M_AXIMM_0_ARADDR),
        .M_AXIMM_0_ARLEN(M_AXIMM_0_ARLEN),
        .M_AXIMM_0_ARSIZE(M_AXIMM_0_ARSIZE),
        .M_AXIMM_0_ARBURST(M_AXIMM_0_ARBURST),
        .M_AXIMM_0_ARLOCK(M_AXIMM_0_ARLOCK),
        .M_AXIMM_0_ARCACHE(M_AXIMM_0_ARCACHE),
        .M_AXIMM_0_ARPROT(M_AXIMM_0_ARPROT),
        .M_AXIMM_0_ARREGION(M_AXIMM_0_ARREGION),
        .M_AXIMM_0_ARQOS(M_AXIMM_0_ARQOS),
        .M_AXIMM_0_ARVALID(M_AXIMM_0_ARVALID),
        .M_AXIMM_0_ARREADY(M_AXIMM_0_ARREADY),
        .M_AXIMM_0_RDATA(M_AXIMM_0_RDATA),
        .M_AXIMM_0_RRESP(M_AXIMM_0_RRESP),
        .M_AXIMM_0_RLAST(M_AXIMM_0_RLAST),
        .M_AXIMM_0_RVALID(M_AXIMM_0_RVALID),
        .M_AXIMM_0_RREADY(M_AXIMM_0_RREADY),
        .AP_AXIMM_1_AWADDR(AP_AXIMM_1_AWADDR),
        .AP_AXIMM_1_AWLEN(AP_AXIMM_1_AWLEN),
        .AP_AXIMM_1_AWSIZE(AP_AXIMM_1_AWSIZE),
        .AP_AXIMM_1_AWBURST(AP_AXIMM_1_AWBURST),
        .AP_AXIMM_1_AWLOCK(AP_AXIMM_1_AWLOCK),
        .AP_AXIMM_1_AWCACHE(AP_AXIMM_1_AWCACHE),
        .AP_AXIMM_1_AWPROT(AP_AXIMM_1_AWPROT),
        .AP_AXIMM_1_AWREGION(AP_AXIMM_1_AWREGION),
        .AP_AXIMM_1_AWQOS(AP_AXIMM_1_AWQOS),
        .AP_AXIMM_1_AWVALID(AP_AXIMM_1_AWVALID),
        .AP_AXIMM_1_AWREADY(AP_AXIMM_1_AWREADY),
        .AP_AXIMM_1_WDATA(AP_AXIMM_1_WDATA),
        .AP_AXIMM_1_WSTRB(AP_AXIMM_1_WSTRB),
        .AP_AXIMM_1_WLAST(AP_AXIMM_1_WLAST),
        .AP_AXIMM_1_WVALID(AP_AXIMM_1_WVALID),
        .AP_AXIMM_1_WREADY(AP_AXIMM_1_WREADY),
        .AP_AXIMM_1_BRESP(AP_AXIMM_1_BRESP),
        .AP_AXIMM_1_BVALID(AP_AXIMM_1_BVALID),
        .AP_AXIMM_1_BREADY(AP_AXIMM_1_BREADY),
        .AP_AXIMM_1_ARADDR(AP_AXIMM_1_ARADDR),
        .AP_AXIMM_1_ARLEN(AP_AXIMM_1_ARLEN),
        .AP_AXIMM_1_ARSIZE(AP_AXIMM_1_ARSIZE),
        .AP_AXIMM_1_ARBURST(AP_AXIMM_1_ARBURST),
        .AP_AXIMM_1_ARLOCK(AP_AXIMM_1_ARLOCK),
        .AP_AXIMM_1_ARCACHE(AP_AXIMM_1_ARCACHE),
        .AP_AXIMM_1_ARPROT(AP_AXIMM_1_ARPROT),
        .AP_AXIMM_1_ARREGION(AP_AXIMM_1_ARREGION),
        .AP_AXIMM_1_ARQOS(AP_AXIMM_1_ARQOS),
        .AP_AXIMM_1_ARVALID(AP_AXIMM_1_ARVALID),
        .AP_AXIMM_1_ARREADY(AP_AXIMM_1_ARREADY),
        .AP_AXIMM_1_RDATA(AP_AXIMM_1_RDATA),
        .AP_AXIMM_1_RRESP(AP_AXIMM_1_RRESP),
        .AP_AXIMM_1_RLAST(AP_AXIMM_1_RLAST),
        .AP_AXIMM_1_RVALID(AP_AXIMM_1_RVALID),
        .AP_AXIMM_1_RREADY(AP_AXIMM_1_RREADY),
        .M_AXIMM_1_AWADDR(M_AXIMM_1_AWADDR),
        .M_AXIMM_1_AWLEN(M_AXIMM_1_AWLEN),
        .M_AXIMM_1_AWSIZE(M_AXIMM_1_AWSIZE),
        .M_AXIMM_1_AWBURST(M_AXIMM_1_AWBURST),
        .M_AXIMM_1_AWLOCK(M_AXIMM_1_AWLOCK),
        .M_AXIMM_1_AWCACHE(M_AXIMM_1_AWCACHE),
        .M_AXIMM_1_AWPROT(M_AXIMM_1_AWPROT),
        .M_AXIMM_1_AWREGION(M_AXIMM_1_AWREGION),
        .M_AXIMM_1_AWQOS(M_AXIMM_1_AWQOS),
        .M_AXIMM_1_AWVALID(M_AXIMM_1_AWVALID),
        .M_AXIMM_1_AWREADY(M_AXIMM_1_AWREADY),
        .M_AXIMM_1_WDATA(M_AXIMM_1_WDATA),
        .M_AXIMM_1_WSTRB(M_AXIMM_1_WSTRB),
        .M_AXIMM_1_WLAST(M_AXIMM_1_WLAST),
        .M_AXIMM_1_WVALID(M_AXIMM_1_WVALID),
        .M_AXIMM_1_WREADY(M_AXIMM_1_WREADY),
        .M_AXIMM_1_BRESP(M_AXIMM_1_BRESP),
        .M_AXIMM_1_BVALID(M_AXIMM_1_BVALID),
        .M_AXIMM_1_BREADY(M_AXIMM_1_BREADY),
        .M_AXIMM_1_ARADDR(M_AXIMM_1_ARADDR),
        .M_AXIMM_1_ARLEN(M_AXIMM_1_ARLEN),
        .M_AXIMM_1_ARSIZE(M_AXIMM_1_ARSIZE),
        .M_AXIMM_1_ARBURST(M_AXIMM_1_ARBURST),
        .M_AXIMM_1_ARLOCK(M_AXIMM_1_ARLOCK),
        .M_AXIMM_1_ARCACHE(M_AXIMM_1_ARCACHE),
        .M_AXIMM_1_ARPROT(M_AXIMM_1_ARPROT),
        .M_AXIMM_1_ARREGION(M_AXIMM_1_ARREGION),
        .M_AXIMM_1_ARQOS(M_AXIMM_1_ARQOS),
        .M_AXIMM_1_ARVALID(M_AXIMM_1_ARVALID),
        .M_AXIMM_1_ARREADY(M_AXIMM_1_ARREADY),
        .M_AXIMM_1_RDATA(M_AXIMM_1_RDATA),
        .M_AXIMM_1_RRESP(M_AXIMM_1_RRESP),
        .M_AXIMM_1_RLAST(M_AXIMM_1_RLAST),
        .M_AXIMM_1_RVALID(M_AXIMM_1_RVALID),
        .M_AXIMM_1_RREADY(M_AXIMM_1_RREADY),
        .AP_AXIMM_2_AWADDR(AP_AXIMM_2_AWADDR),
        .AP_AXIMM_2_AWLEN(AP_AXIMM_2_AWLEN),
        .AP_AXIMM_2_AWSIZE(AP_AXIMM_2_AWSIZE),
        .AP_AXIMM_2_AWBURST(AP_AXIMM_2_AWBURST),
        .AP_AXIMM_2_AWLOCK(AP_AXIMM_2_AWLOCK),
        .AP_AXIMM_2_AWCACHE(AP_AXIMM_2_AWCACHE),
        .AP_AXIMM_2_AWPROT(AP_AXIMM_2_AWPROT),
        .AP_AXIMM_2_AWREGION(AP_AXIMM_2_AWREGION),
        .AP_AXIMM_2_AWQOS(AP_AXIMM_2_AWQOS),
        .AP_AXIMM_2_AWVALID(AP_AXIMM_2_AWVALID),
        .AP_AXIMM_2_AWREADY(AP_AXIMM_2_AWREADY),
        .AP_AXIMM_2_WDATA(AP_AXIMM_2_WDATA),
        .AP_AXIMM_2_WSTRB(AP_AXIMM_2_WSTRB),
        .AP_AXIMM_2_WLAST(AP_AXIMM_2_WLAST),
        .AP_AXIMM_2_WVALID(AP_AXIMM_2_WVALID),
        .AP_AXIMM_2_WREADY(AP_AXIMM_2_WREADY),
        .AP_AXIMM_2_BRESP(AP_AXIMM_2_BRESP),
        .AP_AXIMM_2_BVALID(AP_AXIMM_2_BVALID),
        .AP_AXIMM_2_BREADY(AP_AXIMM_2_BREADY),
        .AP_AXIMM_2_ARADDR(AP_AXIMM_2_ARADDR),
        .AP_AXIMM_2_ARLEN(AP_AXIMM_2_ARLEN),
        .AP_AXIMM_2_ARSIZE(AP_AXIMM_2_ARSIZE),
        .AP_AXIMM_2_ARBURST(AP_AXIMM_2_ARBURST),
        .AP_AXIMM_2_ARLOCK(AP_AXIMM_2_ARLOCK),
        .AP_AXIMM_2_ARCACHE(AP_AXIMM_2_ARCACHE),
        .AP_AXIMM_2_ARPROT(AP_AXIMM_2_ARPROT),
        .AP_AXIMM_2_ARREGION(AP_AXIMM_2_ARREGION),
        .AP_AXIMM_2_ARQOS(AP_AXIMM_2_ARQOS),
        .AP_AXIMM_2_ARVALID(AP_AXIMM_2_ARVALID),
        .AP_AXIMM_2_ARREADY(AP_AXIMM_2_ARREADY),
        .AP_AXIMM_2_RDATA(AP_AXIMM_2_RDATA),
        .AP_AXIMM_2_RRESP(AP_AXIMM_2_RRESP),
        .AP_AXIMM_2_RLAST(AP_AXIMM_2_RLAST),
        .AP_AXIMM_2_RVALID(AP_AXIMM_2_RVALID),
        .AP_AXIMM_2_RREADY(AP_AXIMM_2_RREADY),
        .M_AXIMM_2_AWADDR(M_AXIMM_2_AWADDR),
        .M_AXIMM_2_AWLEN(M_AXIMM_2_AWLEN),
        .M_AXIMM_2_AWSIZE(M_AXIMM_2_AWSIZE),
        .M_AXIMM_2_AWBURST(M_AXIMM_2_AWBURST),
        .M_AXIMM_2_AWLOCK(M_AXIMM_2_AWLOCK),
        .M_AXIMM_2_AWCACHE(M_AXIMM_2_AWCACHE),
        .M_AXIMM_2_AWPROT(M_AXIMM_2_AWPROT),
        .M_AXIMM_2_AWREGION(M_AXIMM_2_AWREGION),
        .M_AXIMM_2_AWQOS(M_AXIMM_2_AWQOS),
        .M_AXIMM_2_AWVALID(M_AXIMM_2_AWVALID),
        .M_AXIMM_2_AWREADY(M_AXIMM_2_AWREADY),
        .M_AXIMM_2_WDATA(M_AXIMM_2_WDATA),
        .M_AXIMM_2_WSTRB(M_AXIMM_2_WSTRB),
        .M_AXIMM_2_WLAST(M_AXIMM_2_WLAST),
        .M_AXIMM_2_WVALID(M_AXIMM_2_WVALID),
        .M_AXIMM_2_WREADY(M_AXIMM_2_WREADY),
        .M_AXIMM_2_BRESP(M_AXIMM_2_BRESP),
        .M_AXIMM_2_BVALID(M_AXIMM_2_BVALID),
        .M_AXIMM_2_BREADY(M_AXIMM_2_BREADY),
        .M_AXIMM_2_ARADDR(M_AXIMM_2_ARADDR),
        .M_AXIMM_2_ARLEN(M_AXIMM_2_ARLEN),
        .M_AXIMM_2_ARSIZE(M_AXIMM_2_ARSIZE),
        .M_AXIMM_2_ARBURST(M_AXIMM_2_ARBURST),
        .M_AXIMM_2_ARLOCK(M_AXIMM_2_ARLOCK),
        .M_AXIMM_2_ARCACHE(M_AXIMM_2_ARCACHE),
        .M_AXIMM_2_ARPROT(M_AXIMM_2_ARPROT),
        .M_AXIMM_2_ARREGION(M_AXIMM_2_ARREGION),
        .M_AXIMM_2_ARQOS(M_AXIMM_2_ARQOS),
        .M_AXIMM_2_ARVALID(M_AXIMM_2_ARVALID),
        .M_AXIMM_2_ARREADY(M_AXIMM_2_ARREADY),
        .M_AXIMM_2_RDATA(M_AXIMM_2_RDATA),
        .M_AXIMM_2_RRESP(M_AXIMM_2_RRESP),
        .M_AXIMM_2_RLAST(M_AXIMM_2_RLAST),
        .M_AXIMM_2_RVALID(M_AXIMM_2_RVALID),
        .M_AXIMM_2_RREADY(M_AXIMM_2_RREADY),
        .AP_AXIMM_3_AWADDR(AP_AXIMM_3_AWADDR),
        .AP_AXIMM_3_AWLEN(AP_AXIMM_3_AWLEN),
        .AP_AXIMM_3_AWSIZE(AP_AXIMM_3_AWSIZE),
        .AP_AXIMM_3_AWBURST(AP_AXIMM_3_AWBURST),
        .AP_AXIMM_3_AWLOCK(AP_AXIMM_3_AWLOCK),
        .AP_AXIMM_3_AWCACHE(AP_AXIMM_3_AWCACHE),
        .AP_AXIMM_3_AWPROT(AP_AXIMM_3_AWPROT),
        .AP_AXIMM_3_AWREGION(AP_AXIMM_3_AWREGION),
        .AP_AXIMM_3_AWQOS(AP_AXIMM_3_AWQOS),
        .AP_AXIMM_3_AWVALID(AP_AXIMM_3_AWVALID),
        .AP_AXIMM_3_AWREADY(AP_AXIMM_3_AWREADY),
        .AP_AXIMM_3_WDATA(AP_AXIMM_3_WDATA),
        .AP_AXIMM_3_WSTRB(AP_AXIMM_3_WSTRB),
        .AP_AXIMM_3_WLAST(AP_AXIMM_3_WLAST),
        .AP_AXIMM_3_WVALID(AP_AXIMM_3_WVALID),
        .AP_AXIMM_3_WREADY(AP_AXIMM_3_WREADY),
        .AP_AXIMM_3_BRESP(AP_AXIMM_3_BRESP),
        .AP_AXIMM_3_BVALID(AP_AXIMM_3_BVALID),
        .AP_AXIMM_3_BREADY(AP_AXIMM_3_BREADY),
        .AP_AXIMM_3_ARADDR(AP_AXIMM_3_ARADDR),
        .AP_AXIMM_3_ARLEN(AP_AXIMM_3_ARLEN),
        .AP_AXIMM_3_ARSIZE(AP_AXIMM_3_ARSIZE),
        .AP_AXIMM_3_ARBURST(AP_AXIMM_3_ARBURST),
        .AP_AXIMM_3_ARLOCK(AP_AXIMM_3_ARLOCK),
        .AP_AXIMM_3_ARCACHE(AP_AXIMM_3_ARCACHE),
        .AP_AXIMM_3_ARPROT(AP_AXIMM_3_ARPROT),
        .AP_AXIMM_3_ARREGION(AP_AXIMM_3_ARREGION),
        .AP_AXIMM_3_ARQOS(AP_AXIMM_3_ARQOS),
        .AP_AXIMM_3_ARVALID(AP_AXIMM_3_ARVALID),
        .AP_AXIMM_3_ARREADY(AP_AXIMM_3_ARREADY),
        .AP_AXIMM_3_RDATA(AP_AXIMM_3_RDATA),
        .AP_AXIMM_3_RRESP(AP_AXIMM_3_RRESP),
        .AP_AXIMM_3_RLAST(AP_AXIMM_3_RLAST),
        .AP_AXIMM_3_RVALID(AP_AXIMM_3_RVALID),
        .AP_AXIMM_3_RREADY(AP_AXIMM_3_RREADY),
        .M_AXIMM_3_AWADDR(M_AXIMM_3_AWADDR),
        .M_AXIMM_3_AWLEN(M_AXIMM_3_AWLEN),
        .M_AXIMM_3_AWSIZE(M_AXIMM_3_AWSIZE),
        .M_AXIMM_3_AWBURST(M_AXIMM_3_AWBURST),
        .M_AXIMM_3_AWLOCK(M_AXIMM_3_AWLOCK),
        .M_AXIMM_3_AWCACHE(M_AXIMM_3_AWCACHE),
        .M_AXIMM_3_AWPROT(M_AXIMM_3_AWPROT),
        .M_AXIMM_3_AWREGION(M_AXIMM_3_AWREGION),
        .M_AXIMM_3_AWQOS(M_AXIMM_3_AWQOS),
        .M_AXIMM_3_AWVALID(M_AXIMM_3_AWVALID),
        .M_AXIMM_3_AWREADY(M_AXIMM_3_AWREADY),
        .M_AXIMM_3_WDATA(M_AXIMM_3_WDATA),
        .M_AXIMM_3_WSTRB(M_AXIMM_3_WSTRB),
        .M_AXIMM_3_WLAST(M_AXIMM_3_WLAST),
        .M_AXIMM_3_WVALID(M_AXIMM_3_WVALID),
        .M_AXIMM_3_WREADY(M_AXIMM_3_WREADY),
        .M_AXIMM_3_BRESP(M_AXIMM_3_BRESP),
        .M_AXIMM_3_BVALID(M_AXIMM_3_BVALID),
        .M_AXIMM_3_BREADY(M_AXIMM_3_BREADY),
        .M_AXIMM_3_ARADDR(M_AXIMM_3_ARADDR),
        .M_AXIMM_3_ARLEN(M_AXIMM_3_ARLEN),
        .M_AXIMM_3_ARSIZE(M_AXIMM_3_ARSIZE),
        .M_AXIMM_3_ARBURST(M_AXIMM_3_ARBURST),
        .M_AXIMM_3_ARLOCK(M_AXIMM_3_ARLOCK),
        .M_AXIMM_3_ARCACHE(M_AXIMM_3_ARCACHE),
        .M_AXIMM_3_ARPROT(M_AXIMM_3_ARPROT),
        .M_AXIMM_3_ARREGION(M_AXIMM_3_ARREGION),
        .M_AXIMM_3_ARQOS(M_AXIMM_3_ARQOS),
        .M_AXIMM_3_ARVALID(M_AXIMM_3_ARVALID),
        .M_AXIMM_3_ARREADY(M_AXIMM_3_ARREADY),
        .M_AXIMM_3_RDATA(M_AXIMM_3_RDATA),
        .M_AXIMM_3_RRESP(M_AXIMM_3_RRESP),
        .M_AXIMM_3_RLAST(M_AXIMM_3_RLAST),
        .M_AXIMM_3_RVALID(M_AXIMM_3_RVALID),
        .M_AXIMM_3_RREADY(M_AXIMM_3_RREADY),
        .AP_AXIMM_4_AWADDR(AP_AXIMM_4_AWADDR),
        .AP_AXIMM_4_AWLEN(AP_AXIMM_4_AWLEN),
        .AP_AXIMM_4_AWSIZE(AP_AXIMM_4_AWSIZE),
        .AP_AXIMM_4_AWBURST(AP_AXIMM_4_AWBURST),
        .AP_AXIMM_4_AWLOCK(AP_AXIMM_4_AWLOCK),
        .AP_AXIMM_4_AWCACHE(AP_AXIMM_4_AWCACHE),
        .AP_AXIMM_4_AWPROT(AP_AXIMM_4_AWPROT),
        .AP_AXIMM_4_AWREGION(AP_AXIMM_4_AWREGION),
        .AP_AXIMM_4_AWQOS(AP_AXIMM_4_AWQOS),
        .AP_AXIMM_4_AWVALID(AP_AXIMM_4_AWVALID),
        .AP_AXIMM_4_AWREADY(AP_AXIMM_4_AWREADY),
        .AP_AXIMM_4_WDATA(AP_AXIMM_4_WDATA),
        .AP_AXIMM_4_WSTRB(AP_AXIMM_4_WSTRB),
        .AP_AXIMM_4_WLAST(AP_AXIMM_4_WLAST),
        .AP_AXIMM_4_WVALID(AP_AXIMM_4_WVALID),
        .AP_AXIMM_4_WREADY(AP_AXIMM_4_WREADY),
        .AP_AXIMM_4_BRESP(AP_AXIMM_4_BRESP),
        .AP_AXIMM_4_BVALID(AP_AXIMM_4_BVALID),
        .AP_AXIMM_4_BREADY(AP_AXIMM_4_BREADY),
        .AP_AXIMM_4_ARADDR(AP_AXIMM_4_ARADDR),
        .AP_AXIMM_4_ARLEN(AP_AXIMM_4_ARLEN),
        .AP_AXIMM_4_ARSIZE(AP_AXIMM_4_ARSIZE),
        .AP_AXIMM_4_ARBURST(AP_AXIMM_4_ARBURST),
        .AP_AXIMM_4_ARLOCK(AP_AXIMM_4_ARLOCK),
        .AP_AXIMM_4_ARCACHE(AP_AXIMM_4_ARCACHE),
        .AP_AXIMM_4_ARPROT(AP_AXIMM_4_ARPROT),
        .AP_AXIMM_4_ARREGION(AP_AXIMM_4_ARREGION),
        .AP_AXIMM_4_ARQOS(AP_AXIMM_4_ARQOS),
        .AP_AXIMM_4_ARVALID(AP_AXIMM_4_ARVALID),
        .AP_AXIMM_4_ARREADY(AP_AXIMM_4_ARREADY),
        .AP_AXIMM_4_RDATA(AP_AXIMM_4_RDATA),
        .AP_AXIMM_4_RRESP(AP_AXIMM_4_RRESP),
        .AP_AXIMM_4_RLAST(AP_AXIMM_4_RLAST),
        .AP_AXIMM_4_RVALID(AP_AXIMM_4_RVALID),
        .AP_AXIMM_4_RREADY(AP_AXIMM_4_RREADY),
        .M_AXIMM_4_AWADDR(M_AXIMM_4_AWADDR),
        .M_AXIMM_4_AWLEN(M_AXIMM_4_AWLEN),
        .M_AXIMM_4_AWSIZE(M_AXIMM_4_AWSIZE),
        .M_AXIMM_4_AWBURST(M_AXIMM_4_AWBURST),
        .M_AXIMM_4_AWLOCK(M_AXIMM_4_AWLOCK),
        .M_AXIMM_4_AWCACHE(M_AXIMM_4_AWCACHE),
        .M_AXIMM_4_AWPROT(M_AXIMM_4_AWPROT),
        .M_AXIMM_4_AWREGION(M_AXIMM_4_AWREGION),
        .M_AXIMM_4_AWQOS(M_AXIMM_4_AWQOS),
        .M_AXIMM_4_AWVALID(M_AXIMM_4_AWVALID),
        .M_AXIMM_4_AWREADY(M_AXIMM_4_AWREADY),
        .M_AXIMM_4_WDATA(M_AXIMM_4_WDATA),
        .M_AXIMM_4_WSTRB(M_AXIMM_4_WSTRB),
        .M_AXIMM_4_WLAST(M_AXIMM_4_WLAST),
        .M_AXIMM_4_WVALID(M_AXIMM_4_WVALID),
        .M_AXIMM_4_WREADY(M_AXIMM_4_WREADY),
        .M_AXIMM_4_BRESP(M_AXIMM_4_BRESP),
        .M_AXIMM_4_BVALID(M_AXIMM_4_BVALID),
        .M_AXIMM_4_BREADY(M_AXIMM_4_BREADY),
        .M_AXIMM_4_ARADDR(M_AXIMM_4_ARADDR),
        .M_AXIMM_4_ARLEN(M_AXIMM_4_ARLEN),
        .M_AXIMM_4_ARSIZE(M_AXIMM_4_ARSIZE),
        .M_AXIMM_4_ARBURST(M_AXIMM_4_ARBURST),
        .M_AXIMM_4_ARLOCK(M_AXIMM_4_ARLOCK),
        .M_AXIMM_4_ARCACHE(M_AXIMM_4_ARCACHE),
        .M_AXIMM_4_ARPROT(M_AXIMM_4_ARPROT),
        .M_AXIMM_4_ARREGION(M_AXIMM_4_ARREGION),
        .M_AXIMM_4_ARQOS(M_AXIMM_4_ARQOS),
        .M_AXIMM_4_ARVALID(M_AXIMM_4_ARVALID),
        .M_AXIMM_4_ARREADY(M_AXIMM_4_ARREADY),
        .M_AXIMM_4_RDATA(M_AXIMM_4_RDATA),
        .M_AXIMM_4_RRESP(M_AXIMM_4_RRESP),
        .M_AXIMM_4_RLAST(M_AXIMM_4_RLAST),
        .M_AXIMM_4_RVALID(M_AXIMM_4_RVALID),
        .M_AXIMM_4_RREADY(M_AXIMM_4_RREADY),
        .AP_AXIMM_5_AWADDR(AP_AXIMM_5_AWADDR),
        .AP_AXIMM_5_AWLEN(AP_AXIMM_5_AWLEN),
        .AP_AXIMM_5_AWSIZE(AP_AXIMM_5_AWSIZE),
        .AP_AXIMM_5_AWBURST(AP_AXIMM_5_AWBURST),
        .AP_AXIMM_5_AWLOCK(AP_AXIMM_5_AWLOCK),
        .AP_AXIMM_5_AWCACHE(AP_AXIMM_5_AWCACHE),
        .AP_AXIMM_5_AWPROT(AP_AXIMM_5_AWPROT),
        .AP_AXIMM_5_AWREGION(AP_AXIMM_5_AWREGION),
        .AP_AXIMM_5_AWQOS(AP_AXIMM_5_AWQOS),
        .AP_AXIMM_5_AWVALID(AP_AXIMM_5_AWVALID),
        .AP_AXIMM_5_AWREADY(AP_AXIMM_5_AWREADY),
        .AP_AXIMM_5_WDATA(AP_AXIMM_5_WDATA),
        .AP_AXIMM_5_WSTRB(AP_AXIMM_5_WSTRB),
        .AP_AXIMM_5_WLAST(AP_AXIMM_5_WLAST),
        .AP_AXIMM_5_WVALID(AP_AXIMM_5_WVALID),
        .AP_AXIMM_5_WREADY(AP_AXIMM_5_WREADY),
        .AP_AXIMM_5_BRESP(AP_AXIMM_5_BRESP),
        .AP_AXIMM_5_BVALID(AP_AXIMM_5_BVALID),
        .AP_AXIMM_5_BREADY(AP_AXIMM_5_BREADY),
        .AP_AXIMM_5_ARADDR(AP_AXIMM_5_ARADDR),
        .AP_AXIMM_5_ARLEN(AP_AXIMM_5_ARLEN),
        .AP_AXIMM_5_ARSIZE(AP_AXIMM_5_ARSIZE),
        .AP_AXIMM_5_ARBURST(AP_AXIMM_5_ARBURST),
        .AP_AXIMM_5_ARLOCK(AP_AXIMM_5_ARLOCK),
        .AP_AXIMM_5_ARCACHE(AP_AXIMM_5_ARCACHE),
        .AP_AXIMM_5_ARPROT(AP_AXIMM_5_ARPROT),
        .AP_AXIMM_5_ARREGION(AP_AXIMM_5_ARREGION),
        .AP_AXIMM_5_ARQOS(AP_AXIMM_5_ARQOS),
        .AP_AXIMM_5_ARVALID(AP_AXIMM_5_ARVALID),
        .AP_AXIMM_5_ARREADY(AP_AXIMM_5_ARREADY),
        .AP_AXIMM_5_RDATA(AP_AXIMM_5_RDATA),
        .AP_AXIMM_5_RRESP(AP_AXIMM_5_RRESP),
        .AP_AXIMM_5_RLAST(AP_AXIMM_5_RLAST),
        .AP_AXIMM_5_RVALID(AP_AXIMM_5_RVALID),
        .AP_AXIMM_5_RREADY(AP_AXIMM_5_RREADY),
        .M_AXIMM_5_AWADDR(M_AXIMM_5_AWADDR),
        .M_AXIMM_5_AWLEN(M_AXIMM_5_AWLEN),
        .M_AXIMM_5_AWSIZE(M_AXIMM_5_AWSIZE),
        .M_AXIMM_5_AWBURST(M_AXIMM_5_AWBURST),
        .M_AXIMM_5_AWLOCK(M_AXIMM_5_AWLOCK),
        .M_AXIMM_5_AWCACHE(M_AXIMM_5_AWCACHE),
        .M_AXIMM_5_AWPROT(M_AXIMM_5_AWPROT),
        .M_AXIMM_5_AWREGION(M_AXIMM_5_AWREGION),
        .M_AXIMM_5_AWQOS(M_AXIMM_5_AWQOS),
        .M_AXIMM_5_AWVALID(M_AXIMM_5_AWVALID),
        .M_AXIMM_5_AWREADY(M_AXIMM_5_AWREADY),
        .M_AXIMM_5_WDATA(M_AXIMM_5_WDATA),
        .M_AXIMM_5_WSTRB(M_AXIMM_5_WSTRB),
        .M_AXIMM_5_WLAST(M_AXIMM_5_WLAST),
        .M_AXIMM_5_WVALID(M_AXIMM_5_WVALID),
        .M_AXIMM_5_WREADY(M_AXIMM_5_WREADY),
        .M_AXIMM_5_BRESP(M_AXIMM_5_BRESP),
        .M_AXIMM_5_BVALID(M_AXIMM_5_BVALID),
        .M_AXIMM_5_BREADY(M_AXIMM_5_BREADY),
        .M_AXIMM_5_ARADDR(M_AXIMM_5_ARADDR),
        .M_AXIMM_5_ARLEN(M_AXIMM_5_ARLEN),
        .M_AXIMM_5_ARSIZE(M_AXIMM_5_ARSIZE),
        .M_AXIMM_5_ARBURST(M_AXIMM_5_ARBURST),
        .M_AXIMM_5_ARLOCK(M_AXIMM_5_ARLOCK),
        .M_AXIMM_5_ARCACHE(M_AXIMM_5_ARCACHE),
        .M_AXIMM_5_ARPROT(M_AXIMM_5_ARPROT),
        .M_AXIMM_5_ARREGION(M_AXIMM_5_ARREGION),
        .M_AXIMM_5_ARQOS(M_AXIMM_5_ARQOS),
        .M_AXIMM_5_ARVALID(M_AXIMM_5_ARVALID),
        .M_AXIMM_5_ARREADY(M_AXIMM_5_ARREADY),
        .M_AXIMM_5_RDATA(M_AXIMM_5_RDATA),
        .M_AXIMM_5_RRESP(M_AXIMM_5_RRESP),
        .M_AXIMM_5_RLAST(M_AXIMM_5_RLAST),
        .M_AXIMM_5_RVALID(M_AXIMM_5_RVALID),
        .M_AXIMM_5_RREADY(M_AXIMM_5_RREADY),
        .AP_AXIMM_6_AWADDR(AP_AXIMM_6_AWADDR),
        .AP_AXIMM_6_AWLEN(AP_AXIMM_6_AWLEN),
        .AP_AXIMM_6_AWSIZE(AP_AXIMM_6_AWSIZE),
        .AP_AXIMM_6_AWBURST(AP_AXIMM_6_AWBURST),
        .AP_AXIMM_6_AWLOCK(AP_AXIMM_6_AWLOCK),
        .AP_AXIMM_6_AWCACHE(AP_AXIMM_6_AWCACHE),
        .AP_AXIMM_6_AWPROT(AP_AXIMM_6_AWPROT),
        .AP_AXIMM_6_AWREGION(AP_AXIMM_6_AWREGION),
        .AP_AXIMM_6_AWQOS(AP_AXIMM_6_AWQOS),
        .AP_AXIMM_6_AWVALID(AP_AXIMM_6_AWVALID),
        .AP_AXIMM_6_AWREADY(AP_AXIMM_6_AWREADY),
        .AP_AXIMM_6_WDATA(AP_AXIMM_6_WDATA),
        .AP_AXIMM_6_WSTRB(AP_AXIMM_6_WSTRB),
        .AP_AXIMM_6_WLAST(AP_AXIMM_6_WLAST),
        .AP_AXIMM_6_WVALID(AP_AXIMM_6_WVALID),
        .AP_AXIMM_6_WREADY(AP_AXIMM_6_WREADY),
        .AP_AXIMM_6_BRESP(AP_AXIMM_6_BRESP),
        .AP_AXIMM_6_BVALID(AP_AXIMM_6_BVALID),
        .AP_AXIMM_6_BREADY(AP_AXIMM_6_BREADY),
        .AP_AXIMM_6_ARADDR(AP_AXIMM_6_ARADDR),
        .AP_AXIMM_6_ARLEN(AP_AXIMM_6_ARLEN),
        .AP_AXIMM_6_ARSIZE(AP_AXIMM_6_ARSIZE),
        .AP_AXIMM_6_ARBURST(AP_AXIMM_6_ARBURST),
        .AP_AXIMM_6_ARLOCK(AP_AXIMM_6_ARLOCK),
        .AP_AXIMM_6_ARCACHE(AP_AXIMM_6_ARCACHE),
        .AP_AXIMM_6_ARPROT(AP_AXIMM_6_ARPROT),
        .AP_AXIMM_6_ARREGION(AP_AXIMM_6_ARREGION),
        .AP_AXIMM_6_ARQOS(AP_AXIMM_6_ARQOS),
        .AP_AXIMM_6_ARVALID(AP_AXIMM_6_ARVALID),
        .AP_AXIMM_6_ARREADY(AP_AXIMM_6_ARREADY),
        .AP_AXIMM_6_RDATA(AP_AXIMM_6_RDATA),
        .AP_AXIMM_6_RRESP(AP_AXIMM_6_RRESP),
        .AP_AXIMM_6_RLAST(AP_AXIMM_6_RLAST),
        .AP_AXIMM_6_RVALID(AP_AXIMM_6_RVALID),
        .AP_AXIMM_6_RREADY(AP_AXIMM_6_RREADY),
        .M_AXIMM_6_AWADDR(M_AXIMM_6_AWADDR),
        .M_AXIMM_6_AWLEN(M_AXIMM_6_AWLEN),
        .M_AXIMM_6_AWSIZE(M_AXIMM_6_AWSIZE),
        .M_AXIMM_6_AWBURST(M_AXIMM_6_AWBURST),
        .M_AXIMM_6_AWLOCK(M_AXIMM_6_AWLOCK),
        .M_AXIMM_6_AWCACHE(M_AXIMM_6_AWCACHE),
        .M_AXIMM_6_AWPROT(M_AXIMM_6_AWPROT),
        .M_AXIMM_6_AWREGION(M_AXIMM_6_AWREGION),
        .M_AXIMM_6_AWQOS(M_AXIMM_6_AWQOS),
        .M_AXIMM_6_AWVALID(M_AXIMM_6_AWVALID),
        .M_AXIMM_6_AWREADY(M_AXIMM_6_AWREADY),
        .M_AXIMM_6_WDATA(M_AXIMM_6_WDATA),
        .M_AXIMM_6_WSTRB(M_AXIMM_6_WSTRB),
        .M_AXIMM_6_WLAST(M_AXIMM_6_WLAST),
        .M_AXIMM_6_WVALID(M_AXIMM_6_WVALID),
        .M_AXIMM_6_WREADY(M_AXIMM_6_WREADY),
        .M_AXIMM_6_BRESP(M_AXIMM_6_BRESP),
        .M_AXIMM_6_BVALID(M_AXIMM_6_BVALID),
        .M_AXIMM_6_BREADY(M_AXIMM_6_BREADY),
        .M_AXIMM_6_ARADDR(M_AXIMM_6_ARADDR),
        .M_AXIMM_6_ARLEN(M_AXIMM_6_ARLEN),
        .M_AXIMM_6_ARSIZE(M_AXIMM_6_ARSIZE),
        .M_AXIMM_6_ARBURST(M_AXIMM_6_ARBURST),
        .M_AXIMM_6_ARLOCK(M_AXIMM_6_ARLOCK),
        .M_AXIMM_6_ARCACHE(M_AXIMM_6_ARCACHE),
        .M_AXIMM_6_ARPROT(M_AXIMM_6_ARPROT),
        .M_AXIMM_6_ARREGION(M_AXIMM_6_ARREGION),
        .M_AXIMM_6_ARQOS(M_AXIMM_6_ARQOS),
        .M_AXIMM_6_ARVALID(M_AXIMM_6_ARVALID),
        .M_AXIMM_6_ARREADY(M_AXIMM_6_ARREADY),
        .M_AXIMM_6_RDATA(M_AXIMM_6_RDATA),
        .M_AXIMM_6_RRESP(M_AXIMM_6_RRESP),
        .M_AXIMM_6_RLAST(M_AXIMM_6_RLAST),
        .M_AXIMM_6_RVALID(M_AXIMM_6_RVALID),
        .M_AXIMM_6_RREADY(M_AXIMM_6_RREADY),
        .AP_AXIMM_7_AWADDR(AP_AXIMM_7_AWADDR),
        .AP_AXIMM_7_AWLEN(AP_AXIMM_7_AWLEN),
        .AP_AXIMM_7_AWSIZE(AP_AXIMM_7_AWSIZE),
        .AP_AXIMM_7_AWBURST(AP_AXIMM_7_AWBURST),
        .AP_AXIMM_7_AWLOCK(AP_AXIMM_7_AWLOCK),
        .AP_AXIMM_7_AWCACHE(AP_AXIMM_7_AWCACHE),
        .AP_AXIMM_7_AWPROT(AP_AXIMM_7_AWPROT),
        .AP_AXIMM_7_AWREGION(AP_AXIMM_7_AWREGION),
        .AP_AXIMM_7_AWQOS(AP_AXIMM_7_AWQOS),
        .AP_AXIMM_7_AWVALID(AP_AXIMM_7_AWVALID),
        .AP_AXIMM_7_AWREADY(AP_AXIMM_7_AWREADY),
        .AP_AXIMM_7_WDATA(AP_AXIMM_7_WDATA),
        .AP_AXIMM_7_WSTRB(AP_AXIMM_7_WSTRB),
        .AP_AXIMM_7_WLAST(AP_AXIMM_7_WLAST),
        .AP_AXIMM_7_WVALID(AP_AXIMM_7_WVALID),
        .AP_AXIMM_7_WREADY(AP_AXIMM_7_WREADY),
        .AP_AXIMM_7_BRESP(AP_AXIMM_7_BRESP),
        .AP_AXIMM_7_BVALID(AP_AXIMM_7_BVALID),
        .AP_AXIMM_7_BREADY(AP_AXIMM_7_BREADY),
        .AP_AXIMM_7_ARADDR(AP_AXIMM_7_ARADDR),
        .AP_AXIMM_7_ARLEN(AP_AXIMM_7_ARLEN),
        .AP_AXIMM_7_ARSIZE(AP_AXIMM_7_ARSIZE),
        .AP_AXIMM_7_ARBURST(AP_AXIMM_7_ARBURST),
        .AP_AXIMM_7_ARLOCK(AP_AXIMM_7_ARLOCK),
        .AP_AXIMM_7_ARCACHE(AP_AXIMM_7_ARCACHE),
        .AP_AXIMM_7_ARPROT(AP_AXIMM_7_ARPROT),
        .AP_AXIMM_7_ARREGION(AP_AXIMM_7_ARREGION),
        .AP_AXIMM_7_ARQOS(AP_AXIMM_7_ARQOS),
        .AP_AXIMM_7_ARVALID(AP_AXIMM_7_ARVALID),
        .AP_AXIMM_7_ARREADY(AP_AXIMM_7_ARREADY),
        .AP_AXIMM_7_RDATA(AP_AXIMM_7_RDATA),
        .AP_AXIMM_7_RRESP(AP_AXIMM_7_RRESP),
        .AP_AXIMM_7_RLAST(AP_AXIMM_7_RLAST),
        .AP_AXIMM_7_RVALID(AP_AXIMM_7_RVALID),
        .AP_AXIMM_7_RREADY(AP_AXIMM_7_RREADY),
        .M_AXIMM_7_AWADDR(M_AXIMM_7_AWADDR),
        .M_AXIMM_7_AWLEN(M_AXIMM_7_AWLEN),
        .M_AXIMM_7_AWSIZE(M_AXIMM_7_AWSIZE),
        .M_AXIMM_7_AWBURST(M_AXIMM_7_AWBURST),
        .M_AXIMM_7_AWLOCK(M_AXIMM_7_AWLOCK),
        .M_AXIMM_7_AWCACHE(M_AXIMM_7_AWCACHE),
        .M_AXIMM_7_AWPROT(M_AXIMM_7_AWPROT),
        .M_AXIMM_7_AWREGION(M_AXIMM_7_AWREGION),
        .M_AXIMM_7_AWQOS(M_AXIMM_7_AWQOS),
        .M_AXIMM_7_AWVALID(M_AXIMM_7_AWVALID),
        .M_AXIMM_7_AWREADY(M_AXIMM_7_AWREADY),
        .M_AXIMM_7_WDATA(M_AXIMM_7_WDATA),
        .M_AXIMM_7_WSTRB(M_AXIMM_7_WSTRB),
        .M_AXIMM_7_WLAST(M_AXIMM_7_WLAST),
        .M_AXIMM_7_WVALID(M_AXIMM_7_WVALID),
        .M_AXIMM_7_WREADY(M_AXIMM_7_WREADY),
        .M_AXIMM_7_BRESP(M_AXIMM_7_BRESP),
        .M_AXIMM_7_BVALID(M_AXIMM_7_BVALID),
        .M_AXIMM_7_BREADY(M_AXIMM_7_BREADY),
        .M_AXIMM_7_ARADDR(M_AXIMM_7_ARADDR),
        .M_AXIMM_7_ARLEN(M_AXIMM_7_ARLEN),
        .M_AXIMM_7_ARSIZE(M_AXIMM_7_ARSIZE),
        .M_AXIMM_7_ARBURST(M_AXIMM_7_ARBURST),
        .M_AXIMM_7_ARLOCK(M_AXIMM_7_ARLOCK),
        .M_AXIMM_7_ARCACHE(M_AXIMM_7_ARCACHE),
        .M_AXIMM_7_ARPROT(M_AXIMM_7_ARPROT),
        .M_AXIMM_7_ARREGION(M_AXIMM_7_ARREGION),
        .M_AXIMM_7_ARQOS(M_AXIMM_7_ARQOS),
        .M_AXIMM_7_ARVALID(M_AXIMM_7_ARVALID),
        .M_AXIMM_7_ARREADY(M_AXIMM_7_ARREADY),
        .M_AXIMM_7_RDATA(M_AXIMM_7_RDATA),
        .M_AXIMM_7_RRESP(M_AXIMM_7_RRESP),
        .M_AXIMM_7_RLAST(M_AXIMM_7_RLAST),
        .M_AXIMM_7_RVALID(M_AXIMM_7_RVALID),
        .M_AXIMM_7_RREADY(M_AXIMM_7_RREADY),
        .AP_AXIMM_8_AWADDR(AP_AXIMM_8_AWADDR),
        .AP_AXIMM_8_AWLEN(AP_AXIMM_8_AWLEN),
        .AP_AXIMM_8_AWSIZE(AP_AXIMM_8_AWSIZE),
        .AP_AXIMM_8_AWBURST(AP_AXIMM_8_AWBURST),
        .AP_AXIMM_8_AWLOCK(AP_AXIMM_8_AWLOCK),
        .AP_AXIMM_8_AWCACHE(AP_AXIMM_8_AWCACHE),
        .AP_AXIMM_8_AWPROT(AP_AXIMM_8_AWPROT),
        .AP_AXIMM_8_AWREGION(AP_AXIMM_8_AWREGION),
        .AP_AXIMM_8_AWQOS(AP_AXIMM_8_AWQOS),
        .AP_AXIMM_8_AWVALID(AP_AXIMM_8_AWVALID),
        .AP_AXIMM_8_AWREADY(AP_AXIMM_8_AWREADY),
        .AP_AXIMM_8_WDATA(AP_AXIMM_8_WDATA),
        .AP_AXIMM_8_WSTRB(AP_AXIMM_8_WSTRB),
        .AP_AXIMM_8_WLAST(AP_AXIMM_8_WLAST),
        .AP_AXIMM_8_WVALID(AP_AXIMM_8_WVALID),
        .AP_AXIMM_8_WREADY(AP_AXIMM_8_WREADY),
        .AP_AXIMM_8_BRESP(AP_AXIMM_8_BRESP),
        .AP_AXIMM_8_BVALID(AP_AXIMM_8_BVALID),
        .AP_AXIMM_8_BREADY(AP_AXIMM_8_BREADY),
        .AP_AXIMM_8_ARADDR(AP_AXIMM_8_ARADDR),
        .AP_AXIMM_8_ARLEN(AP_AXIMM_8_ARLEN),
        .AP_AXIMM_8_ARSIZE(AP_AXIMM_8_ARSIZE),
        .AP_AXIMM_8_ARBURST(AP_AXIMM_8_ARBURST),
        .AP_AXIMM_8_ARLOCK(AP_AXIMM_8_ARLOCK),
        .AP_AXIMM_8_ARCACHE(AP_AXIMM_8_ARCACHE),
        .AP_AXIMM_8_ARPROT(AP_AXIMM_8_ARPROT),
        .AP_AXIMM_8_ARREGION(AP_AXIMM_8_ARREGION),
        .AP_AXIMM_8_ARQOS(AP_AXIMM_8_ARQOS),
        .AP_AXIMM_8_ARVALID(AP_AXIMM_8_ARVALID),
        .AP_AXIMM_8_ARREADY(AP_AXIMM_8_ARREADY),
        .AP_AXIMM_8_RDATA(AP_AXIMM_8_RDATA),
        .AP_AXIMM_8_RRESP(AP_AXIMM_8_RRESP),
        .AP_AXIMM_8_RLAST(AP_AXIMM_8_RLAST),
        .AP_AXIMM_8_RVALID(AP_AXIMM_8_RVALID),
        .AP_AXIMM_8_RREADY(AP_AXIMM_8_RREADY),
        .M_AXIMM_8_AWADDR(M_AXIMM_8_AWADDR),
        .M_AXIMM_8_AWLEN(M_AXIMM_8_AWLEN),
        .M_AXIMM_8_AWSIZE(M_AXIMM_8_AWSIZE),
        .M_AXIMM_8_AWBURST(M_AXIMM_8_AWBURST),
        .M_AXIMM_8_AWLOCK(M_AXIMM_8_AWLOCK),
        .M_AXIMM_8_AWCACHE(M_AXIMM_8_AWCACHE),
        .M_AXIMM_8_AWPROT(M_AXIMM_8_AWPROT),
        .M_AXIMM_8_AWREGION(M_AXIMM_8_AWREGION),
        .M_AXIMM_8_AWQOS(M_AXIMM_8_AWQOS),
        .M_AXIMM_8_AWVALID(M_AXIMM_8_AWVALID),
        .M_AXIMM_8_AWREADY(M_AXIMM_8_AWREADY),
        .M_AXIMM_8_WDATA(M_AXIMM_8_WDATA),
        .M_AXIMM_8_WSTRB(M_AXIMM_8_WSTRB),
        .M_AXIMM_8_WLAST(M_AXIMM_8_WLAST),
        .M_AXIMM_8_WVALID(M_AXIMM_8_WVALID),
        .M_AXIMM_8_WREADY(M_AXIMM_8_WREADY),
        .M_AXIMM_8_BRESP(M_AXIMM_8_BRESP),
        .M_AXIMM_8_BVALID(M_AXIMM_8_BVALID),
        .M_AXIMM_8_BREADY(M_AXIMM_8_BREADY),
        .M_AXIMM_8_ARADDR(M_AXIMM_8_ARADDR),
        .M_AXIMM_8_ARLEN(M_AXIMM_8_ARLEN),
        .M_AXIMM_8_ARSIZE(M_AXIMM_8_ARSIZE),
        .M_AXIMM_8_ARBURST(M_AXIMM_8_ARBURST),
        .M_AXIMM_8_ARLOCK(M_AXIMM_8_ARLOCK),
        .M_AXIMM_8_ARCACHE(M_AXIMM_8_ARCACHE),
        .M_AXIMM_8_ARPROT(M_AXIMM_8_ARPROT),
        .M_AXIMM_8_ARREGION(M_AXIMM_8_ARREGION),
        .M_AXIMM_8_ARQOS(M_AXIMM_8_ARQOS),
        .M_AXIMM_8_ARVALID(M_AXIMM_8_ARVALID),
        .M_AXIMM_8_ARREADY(M_AXIMM_8_ARREADY),
        .M_AXIMM_8_RDATA(M_AXIMM_8_RDATA),
        .M_AXIMM_8_RRESP(M_AXIMM_8_RRESP),
        .M_AXIMM_8_RLAST(M_AXIMM_8_RLAST),
        .M_AXIMM_8_RVALID(M_AXIMM_8_RVALID),
        .M_AXIMM_8_RREADY(M_AXIMM_8_RREADY),
        .AP_AXIMM_9_AWADDR(AP_AXIMM_9_AWADDR),
        .AP_AXIMM_9_AWLEN(AP_AXIMM_9_AWLEN),
        .AP_AXIMM_9_AWSIZE(AP_AXIMM_9_AWSIZE),
        .AP_AXIMM_9_AWBURST(AP_AXIMM_9_AWBURST),
        .AP_AXIMM_9_AWLOCK(AP_AXIMM_9_AWLOCK),
        .AP_AXIMM_9_AWCACHE(AP_AXIMM_9_AWCACHE),
        .AP_AXIMM_9_AWPROT(AP_AXIMM_9_AWPROT),
        .AP_AXIMM_9_AWREGION(AP_AXIMM_9_AWREGION),
        .AP_AXIMM_9_AWQOS(AP_AXIMM_9_AWQOS),
        .AP_AXIMM_9_AWVALID(AP_AXIMM_9_AWVALID),
        .AP_AXIMM_9_AWREADY(AP_AXIMM_9_AWREADY),
        .AP_AXIMM_9_WDATA(AP_AXIMM_9_WDATA),
        .AP_AXIMM_9_WSTRB(AP_AXIMM_9_WSTRB),
        .AP_AXIMM_9_WLAST(AP_AXIMM_9_WLAST),
        .AP_AXIMM_9_WVALID(AP_AXIMM_9_WVALID),
        .AP_AXIMM_9_WREADY(AP_AXIMM_9_WREADY),
        .AP_AXIMM_9_BRESP(AP_AXIMM_9_BRESP),
        .AP_AXIMM_9_BVALID(AP_AXIMM_9_BVALID),
        .AP_AXIMM_9_BREADY(AP_AXIMM_9_BREADY),
        .AP_AXIMM_9_ARADDR(AP_AXIMM_9_ARADDR),
        .AP_AXIMM_9_ARLEN(AP_AXIMM_9_ARLEN),
        .AP_AXIMM_9_ARSIZE(AP_AXIMM_9_ARSIZE),
        .AP_AXIMM_9_ARBURST(AP_AXIMM_9_ARBURST),
        .AP_AXIMM_9_ARLOCK(AP_AXIMM_9_ARLOCK),
        .AP_AXIMM_9_ARCACHE(AP_AXIMM_9_ARCACHE),
        .AP_AXIMM_9_ARPROT(AP_AXIMM_9_ARPROT),
        .AP_AXIMM_9_ARREGION(AP_AXIMM_9_ARREGION),
        .AP_AXIMM_9_ARQOS(AP_AXIMM_9_ARQOS),
        .AP_AXIMM_9_ARVALID(AP_AXIMM_9_ARVALID),
        .AP_AXIMM_9_ARREADY(AP_AXIMM_9_ARREADY),
        .AP_AXIMM_9_RDATA(AP_AXIMM_9_RDATA),
        .AP_AXIMM_9_RRESP(AP_AXIMM_9_RRESP),
        .AP_AXIMM_9_RLAST(AP_AXIMM_9_RLAST),
        .AP_AXIMM_9_RVALID(AP_AXIMM_9_RVALID),
        .AP_AXIMM_9_RREADY(AP_AXIMM_9_RREADY),
        .M_AXIMM_9_AWADDR(M_AXIMM_9_AWADDR),
        .M_AXIMM_9_AWLEN(M_AXIMM_9_AWLEN),
        .M_AXIMM_9_AWSIZE(M_AXIMM_9_AWSIZE),
        .M_AXIMM_9_AWBURST(M_AXIMM_9_AWBURST),
        .M_AXIMM_9_AWLOCK(M_AXIMM_9_AWLOCK),
        .M_AXIMM_9_AWCACHE(M_AXIMM_9_AWCACHE),
        .M_AXIMM_9_AWPROT(M_AXIMM_9_AWPROT),
        .M_AXIMM_9_AWREGION(M_AXIMM_9_AWREGION),
        .M_AXIMM_9_AWQOS(M_AXIMM_9_AWQOS),
        .M_AXIMM_9_AWVALID(M_AXIMM_9_AWVALID),
        .M_AXIMM_9_AWREADY(M_AXIMM_9_AWREADY),
        .M_AXIMM_9_WDATA(M_AXIMM_9_WDATA),
        .M_AXIMM_9_WSTRB(M_AXIMM_9_WSTRB),
        .M_AXIMM_9_WLAST(M_AXIMM_9_WLAST),
        .M_AXIMM_9_WVALID(M_AXIMM_9_WVALID),
        .M_AXIMM_9_WREADY(M_AXIMM_9_WREADY),
        .M_AXIMM_9_BRESP(M_AXIMM_9_BRESP),
        .M_AXIMM_9_BVALID(M_AXIMM_9_BVALID),
        .M_AXIMM_9_BREADY(M_AXIMM_9_BREADY),
        .M_AXIMM_9_ARADDR(M_AXIMM_9_ARADDR),
        .M_AXIMM_9_ARLEN(M_AXIMM_9_ARLEN),
        .M_AXIMM_9_ARSIZE(M_AXIMM_9_ARSIZE),
        .M_AXIMM_9_ARBURST(M_AXIMM_9_ARBURST),
        .M_AXIMM_9_ARLOCK(M_AXIMM_9_ARLOCK),
        .M_AXIMM_9_ARCACHE(M_AXIMM_9_ARCACHE),
        .M_AXIMM_9_ARPROT(M_AXIMM_9_ARPROT),
        .M_AXIMM_9_ARREGION(M_AXIMM_9_ARREGION),
        .M_AXIMM_9_ARQOS(M_AXIMM_9_ARQOS),
        .M_AXIMM_9_ARVALID(M_AXIMM_9_ARVALID),
        .M_AXIMM_9_ARREADY(M_AXIMM_9_ARREADY),
        .M_AXIMM_9_RDATA(M_AXIMM_9_RDATA),
        .M_AXIMM_9_RRESP(M_AXIMM_9_RRESP),
        .M_AXIMM_9_RLAST(M_AXIMM_9_RLAST),
        .M_AXIMM_9_RVALID(M_AXIMM_9_RVALID),
        .M_AXIMM_9_RREADY(M_AXIMM_9_RREADY),
        .AP_AXIMM_10_AWADDR(AP_AXIMM_10_AWADDR),
        .AP_AXIMM_10_AWLEN(AP_AXIMM_10_AWLEN),
        .AP_AXIMM_10_AWSIZE(AP_AXIMM_10_AWSIZE),
        .AP_AXIMM_10_AWBURST(AP_AXIMM_10_AWBURST),
        .AP_AXIMM_10_AWLOCK(AP_AXIMM_10_AWLOCK),
        .AP_AXIMM_10_AWCACHE(AP_AXIMM_10_AWCACHE),
        .AP_AXIMM_10_AWPROT(AP_AXIMM_10_AWPROT),
        .AP_AXIMM_10_AWREGION(AP_AXIMM_10_AWREGION),
        .AP_AXIMM_10_AWQOS(AP_AXIMM_10_AWQOS),
        .AP_AXIMM_10_AWVALID(AP_AXIMM_10_AWVALID),
        .AP_AXIMM_10_AWREADY(AP_AXIMM_10_AWREADY),
        .AP_AXIMM_10_WDATA(AP_AXIMM_10_WDATA),
        .AP_AXIMM_10_WSTRB(AP_AXIMM_10_WSTRB),
        .AP_AXIMM_10_WLAST(AP_AXIMM_10_WLAST),
        .AP_AXIMM_10_WVALID(AP_AXIMM_10_WVALID),
        .AP_AXIMM_10_WREADY(AP_AXIMM_10_WREADY),
        .AP_AXIMM_10_BRESP(AP_AXIMM_10_BRESP),
        .AP_AXIMM_10_BVALID(AP_AXIMM_10_BVALID),
        .AP_AXIMM_10_BREADY(AP_AXIMM_10_BREADY),
        .AP_AXIMM_10_ARADDR(AP_AXIMM_10_ARADDR),
        .AP_AXIMM_10_ARLEN(AP_AXIMM_10_ARLEN),
        .AP_AXIMM_10_ARSIZE(AP_AXIMM_10_ARSIZE),
        .AP_AXIMM_10_ARBURST(AP_AXIMM_10_ARBURST),
        .AP_AXIMM_10_ARLOCK(AP_AXIMM_10_ARLOCK),
        .AP_AXIMM_10_ARCACHE(AP_AXIMM_10_ARCACHE),
        .AP_AXIMM_10_ARPROT(AP_AXIMM_10_ARPROT),
        .AP_AXIMM_10_ARREGION(AP_AXIMM_10_ARREGION),
        .AP_AXIMM_10_ARQOS(AP_AXIMM_10_ARQOS),
        .AP_AXIMM_10_ARVALID(AP_AXIMM_10_ARVALID),
        .AP_AXIMM_10_ARREADY(AP_AXIMM_10_ARREADY),
        .AP_AXIMM_10_RDATA(AP_AXIMM_10_RDATA),
        .AP_AXIMM_10_RRESP(AP_AXIMM_10_RRESP),
        .AP_AXIMM_10_RLAST(AP_AXIMM_10_RLAST),
        .AP_AXIMM_10_RVALID(AP_AXIMM_10_RVALID),
        .AP_AXIMM_10_RREADY(AP_AXIMM_10_RREADY),
        .M_AXIMM_10_AWADDR(M_AXIMM_10_AWADDR),
        .M_AXIMM_10_AWLEN(M_AXIMM_10_AWLEN),
        .M_AXIMM_10_AWSIZE(M_AXIMM_10_AWSIZE),
        .M_AXIMM_10_AWBURST(M_AXIMM_10_AWBURST),
        .M_AXIMM_10_AWLOCK(M_AXIMM_10_AWLOCK),
        .M_AXIMM_10_AWCACHE(M_AXIMM_10_AWCACHE),
        .M_AXIMM_10_AWPROT(M_AXIMM_10_AWPROT),
        .M_AXIMM_10_AWREGION(M_AXIMM_10_AWREGION),
        .M_AXIMM_10_AWQOS(M_AXIMM_10_AWQOS),
        .M_AXIMM_10_AWVALID(M_AXIMM_10_AWVALID),
        .M_AXIMM_10_AWREADY(M_AXIMM_10_AWREADY),
        .M_AXIMM_10_WDATA(M_AXIMM_10_WDATA),
        .M_AXIMM_10_WSTRB(M_AXIMM_10_WSTRB),
        .M_AXIMM_10_WLAST(M_AXIMM_10_WLAST),
        .M_AXIMM_10_WVALID(M_AXIMM_10_WVALID),
        .M_AXIMM_10_WREADY(M_AXIMM_10_WREADY),
        .M_AXIMM_10_BRESP(M_AXIMM_10_BRESP),
        .M_AXIMM_10_BVALID(M_AXIMM_10_BVALID),
        .M_AXIMM_10_BREADY(M_AXIMM_10_BREADY),
        .M_AXIMM_10_ARADDR(M_AXIMM_10_ARADDR),
        .M_AXIMM_10_ARLEN(M_AXIMM_10_ARLEN),
        .M_AXIMM_10_ARSIZE(M_AXIMM_10_ARSIZE),
        .M_AXIMM_10_ARBURST(M_AXIMM_10_ARBURST),
        .M_AXIMM_10_ARLOCK(M_AXIMM_10_ARLOCK),
        .M_AXIMM_10_ARCACHE(M_AXIMM_10_ARCACHE),
        .M_AXIMM_10_ARPROT(M_AXIMM_10_ARPROT),
        .M_AXIMM_10_ARREGION(M_AXIMM_10_ARREGION),
        .M_AXIMM_10_ARQOS(M_AXIMM_10_ARQOS),
        .M_AXIMM_10_ARVALID(M_AXIMM_10_ARVALID),
        .M_AXIMM_10_ARREADY(M_AXIMM_10_ARREADY),
        .M_AXIMM_10_RDATA(M_AXIMM_10_RDATA),
        .M_AXIMM_10_RRESP(M_AXIMM_10_RRESP),
        .M_AXIMM_10_RLAST(M_AXIMM_10_RLAST),
        .M_AXIMM_10_RVALID(M_AXIMM_10_RVALID),
        .M_AXIMM_10_RREADY(M_AXIMM_10_RREADY),
        .AP_AXIMM_11_AWADDR(AP_AXIMM_11_AWADDR),
        .AP_AXIMM_11_AWLEN(AP_AXIMM_11_AWLEN),
        .AP_AXIMM_11_AWSIZE(AP_AXIMM_11_AWSIZE),
        .AP_AXIMM_11_AWBURST(AP_AXIMM_11_AWBURST),
        .AP_AXIMM_11_AWLOCK(AP_AXIMM_11_AWLOCK),
        .AP_AXIMM_11_AWCACHE(AP_AXIMM_11_AWCACHE),
        .AP_AXIMM_11_AWPROT(AP_AXIMM_11_AWPROT),
        .AP_AXIMM_11_AWREGION(AP_AXIMM_11_AWREGION),
        .AP_AXIMM_11_AWQOS(AP_AXIMM_11_AWQOS),
        .AP_AXIMM_11_AWVALID(AP_AXIMM_11_AWVALID),
        .AP_AXIMM_11_AWREADY(AP_AXIMM_11_AWREADY),
        .AP_AXIMM_11_WDATA(AP_AXIMM_11_WDATA),
        .AP_AXIMM_11_WSTRB(AP_AXIMM_11_WSTRB),
        .AP_AXIMM_11_WLAST(AP_AXIMM_11_WLAST),
        .AP_AXIMM_11_WVALID(AP_AXIMM_11_WVALID),
        .AP_AXIMM_11_WREADY(AP_AXIMM_11_WREADY),
        .AP_AXIMM_11_BRESP(AP_AXIMM_11_BRESP),
        .AP_AXIMM_11_BVALID(AP_AXIMM_11_BVALID),
        .AP_AXIMM_11_BREADY(AP_AXIMM_11_BREADY),
        .AP_AXIMM_11_ARADDR(AP_AXIMM_11_ARADDR),
        .AP_AXIMM_11_ARLEN(AP_AXIMM_11_ARLEN),
        .AP_AXIMM_11_ARSIZE(AP_AXIMM_11_ARSIZE),
        .AP_AXIMM_11_ARBURST(AP_AXIMM_11_ARBURST),
        .AP_AXIMM_11_ARLOCK(AP_AXIMM_11_ARLOCK),
        .AP_AXIMM_11_ARCACHE(AP_AXIMM_11_ARCACHE),
        .AP_AXIMM_11_ARPROT(AP_AXIMM_11_ARPROT),
        .AP_AXIMM_11_ARREGION(AP_AXIMM_11_ARREGION),
        .AP_AXIMM_11_ARQOS(AP_AXIMM_11_ARQOS),
        .AP_AXIMM_11_ARVALID(AP_AXIMM_11_ARVALID),
        .AP_AXIMM_11_ARREADY(AP_AXIMM_11_ARREADY),
        .AP_AXIMM_11_RDATA(AP_AXIMM_11_RDATA),
        .AP_AXIMM_11_RRESP(AP_AXIMM_11_RRESP),
        .AP_AXIMM_11_RLAST(AP_AXIMM_11_RLAST),
        .AP_AXIMM_11_RVALID(AP_AXIMM_11_RVALID),
        .AP_AXIMM_11_RREADY(AP_AXIMM_11_RREADY),
        .M_AXIMM_11_AWADDR(M_AXIMM_11_AWADDR),
        .M_AXIMM_11_AWLEN(M_AXIMM_11_AWLEN),
        .M_AXIMM_11_AWSIZE(M_AXIMM_11_AWSIZE),
        .M_AXIMM_11_AWBURST(M_AXIMM_11_AWBURST),
        .M_AXIMM_11_AWLOCK(M_AXIMM_11_AWLOCK),
        .M_AXIMM_11_AWCACHE(M_AXIMM_11_AWCACHE),
        .M_AXIMM_11_AWPROT(M_AXIMM_11_AWPROT),
        .M_AXIMM_11_AWREGION(M_AXIMM_11_AWREGION),
        .M_AXIMM_11_AWQOS(M_AXIMM_11_AWQOS),
        .M_AXIMM_11_AWVALID(M_AXIMM_11_AWVALID),
        .M_AXIMM_11_AWREADY(M_AXIMM_11_AWREADY),
        .M_AXIMM_11_WDATA(M_AXIMM_11_WDATA),
        .M_AXIMM_11_WSTRB(M_AXIMM_11_WSTRB),
        .M_AXIMM_11_WLAST(M_AXIMM_11_WLAST),
        .M_AXIMM_11_WVALID(M_AXIMM_11_WVALID),
        .M_AXIMM_11_WREADY(M_AXIMM_11_WREADY),
        .M_AXIMM_11_BRESP(M_AXIMM_11_BRESP),
        .M_AXIMM_11_BVALID(M_AXIMM_11_BVALID),
        .M_AXIMM_11_BREADY(M_AXIMM_11_BREADY),
        .M_AXIMM_11_ARADDR(M_AXIMM_11_ARADDR),
        .M_AXIMM_11_ARLEN(M_AXIMM_11_ARLEN),
        .M_AXIMM_11_ARSIZE(M_AXIMM_11_ARSIZE),
        .M_AXIMM_11_ARBURST(M_AXIMM_11_ARBURST),
        .M_AXIMM_11_ARLOCK(M_AXIMM_11_ARLOCK),
        .M_AXIMM_11_ARCACHE(M_AXIMM_11_ARCACHE),
        .M_AXIMM_11_ARPROT(M_AXIMM_11_ARPROT),
        .M_AXIMM_11_ARREGION(M_AXIMM_11_ARREGION),
        .M_AXIMM_11_ARQOS(M_AXIMM_11_ARQOS),
        .M_AXIMM_11_ARVALID(M_AXIMM_11_ARVALID),
        .M_AXIMM_11_ARREADY(M_AXIMM_11_ARREADY),
        .M_AXIMM_11_RDATA(M_AXIMM_11_RDATA),
        .M_AXIMM_11_RRESP(M_AXIMM_11_RRESP),
        .M_AXIMM_11_RLAST(M_AXIMM_11_RLAST),
        .M_AXIMM_11_RVALID(M_AXIMM_11_RVALID),
        .M_AXIMM_11_RREADY(M_AXIMM_11_RREADY),
        .AP_AXIMM_12_AWADDR(AP_AXIMM_12_AWADDR),
        .AP_AXIMM_12_AWLEN(AP_AXIMM_12_AWLEN),
        .AP_AXIMM_12_AWSIZE(AP_AXIMM_12_AWSIZE),
        .AP_AXIMM_12_AWBURST(AP_AXIMM_12_AWBURST),
        .AP_AXIMM_12_AWLOCK(AP_AXIMM_12_AWLOCK),
        .AP_AXIMM_12_AWCACHE(AP_AXIMM_12_AWCACHE),
        .AP_AXIMM_12_AWPROT(AP_AXIMM_12_AWPROT),
        .AP_AXIMM_12_AWREGION(AP_AXIMM_12_AWREGION),
        .AP_AXIMM_12_AWQOS(AP_AXIMM_12_AWQOS),
        .AP_AXIMM_12_AWVALID(AP_AXIMM_12_AWVALID),
        .AP_AXIMM_12_AWREADY(AP_AXIMM_12_AWREADY),
        .AP_AXIMM_12_WDATA(AP_AXIMM_12_WDATA),
        .AP_AXIMM_12_WSTRB(AP_AXIMM_12_WSTRB),
        .AP_AXIMM_12_WLAST(AP_AXIMM_12_WLAST),
        .AP_AXIMM_12_WVALID(AP_AXIMM_12_WVALID),
        .AP_AXIMM_12_WREADY(AP_AXIMM_12_WREADY),
        .AP_AXIMM_12_BRESP(AP_AXIMM_12_BRESP),
        .AP_AXIMM_12_BVALID(AP_AXIMM_12_BVALID),
        .AP_AXIMM_12_BREADY(AP_AXIMM_12_BREADY),
        .AP_AXIMM_12_ARADDR(AP_AXIMM_12_ARADDR),
        .AP_AXIMM_12_ARLEN(AP_AXIMM_12_ARLEN),
        .AP_AXIMM_12_ARSIZE(AP_AXIMM_12_ARSIZE),
        .AP_AXIMM_12_ARBURST(AP_AXIMM_12_ARBURST),
        .AP_AXIMM_12_ARLOCK(AP_AXIMM_12_ARLOCK),
        .AP_AXIMM_12_ARCACHE(AP_AXIMM_12_ARCACHE),
        .AP_AXIMM_12_ARPROT(AP_AXIMM_12_ARPROT),
        .AP_AXIMM_12_ARREGION(AP_AXIMM_12_ARREGION),
        .AP_AXIMM_12_ARQOS(AP_AXIMM_12_ARQOS),
        .AP_AXIMM_12_ARVALID(AP_AXIMM_12_ARVALID),
        .AP_AXIMM_12_ARREADY(AP_AXIMM_12_ARREADY),
        .AP_AXIMM_12_RDATA(AP_AXIMM_12_RDATA),
        .AP_AXIMM_12_RRESP(AP_AXIMM_12_RRESP),
        .AP_AXIMM_12_RLAST(AP_AXIMM_12_RLAST),
        .AP_AXIMM_12_RVALID(AP_AXIMM_12_RVALID),
        .AP_AXIMM_12_RREADY(AP_AXIMM_12_RREADY),
        .M_AXIMM_12_AWADDR(M_AXIMM_12_AWADDR),
        .M_AXIMM_12_AWLEN(M_AXIMM_12_AWLEN),
        .M_AXIMM_12_AWSIZE(M_AXIMM_12_AWSIZE),
        .M_AXIMM_12_AWBURST(M_AXIMM_12_AWBURST),
        .M_AXIMM_12_AWLOCK(M_AXIMM_12_AWLOCK),
        .M_AXIMM_12_AWCACHE(M_AXIMM_12_AWCACHE),
        .M_AXIMM_12_AWPROT(M_AXIMM_12_AWPROT),
        .M_AXIMM_12_AWREGION(M_AXIMM_12_AWREGION),
        .M_AXIMM_12_AWQOS(M_AXIMM_12_AWQOS),
        .M_AXIMM_12_AWVALID(M_AXIMM_12_AWVALID),
        .M_AXIMM_12_AWREADY(M_AXIMM_12_AWREADY),
        .M_AXIMM_12_WDATA(M_AXIMM_12_WDATA),
        .M_AXIMM_12_WSTRB(M_AXIMM_12_WSTRB),
        .M_AXIMM_12_WLAST(M_AXIMM_12_WLAST),
        .M_AXIMM_12_WVALID(M_AXIMM_12_WVALID),
        .M_AXIMM_12_WREADY(M_AXIMM_12_WREADY),
        .M_AXIMM_12_BRESP(M_AXIMM_12_BRESP),
        .M_AXIMM_12_BVALID(M_AXIMM_12_BVALID),
        .M_AXIMM_12_BREADY(M_AXIMM_12_BREADY),
        .M_AXIMM_12_ARADDR(M_AXIMM_12_ARADDR),
        .M_AXIMM_12_ARLEN(M_AXIMM_12_ARLEN),
        .M_AXIMM_12_ARSIZE(M_AXIMM_12_ARSIZE),
        .M_AXIMM_12_ARBURST(M_AXIMM_12_ARBURST),
        .M_AXIMM_12_ARLOCK(M_AXIMM_12_ARLOCK),
        .M_AXIMM_12_ARCACHE(M_AXIMM_12_ARCACHE),
        .M_AXIMM_12_ARPROT(M_AXIMM_12_ARPROT),
        .M_AXIMM_12_ARREGION(M_AXIMM_12_ARREGION),
        .M_AXIMM_12_ARQOS(M_AXIMM_12_ARQOS),
        .M_AXIMM_12_ARVALID(M_AXIMM_12_ARVALID),
        .M_AXIMM_12_ARREADY(M_AXIMM_12_ARREADY),
        .M_AXIMM_12_RDATA(M_AXIMM_12_RDATA),
        .M_AXIMM_12_RRESP(M_AXIMM_12_RRESP),
        .M_AXIMM_12_RLAST(M_AXIMM_12_RLAST),
        .M_AXIMM_12_RVALID(M_AXIMM_12_RVALID),
        .M_AXIMM_12_RREADY(M_AXIMM_12_RREADY),
        .AP_AXIMM_13_AWADDR(AP_AXIMM_13_AWADDR),
        .AP_AXIMM_13_AWLEN(AP_AXIMM_13_AWLEN),
        .AP_AXIMM_13_AWSIZE(AP_AXIMM_13_AWSIZE),
        .AP_AXIMM_13_AWBURST(AP_AXIMM_13_AWBURST),
        .AP_AXIMM_13_AWLOCK(AP_AXIMM_13_AWLOCK),
        .AP_AXIMM_13_AWCACHE(AP_AXIMM_13_AWCACHE),
        .AP_AXIMM_13_AWPROT(AP_AXIMM_13_AWPROT),
        .AP_AXIMM_13_AWREGION(AP_AXIMM_13_AWREGION),
        .AP_AXIMM_13_AWQOS(AP_AXIMM_13_AWQOS),
        .AP_AXIMM_13_AWVALID(AP_AXIMM_13_AWVALID),
        .AP_AXIMM_13_AWREADY(AP_AXIMM_13_AWREADY),
        .AP_AXIMM_13_WDATA(AP_AXIMM_13_WDATA),
        .AP_AXIMM_13_WSTRB(AP_AXIMM_13_WSTRB),
        .AP_AXIMM_13_WLAST(AP_AXIMM_13_WLAST),
        .AP_AXIMM_13_WVALID(AP_AXIMM_13_WVALID),
        .AP_AXIMM_13_WREADY(AP_AXIMM_13_WREADY),
        .AP_AXIMM_13_BRESP(AP_AXIMM_13_BRESP),
        .AP_AXIMM_13_BVALID(AP_AXIMM_13_BVALID),
        .AP_AXIMM_13_BREADY(AP_AXIMM_13_BREADY),
        .AP_AXIMM_13_ARADDR(AP_AXIMM_13_ARADDR),
        .AP_AXIMM_13_ARLEN(AP_AXIMM_13_ARLEN),
        .AP_AXIMM_13_ARSIZE(AP_AXIMM_13_ARSIZE),
        .AP_AXIMM_13_ARBURST(AP_AXIMM_13_ARBURST),
        .AP_AXIMM_13_ARLOCK(AP_AXIMM_13_ARLOCK),
        .AP_AXIMM_13_ARCACHE(AP_AXIMM_13_ARCACHE),
        .AP_AXIMM_13_ARPROT(AP_AXIMM_13_ARPROT),
        .AP_AXIMM_13_ARREGION(AP_AXIMM_13_ARREGION),
        .AP_AXIMM_13_ARQOS(AP_AXIMM_13_ARQOS),
        .AP_AXIMM_13_ARVALID(AP_AXIMM_13_ARVALID),
        .AP_AXIMM_13_ARREADY(AP_AXIMM_13_ARREADY),
        .AP_AXIMM_13_RDATA(AP_AXIMM_13_RDATA),
        .AP_AXIMM_13_RRESP(AP_AXIMM_13_RRESP),
        .AP_AXIMM_13_RLAST(AP_AXIMM_13_RLAST),
        .AP_AXIMM_13_RVALID(AP_AXIMM_13_RVALID),
        .AP_AXIMM_13_RREADY(AP_AXIMM_13_RREADY),
        .M_AXIMM_13_AWADDR(M_AXIMM_13_AWADDR),
        .M_AXIMM_13_AWLEN(M_AXIMM_13_AWLEN),
        .M_AXIMM_13_AWSIZE(M_AXIMM_13_AWSIZE),
        .M_AXIMM_13_AWBURST(M_AXIMM_13_AWBURST),
        .M_AXIMM_13_AWLOCK(M_AXIMM_13_AWLOCK),
        .M_AXIMM_13_AWCACHE(M_AXIMM_13_AWCACHE),
        .M_AXIMM_13_AWPROT(M_AXIMM_13_AWPROT),
        .M_AXIMM_13_AWREGION(M_AXIMM_13_AWREGION),
        .M_AXIMM_13_AWQOS(M_AXIMM_13_AWQOS),
        .M_AXIMM_13_AWVALID(M_AXIMM_13_AWVALID),
        .M_AXIMM_13_AWREADY(M_AXIMM_13_AWREADY),
        .M_AXIMM_13_WDATA(M_AXIMM_13_WDATA),
        .M_AXIMM_13_WSTRB(M_AXIMM_13_WSTRB),
        .M_AXIMM_13_WLAST(M_AXIMM_13_WLAST),
        .M_AXIMM_13_WVALID(M_AXIMM_13_WVALID),
        .M_AXIMM_13_WREADY(M_AXIMM_13_WREADY),
        .M_AXIMM_13_BRESP(M_AXIMM_13_BRESP),
        .M_AXIMM_13_BVALID(M_AXIMM_13_BVALID),
        .M_AXIMM_13_BREADY(M_AXIMM_13_BREADY),
        .M_AXIMM_13_ARADDR(M_AXIMM_13_ARADDR),
        .M_AXIMM_13_ARLEN(M_AXIMM_13_ARLEN),
        .M_AXIMM_13_ARSIZE(M_AXIMM_13_ARSIZE),
        .M_AXIMM_13_ARBURST(M_AXIMM_13_ARBURST),
        .M_AXIMM_13_ARLOCK(M_AXIMM_13_ARLOCK),
        .M_AXIMM_13_ARCACHE(M_AXIMM_13_ARCACHE),
        .M_AXIMM_13_ARPROT(M_AXIMM_13_ARPROT),
        .M_AXIMM_13_ARREGION(M_AXIMM_13_ARREGION),
        .M_AXIMM_13_ARQOS(M_AXIMM_13_ARQOS),
        .M_AXIMM_13_ARVALID(M_AXIMM_13_ARVALID),
        .M_AXIMM_13_ARREADY(M_AXIMM_13_ARREADY),
        .M_AXIMM_13_RDATA(M_AXIMM_13_RDATA),
        .M_AXIMM_13_RRESP(M_AXIMM_13_RRESP),
        .M_AXIMM_13_RLAST(M_AXIMM_13_RLAST),
        .M_AXIMM_13_RVALID(M_AXIMM_13_RVALID),
        .M_AXIMM_13_RREADY(M_AXIMM_13_RREADY),
        .AP_AXIMM_14_AWADDR(AP_AXIMM_14_AWADDR),
        .AP_AXIMM_14_AWLEN(AP_AXIMM_14_AWLEN),
        .AP_AXIMM_14_AWSIZE(AP_AXIMM_14_AWSIZE),
        .AP_AXIMM_14_AWBURST(AP_AXIMM_14_AWBURST),
        .AP_AXIMM_14_AWLOCK(AP_AXIMM_14_AWLOCK),
        .AP_AXIMM_14_AWCACHE(AP_AXIMM_14_AWCACHE),
        .AP_AXIMM_14_AWPROT(AP_AXIMM_14_AWPROT),
        .AP_AXIMM_14_AWREGION(AP_AXIMM_14_AWREGION),
        .AP_AXIMM_14_AWQOS(AP_AXIMM_14_AWQOS),
        .AP_AXIMM_14_AWVALID(AP_AXIMM_14_AWVALID),
        .AP_AXIMM_14_AWREADY(AP_AXIMM_14_AWREADY),
        .AP_AXIMM_14_WDATA(AP_AXIMM_14_WDATA),
        .AP_AXIMM_14_WSTRB(AP_AXIMM_14_WSTRB),
        .AP_AXIMM_14_WLAST(AP_AXIMM_14_WLAST),
        .AP_AXIMM_14_WVALID(AP_AXIMM_14_WVALID),
        .AP_AXIMM_14_WREADY(AP_AXIMM_14_WREADY),
        .AP_AXIMM_14_BRESP(AP_AXIMM_14_BRESP),
        .AP_AXIMM_14_BVALID(AP_AXIMM_14_BVALID),
        .AP_AXIMM_14_BREADY(AP_AXIMM_14_BREADY),
        .AP_AXIMM_14_ARADDR(AP_AXIMM_14_ARADDR),
        .AP_AXIMM_14_ARLEN(AP_AXIMM_14_ARLEN),
        .AP_AXIMM_14_ARSIZE(AP_AXIMM_14_ARSIZE),
        .AP_AXIMM_14_ARBURST(AP_AXIMM_14_ARBURST),
        .AP_AXIMM_14_ARLOCK(AP_AXIMM_14_ARLOCK),
        .AP_AXIMM_14_ARCACHE(AP_AXIMM_14_ARCACHE),
        .AP_AXIMM_14_ARPROT(AP_AXIMM_14_ARPROT),
        .AP_AXIMM_14_ARREGION(AP_AXIMM_14_ARREGION),
        .AP_AXIMM_14_ARQOS(AP_AXIMM_14_ARQOS),
        .AP_AXIMM_14_ARVALID(AP_AXIMM_14_ARVALID),
        .AP_AXIMM_14_ARREADY(AP_AXIMM_14_ARREADY),
        .AP_AXIMM_14_RDATA(AP_AXIMM_14_RDATA),
        .AP_AXIMM_14_RRESP(AP_AXIMM_14_RRESP),
        .AP_AXIMM_14_RLAST(AP_AXIMM_14_RLAST),
        .AP_AXIMM_14_RVALID(AP_AXIMM_14_RVALID),
        .AP_AXIMM_14_RREADY(AP_AXIMM_14_RREADY),
        .M_AXIMM_14_AWADDR(M_AXIMM_14_AWADDR),
        .M_AXIMM_14_AWLEN(M_AXIMM_14_AWLEN),
        .M_AXIMM_14_AWSIZE(M_AXIMM_14_AWSIZE),
        .M_AXIMM_14_AWBURST(M_AXIMM_14_AWBURST),
        .M_AXIMM_14_AWLOCK(M_AXIMM_14_AWLOCK),
        .M_AXIMM_14_AWCACHE(M_AXIMM_14_AWCACHE),
        .M_AXIMM_14_AWPROT(M_AXIMM_14_AWPROT),
        .M_AXIMM_14_AWREGION(M_AXIMM_14_AWREGION),
        .M_AXIMM_14_AWQOS(M_AXIMM_14_AWQOS),
        .M_AXIMM_14_AWVALID(M_AXIMM_14_AWVALID),
        .M_AXIMM_14_AWREADY(M_AXIMM_14_AWREADY),
        .M_AXIMM_14_WDATA(M_AXIMM_14_WDATA),
        .M_AXIMM_14_WSTRB(M_AXIMM_14_WSTRB),
        .M_AXIMM_14_WLAST(M_AXIMM_14_WLAST),
        .M_AXIMM_14_WVALID(M_AXIMM_14_WVALID),
        .M_AXIMM_14_WREADY(M_AXIMM_14_WREADY),
        .M_AXIMM_14_BRESP(M_AXIMM_14_BRESP),
        .M_AXIMM_14_BVALID(M_AXIMM_14_BVALID),
        .M_AXIMM_14_BREADY(M_AXIMM_14_BREADY),
        .M_AXIMM_14_ARADDR(M_AXIMM_14_ARADDR),
        .M_AXIMM_14_ARLEN(M_AXIMM_14_ARLEN),
        .M_AXIMM_14_ARSIZE(M_AXIMM_14_ARSIZE),
        .M_AXIMM_14_ARBURST(M_AXIMM_14_ARBURST),
        .M_AXIMM_14_ARLOCK(M_AXIMM_14_ARLOCK),
        .M_AXIMM_14_ARCACHE(M_AXIMM_14_ARCACHE),
        .M_AXIMM_14_ARPROT(M_AXIMM_14_ARPROT),
        .M_AXIMM_14_ARREGION(M_AXIMM_14_ARREGION),
        .M_AXIMM_14_ARQOS(M_AXIMM_14_ARQOS),
        .M_AXIMM_14_ARVALID(M_AXIMM_14_ARVALID),
        .M_AXIMM_14_ARREADY(M_AXIMM_14_ARREADY),
        .M_AXIMM_14_RDATA(M_AXIMM_14_RDATA),
        .M_AXIMM_14_RRESP(M_AXIMM_14_RRESP),
        .M_AXIMM_14_RLAST(M_AXIMM_14_RLAST),
        .M_AXIMM_14_RVALID(M_AXIMM_14_RVALID),
        .M_AXIMM_14_RREADY(M_AXIMM_14_RREADY),
        .AP_AXIMM_15_AWADDR(AP_AXIMM_15_AWADDR),
        .AP_AXIMM_15_AWLEN(AP_AXIMM_15_AWLEN),
        .AP_AXIMM_15_AWSIZE(AP_AXIMM_15_AWSIZE),
        .AP_AXIMM_15_AWBURST(AP_AXIMM_15_AWBURST),
        .AP_AXIMM_15_AWLOCK(AP_AXIMM_15_AWLOCK),
        .AP_AXIMM_15_AWCACHE(AP_AXIMM_15_AWCACHE),
        .AP_AXIMM_15_AWPROT(AP_AXIMM_15_AWPROT),
        .AP_AXIMM_15_AWREGION(AP_AXIMM_15_AWREGION),
        .AP_AXIMM_15_AWQOS(AP_AXIMM_15_AWQOS),
        .AP_AXIMM_15_AWVALID(AP_AXIMM_15_AWVALID),
        .AP_AXIMM_15_AWREADY(AP_AXIMM_15_AWREADY),
        .AP_AXIMM_15_WDATA(AP_AXIMM_15_WDATA),
        .AP_AXIMM_15_WSTRB(AP_AXIMM_15_WSTRB),
        .AP_AXIMM_15_WLAST(AP_AXIMM_15_WLAST),
        .AP_AXIMM_15_WVALID(AP_AXIMM_15_WVALID),
        .AP_AXIMM_15_WREADY(AP_AXIMM_15_WREADY),
        .AP_AXIMM_15_BRESP(AP_AXIMM_15_BRESP),
        .AP_AXIMM_15_BVALID(AP_AXIMM_15_BVALID),
        .AP_AXIMM_15_BREADY(AP_AXIMM_15_BREADY),
        .AP_AXIMM_15_ARADDR(AP_AXIMM_15_ARADDR),
        .AP_AXIMM_15_ARLEN(AP_AXIMM_15_ARLEN),
        .AP_AXIMM_15_ARSIZE(AP_AXIMM_15_ARSIZE),
        .AP_AXIMM_15_ARBURST(AP_AXIMM_15_ARBURST),
        .AP_AXIMM_15_ARLOCK(AP_AXIMM_15_ARLOCK),
        .AP_AXIMM_15_ARCACHE(AP_AXIMM_15_ARCACHE),
        .AP_AXIMM_15_ARPROT(AP_AXIMM_15_ARPROT),
        .AP_AXIMM_15_ARREGION(AP_AXIMM_15_ARREGION),
        .AP_AXIMM_15_ARQOS(AP_AXIMM_15_ARQOS),
        .AP_AXIMM_15_ARVALID(AP_AXIMM_15_ARVALID),
        .AP_AXIMM_15_ARREADY(AP_AXIMM_15_ARREADY),
        .AP_AXIMM_15_RDATA(AP_AXIMM_15_RDATA),
        .AP_AXIMM_15_RRESP(AP_AXIMM_15_RRESP),
        .AP_AXIMM_15_RLAST(AP_AXIMM_15_RLAST),
        .AP_AXIMM_15_RVALID(AP_AXIMM_15_RVALID),
        .AP_AXIMM_15_RREADY(AP_AXIMM_15_RREADY),
        .M_AXIMM_15_AWADDR(M_AXIMM_15_AWADDR),
        .M_AXIMM_15_AWLEN(M_AXIMM_15_AWLEN),
        .M_AXIMM_15_AWSIZE(M_AXIMM_15_AWSIZE),
        .M_AXIMM_15_AWBURST(M_AXIMM_15_AWBURST),
        .M_AXIMM_15_AWLOCK(M_AXIMM_15_AWLOCK),
        .M_AXIMM_15_AWCACHE(M_AXIMM_15_AWCACHE),
        .M_AXIMM_15_AWPROT(M_AXIMM_15_AWPROT),
        .M_AXIMM_15_AWREGION(M_AXIMM_15_AWREGION),
        .M_AXIMM_15_AWQOS(M_AXIMM_15_AWQOS),
        .M_AXIMM_15_AWVALID(M_AXIMM_15_AWVALID),
        .M_AXIMM_15_AWREADY(M_AXIMM_15_AWREADY),
        .M_AXIMM_15_WDATA(M_AXIMM_15_WDATA),
        .M_AXIMM_15_WSTRB(M_AXIMM_15_WSTRB),
        .M_AXIMM_15_WLAST(M_AXIMM_15_WLAST),
        .M_AXIMM_15_WVALID(M_AXIMM_15_WVALID),
        .M_AXIMM_15_WREADY(M_AXIMM_15_WREADY),
        .M_AXIMM_15_BRESP(M_AXIMM_15_BRESP),
        .M_AXIMM_15_BVALID(M_AXIMM_15_BVALID),
        .M_AXIMM_15_BREADY(M_AXIMM_15_BREADY),
        .M_AXIMM_15_ARADDR(M_AXIMM_15_ARADDR),
        .M_AXIMM_15_ARLEN(M_AXIMM_15_ARLEN),
        .M_AXIMM_15_ARSIZE(M_AXIMM_15_ARSIZE),
        .M_AXIMM_15_ARBURST(M_AXIMM_15_ARBURST),
        .M_AXIMM_15_ARLOCK(M_AXIMM_15_ARLOCK),
        .M_AXIMM_15_ARCACHE(M_AXIMM_15_ARCACHE),
        .M_AXIMM_15_ARPROT(M_AXIMM_15_ARPROT),
        .M_AXIMM_15_ARREGION(M_AXIMM_15_ARREGION),
        .M_AXIMM_15_ARQOS(M_AXIMM_15_ARQOS),
        .M_AXIMM_15_ARVALID(M_AXIMM_15_ARVALID),
        .M_AXIMM_15_ARREADY(M_AXIMM_15_ARREADY),
        .M_AXIMM_15_RDATA(M_AXIMM_15_RDATA),
        .M_AXIMM_15_RRESP(M_AXIMM_15_RRESP),
        .M_AXIMM_15_RLAST(M_AXIMM_15_RLAST),
        .M_AXIMM_15_RVALID(M_AXIMM_15_RVALID),
        .M_AXIMM_15_RREADY(M_AXIMM_15_RREADY),
        .AP_AXIMM_16_AWADDR(AP_AXIMM_16_AWADDR),
        .AP_AXIMM_16_AWLEN(AP_AXIMM_16_AWLEN),
        .AP_AXIMM_16_AWSIZE(AP_AXIMM_16_AWSIZE),
        .AP_AXIMM_16_AWBURST(AP_AXIMM_16_AWBURST),
        .AP_AXIMM_16_AWLOCK(AP_AXIMM_16_AWLOCK),
        .AP_AXIMM_16_AWCACHE(AP_AXIMM_16_AWCACHE),
        .AP_AXIMM_16_AWPROT(AP_AXIMM_16_AWPROT),
        .AP_AXIMM_16_AWREGION(AP_AXIMM_16_AWREGION),
        .AP_AXIMM_16_AWQOS(AP_AXIMM_16_AWQOS),
        .AP_AXIMM_16_AWVALID(AP_AXIMM_16_AWVALID),
        .AP_AXIMM_16_AWREADY(AP_AXIMM_16_AWREADY),
        .AP_AXIMM_16_WDATA(AP_AXIMM_16_WDATA),
        .AP_AXIMM_16_WSTRB(AP_AXIMM_16_WSTRB),
        .AP_AXIMM_16_WLAST(AP_AXIMM_16_WLAST),
        .AP_AXIMM_16_WVALID(AP_AXIMM_16_WVALID),
        .AP_AXIMM_16_WREADY(AP_AXIMM_16_WREADY),
        .AP_AXIMM_16_BRESP(AP_AXIMM_16_BRESP),
        .AP_AXIMM_16_BVALID(AP_AXIMM_16_BVALID),
        .AP_AXIMM_16_BREADY(AP_AXIMM_16_BREADY),
        .AP_AXIMM_16_ARADDR(AP_AXIMM_16_ARADDR),
        .AP_AXIMM_16_ARLEN(AP_AXIMM_16_ARLEN),
        .AP_AXIMM_16_ARSIZE(AP_AXIMM_16_ARSIZE),
        .AP_AXIMM_16_ARBURST(AP_AXIMM_16_ARBURST),
        .AP_AXIMM_16_ARLOCK(AP_AXIMM_16_ARLOCK),
        .AP_AXIMM_16_ARCACHE(AP_AXIMM_16_ARCACHE),
        .AP_AXIMM_16_ARPROT(AP_AXIMM_16_ARPROT),
        .AP_AXIMM_16_ARREGION(AP_AXIMM_16_ARREGION),
        .AP_AXIMM_16_ARQOS(AP_AXIMM_16_ARQOS),
        .AP_AXIMM_16_ARVALID(AP_AXIMM_16_ARVALID),
        .AP_AXIMM_16_ARREADY(AP_AXIMM_16_ARREADY),
        .AP_AXIMM_16_RDATA(AP_AXIMM_16_RDATA),
        .AP_AXIMM_16_RRESP(AP_AXIMM_16_RRESP),
        .AP_AXIMM_16_RLAST(AP_AXIMM_16_RLAST),
        .AP_AXIMM_16_RVALID(AP_AXIMM_16_RVALID),
        .AP_AXIMM_16_RREADY(AP_AXIMM_16_RREADY),
        .M_AXIMM_16_AWADDR(M_AXIMM_16_AWADDR),
        .M_AXIMM_16_AWLEN(M_AXIMM_16_AWLEN),
        .M_AXIMM_16_AWSIZE(M_AXIMM_16_AWSIZE),
        .M_AXIMM_16_AWBURST(M_AXIMM_16_AWBURST),
        .M_AXIMM_16_AWLOCK(M_AXIMM_16_AWLOCK),
        .M_AXIMM_16_AWCACHE(M_AXIMM_16_AWCACHE),
        .M_AXIMM_16_AWPROT(M_AXIMM_16_AWPROT),
        .M_AXIMM_16_AWREGION(M_AXIMM_16_AWREGION),
        .M_AXIMM_16_AWQOS(M_AXIMM_16_AWQOS),
        .M_AXIMM_16_AWVALID(M_AXIMM_16_AWVALID),
        .M_AXIMM_16_AWREADY(M_AXIMM_16_AWREADY),
        .M_AXIMM_16_WDATA(M_AXIMM_16_WDATA),
        .M_AXIMM_16_WSTRB(M_AXIMM_16_WSTRB),
        .M_AXIMM_16_WLAST(M_AXIMM_16_WLAST),
        .M_AXIMM_16_WVALID(M_AXIMM_16_WVALID),
        .M_AXIMM_16_WREADY(M_AXIMM_16_WREADY),
        .M_AXIMM_16_BRESP(M_AXIMM_16_BRESP),
        .M_AXIMM_16_BVALID(M_AXIMM_16_BVALID),
        .M_AXIMM_16_BREADY(M_AXIMM_16_BREADY),
        .M_AXIMM_16_ARADDR(M_AXIMM_16_ARADDR),
        .M_AXIMM_16_ARLEN(M_AXIMM_16_ARLEN),
        .M_AXIMM_16_ARSIZE(M_AXIMM_16_ARSIZE),
        .M_AXIMM_16_ARBURST(M_AXIMM_16_ARBURST),
        .M_AXIMM_16_ARLOCK(M_AXIMM_16_ARLOCK),
        .M_AXIMM_16_ARCACHE(M_AXIMM_16_ARCACHE),
        .M_AXIMM_16_ARPROT(M_AXIMM_16_ARPROT),
        .M_AXIMM_16_ARREGION(M_AXIMM_16_ARREGION),
        .M_AXIMM_16_ARQOS(M_AXIMM_16_ARQOS),
        .M_AXIMM_16_ARVALID(M_AXIMM_16_ARVALID),
        .M_AXIMM_16_ARREADY(M_AXIMM_16_ARREADY),
        .M_AXIMM_16_RDATA(M_AXIMM_16_RDATA),
        .M_AXIMM_16_RRESP(M_AXIMM_16_RRESP),
        .M_AXIMM_16_RLAST(M_AXIMM_16_RLAST),
        .M_AXIMM_16_RVALID(M_AXIMM_16_RVALID),
        .M_AXIMM_16_RREADY(M_AXIMM_16_RREADY),
        .AP_AXIMM_17_AWADDR(AP_AXIMM_17_AWADDR),
        .AP_AXIMM_17_AWLEN(AP_AXIMM_17_AWLEN),
        .AP_AXIMM_17_AWSIZE(AP_AXIMM_17_AWSIZE),
        .AP_AXIMM_17_AWBURST(AP_AXIMM_17_AWBURST),
        .AP_AXIMM_17_AWLOCK(AP_AXIMM_17_AWLOCK),
        .AP_AXIMM_17_AWCACHE(AP_AXIMM_17_AWCACHE),
        .AP_AXIMM_17_AWPROT(AP_AXIMM_17_AWPROT),
        .AP_AXIMM_17_AWREGION(AP_AXIMM_17_AWREGION),
        .AP_AXIMM_17_AWQOS(AP_AXIMM_17_AWQOS),
        .AP_AXIMM_17_AWVALID(AP_AXIMM_17_AWVALID),
        .AP_AXIMM_17_AWREADY(AP_AXIMM_17_AWREADY),
        .AP_AXIMM_17_WDATA(AP_AXIMM_17_WDATA),
        .AP_AXIMM_17_WSTRB(AP_AXIMM_17_WSTRB),
        .AP_AXIMM_17_WLAST(AP_AXIMM_17_WLAST),
        .AP_AXIMM_17_WVALID(AP_AXIMM_17_WVALID),
        .AP_AXIMM_17_WREADY(AP_AXIMM_17_WREADY),
        .AP_AXIMM_17_BRESP(AP_AXIMM_17_BRESP),
        .AP_AXIMM_17_BVALID(AP_AXIMM_17_BVALID),
        .AP_AXIMM_17_BREADY(AP_AXIMM_17_BREADY),
        .AP_AXIMM_17_ARADDR(AP_AXIMM_17_ARADDR),
        .AP_AXIMM_17_ARLEN(AP_AXIMM_17_ARLEN),
        .AP_AXIMM_17_ARSIZE(AP_AXIMM_17_ARSIZE),
        .AP_AXIMM_17_ARBURST(AP_AXIMM_17_ARBURST),
        .AP_AXIMM_17_ARLOCK(AP_AXIMM_17_ARLOCK),
        .AP_AXIMM_17_ARCACHE(AP_AXIMM_17_ARCACHE),
        .AP_AXIMM_17_ARPROT(AP_AXIMM_17_ARPROT),
        .AP_AXIMM_17_ARREGION(AP_AXIMM_17_ARREGION),
        .AP_AXIMM_17_ARQOS(AP_AXIMM_17_ARQOS),
        .AP_AXIMM_17_ARVALID(AP_AXIMM_17_ARVALID),
        .AP_AXIMM_17_ARREADY(AP_AXIMM_17_ARREADY),
        .AP_AXIMM_17_RDATA(AP_AXIMM_17_RDATA),
        .AP_AXIMM_17_RRESP(AP_AXIMM_17_RRESP),
        .AP_AXIMM_17_RLAST(AP_AXIMM_17_RLAST),
        .AP_AXIMM_17_RVALID(AP_AXIMM_17_RVALID),
        .AP_AXIMM_17_RREADY(AP_AXIMM_17_RREADY),
        .M_AXIMM_17_AWADDR(M_AXIMM_17_AWADDR),
        .M_AXIMM_17_AWLEN(M_AXIMM_17_AWLEN),
        .M_AXIMM_17_AWSIZE(M_AXIMM_17_AWSIZE),
        .M_AXIMM_17_AWBURST(M_AXIMM_17_AWBURST),
        .M_AXIMM_17_AWLOCK(M_AXIMM_17_AWLOCK),
        .M_AXIMM_17_AWCACHE(M_AXIMM_17_AWCACHE),
        .M_AXIMM_17_AWPROT(M_AXIMM_17_AWPROT),
        .M_AXIMM_17_AWREGION(M_AXIMM_17_AWREGION),
        .M_AXIMM_17_AWQOS(M_AXIMM_17_AWQOS),
        .M_AXIMM_17_AWVALID(M_AXIMM_17_AWVALID),
        .M_AXIMM_17_AWREADY(M_AXIMM_17_AWREADY),
        .M_AXIMM_17_WDATA(M_AXIMM_17_WDATA),
        .M_AXIMM_17_WSTRB(M_AXIMM_17_WSTRB),
        .M_AXIMM_17_WLAST(M_AXIMM_17_WLAST),
        .M_AXIMM_17_WVALID(M_AXIMM_17_WVALID),
        .M_AXIMM_17_WREADY(M_AXIMM_17_WREADY),
        .M_AXIMM_17_BRESP(M_AXIMM_17_BRESP),
        .M_AXIMM_17_BVALID(M_AXIMM_17_BVALID),
        .M_AXIMM_17_BREADY(M_AXIMM_17_BREADY),
        .M_AXIMM_17_ARADDR(M_AXIMM_17_ARADDR),
        .M_AXIMM_17_ARLEN(M_AXIMM_17_ARLEN),
        .M_AXIMM_17_ARSIZE(M_AXIMM_17_ARSIZE),
        .M_AXIMM_17_ARBURST(M_AXIMM_17_ARBURST),
        .M_AXIMM_17_ARLOCK(M_AXIMM_17_ARLOCK),
        .M_AXIMM_17_ARCACHE(M_AXIMM_17_ARCACHE),
        .M_AXIMM_17_ARPROT(M_AXIMM_17_ARPROT),
        .M_AXIMM_17_ARREGION(M_AXIMM_17_ARREGION),
        .M_AXIMM_17_ARQOS(M_AXIMM_17_ARQOS),
        .M_AXIMM_17_ARVALID(M_AXIMM_17_ARVALID),
        .M_AXIMM_17_ARREADY(M_AXIMM_17_ARREADY),
        .M_AXIMM_17_RDATA(M_AXIMM_17_RDATA),
        .M_AXIMM_17_RRESP(M_AXIMM_17_RRESP),
        .M_AXIMM_17_RLAST(M_AXIMM_17_RLAST),
        .M_AXIMM_17_RVALID(M_AXIMM_17_RVALID),
        .M_AXIMM_17_RREADY(M_AXIMM_17_RREADY),
        .AP_AXIMM_18_AWADDR(AP_AXIMM_18_AWADDR),
        .AP_AXIMM_18_AWLEN(AP_AXIMM_18_AWLEN),
        .AP_AXIMM_18_AWSIZE(AP_AXIMM_18_AWSIZE),
        .AP_AXIMM_18_AWBURST(AP_AXIMM_18_AWBURST),
        .AP_AXIMM_18_AWLOCK(AP_AXIMM_18_AWLOCK),
        .AP_AXIMM_18_AWCACHE(AP_AXIMM_18_AWCACHE),
        .AP_AXIMM_18_AWPROT(AP_AXIMM_18_AWPROT),
        .AP_AXIMM_18_AWREGION(AP_AXIMM_18_AWREGION),
        .AP_AXIMM_18_AWQOS(AP_AXIMM_18_AWQOS),
        .AP_AXIMM_18_AWVALID(AP_AXIMM_18_AWVALID),
        .AP_AXIMM_18_AWREADY(AP_AXIMM_18_AWREADY),
        .AP_AXIMM_18_WDATA(AP_AXIMM_18_WDATA),
        .AP_AXIMM_18_WSTRB(AP_AXIMM_18_WSTRB),
        .AP_AXIMM_18_WLAST(AP_AXIMM_18_WLAST),
        .AP_AXIMM_18_WVALID(AP_AXIMM_18_WVALID),
        .AP_AXIMM_18_WREADY(AP_AXIMM_18_WREADY),
        .AP_AXIMM_18_BRESP(AP_AXIMM_18_BRESP),
        .AP_AXIMM_18_BVALID(AP_AXIMM_18_BVALID),
        .AP_AXIMM_18_BREADY(AP_AXIMM_18_BREADY),
        .AP_AXIMM_18_ARADDR(AP_AXIMM_18_ARADDR),
        .AP_AXIMM_18_ARLEN(AP_AXIMM_18_ARLEN),
        .AP_AXIMM_18_ARSIZE(AP_AXIMM_18_ARSIZE),
        .AP_AXIMM_18_ARBURST(AP_AXIMM_18_ARBURST),
        .AP_AXIMM_18_ARLOCK(AP_AXIMM_18_ARLOCK),
        .AP_AXIMM_18_ARCACHE(AP_AXIMM_18_ARCACHE),
        .AP_AXIMM_18_ARPROT(AP_AXIMM_18_ARPROT),
        .AP_AXIMM_18_ARREGION(AP_AXIMM_18_ARREGION),
        .AP_AXIMM_18_ARQOS(AP_AXIMM_18_ARQOS),
        .AP_AXIMM_18_ARVALID(AP_AXIMM_18_ARVALID),
        .AP_AXIMM_18_ARREADY(AP_AXIMM_18_ARREADY),
        .AP_AXIMM_18_RDATA(AP_AXIMM_18_RDATA),
        .AP_AXIMM_18_RRESP(AP_AXIMM_18_RRESP),
        .AP_AXIMM_18_RLAST(AP_AXIMM_18_RLAST),
        .AP_AXIMM_18_RVALID(AP_AXIMM_18_RVALID),
        .AP_AXIMM_18_RREADY(AP_AXIMM_18_RREADY),
        .M_AXIMM_18_AWADDR(M_AXIMM_18_AWADDR),
        .M_AXIMM_18_AWLEN(M_AXIMM_18_AWLEN),
        .M_AXIMM_18_AWSIZE(M_AXIMM_18_AWSIZE),
        .M_AXIMM_18_AWBURST(M_AXIMM_18_AWBURST),
        .M_AXIMM_18_AWLOCK(M_AXIMM_18_AWLOCK),
        .M_AXIMM_18_AWCACHE(M_AXIMM_18_AWCACHE),
        .M_AXIMM_18_AWPROT(M_AXIMM_18_AWPROT),
        .M_AXIMM_18_AWREGION(M_AXIMM_18_AWREGION),
        .M_AXIMM_18_AWQOS(M_AXIMM_18_AWQOS),
        .M_AXIMM_18_AWVALID(M_AXIMM_18_AWVALID),
        .M_AXIMM_18_AWREADY(M_AXIMM_18_AWREADY),
        .M_AXIMM_18_WDATA(M_AXIMM_18_WDATA),
        .M_AXIMM_18_WSTRB(M_AXIMM_18_WSTRB),
        .M_AXIMM_18_WLAST(M_AXIMM_18_WLAST),
        .M_AXIMM_18_WVALID(M_AXIMM_18_WVALID),
        .M_AXIMM_18_WREADY(M_AXIMM_18_WREADY),
        .M_AXIMM_18_BRESP(M_AXIMM_18_BRESP),
        .M_AXIMM_18_BVALID(M_AXIMM_18_BVALID),
        .M_AXIMM_18_BREADY(M_AXIMM_18_BREADY),
        .M_AXIMM_18_ARADDR(M_AXIMM_18_ARADDR),
        .M_AXIMM_18_ARLEN(M_AXIMM_18_ARLEN),
        .M_AXIMM_18_ARSIZE(M_AXIMM_18_ARSIZE),
        .M_AXIMM_18_ARBURST(M_AXIMM_18_ARBURST),
        .M_AXIMM_18_ARLOCK(M_AXIMM_18_ARLOCK),
        .M_AXIMM_18_ARCACHE(M_AXIMM_18_ARCACHE),
        .M_AXIMM_18_ARPROT(M_AXIMM_18_ARPROT),
        .M_AXIMM_18_ARREGION(M_AXIMM_18_ARREGION),
        .M_AXIMM_18_ARQOS(M_AXIMM_18_ARQOS),
        .M_AXIMM_18_ARVALID(M_AXIMM_18_ARVALID),
        .M_AXIMM_18_ARREADY(M_AXIMM_18_ARREADY),
        .M_AXIMM_18_RDATA(M_AXIMM_18_RDATA),
        .M_AXIMM_18_RRESP(M_AXIMM_18_RRESP),
        .M_AXIMM_18_RLAST(M_AXIMM_18_RLAST),
        .M_AXIMM_18_RVALID(M_AXIMM_18_RVALID),
        .M_AXIMM_18_RREADY(M_AXIMM_18_RREADY),
        .AP_AXIMM_19_AWADDR(AP_AXIMM_19_AWADDR),
        .AP_AXIMM_19_AWLEN(AP_AXIMM_19_AWLEN),
        .AP_AXIMM_19_AWSIZE(AP_AXIMM_19_AWSIZE),
        .AP_AXIMM_19_AWBURST(AP_AXIMM_19_AWBURST),
        .AP_AXIMM_19_AWLOCK(AP_AXIMM_19_AWLOCK),
        .AP_AXIMM_19_AWCACHE(AP_AXIMM_19_AWCACHE),
        .AP_AXIMM_19_AWPROT(AP_AXIMM_19_AWPROT),
        .AP_AXIMM_19_AWREGION(AP_AXIMM_19_AWREGION),
        .AP_AXIMM_19_AWQOS(AP_AXIMM_19_AWQOS),
        .AP_AXIMM_19_AWVALID(AP_AXIMM_19_AWVALID),
        .AP_AXIMM_19_AWREADY(AP_AXIMM_19_AWREADY),
        .AP_AXIMM_19_WDATA(AP_AXIMM_19_WDATA),
        .AP_AXIMM_19_WSTRB(AP_AXIMM_19_WSTRB),
        .AP_AXIMM_19_WLAST(AP_AXIMM_19_WLAST),
        .AP_AXIMM_19_WVALID(AP_AXIMM_19_WVALID),
        .AP_AXIMM_19_WREADY(AP_AXIMM_19_WREADY),
        .AP_AXIMM_19_BRESP(AP_AXIMM_19_BRESP),
        .AP_AXIMM_19_BVALID(AP_AXIMM_19_BVALID),
        .AP_AXIMM_19_BREADY(AP_AXIMM_19_BREADY),
        .AP_AXIMM_19_ARADDR(AP_AXIMM_19_ARADDR),
        .AP_AXIMM_19_ARLEN(AP_AXIMM_19_ARLEN),
        .AP_AXIMM_19_ARSIZE(AP_AXIMM_19_ARSIZE),
        .AP_AXIMM_19_ARBURST(AP_AXIMM_19_ARBURST),
        .AP_AXIMM_19_ARLOCK(AP_AXIMM_19_ARLOCK),
        .AP_AXIMM_19_ARCACHE(AP_AXIMM_19_ARCACHE),
        .AP_AXIMM_19_ARPROT(AP_AXIMM_19_ARPROT),
        .AP_AXIMM_19_ARREGION(AP_AXIMM_19_ARREGION),
        .AP_AXIMM_19_ARQOS(AP_AXIMM_19_ARQOS),
        .AP_AXIMM_19_ARVALID(AP_AXIMM_19_ARVALID),
        .AP_AXIMM_19_ARREADY(AP_AXIMM_19_ARREADY),
        .AP_AXIMM_19_RDATA(AP_AXIMM_19_RDATA),
        .AP_AXIMM_19_RRESP(AP_AXIMM_19_RRESP),
        .AP_AXIMM_19_RLAST(AP_AXIMM_19_RLAST),
        .AP_AXIMM_19_RVALID(AP_AXIMM_19_RVALID),
        .AP_AXIMM_19_RREADY(AP_AXIMM_19_RREADY),
        .M_AXIMM_19_AWADDR(M_AXIMM_19_AWADDR),
        .M_AXIMM_19_AWLEN(M_AXIMM_19_AWLEN),
        .M_AXIMM_19_AWSIZE(M_AXIMM_19_AWSIZE),
        .M_AXIMM_19_AWBURST(M_AXIMM_19_AWBURST),
        .M_AXIMM_19_AWLOCK(M_AXIMM_19_AWLOCK),
        .M_AXIMM_19_AWCACHE(M_AXIMM_19_AWCACHE),
        .M_AXIMM_19_AWPROT(M_AXIMM_19_AWPROT),
        .M_AXIMM_19_AWREGION(M_AXIMM_19_AWREGION),
        .M_AXIMM_19_AWQOS(M_AXIMM_19_AWQOS),
        .M_AXIMM_19_AWVALID(M_AXIMM_19_AWVALID),
        .M_AXIMM_19_AWREADY(M_AXIMM_19_AWREADY),
        .M_AXIMM_19_WDATA(M_AXIMM_19_WDATA),
        .M_AXIMM_19_WSTRB(M_AXIMM_19_WSTRB),
        .M_AXIMM_19_WLAST(M_AXIMM_19_WLAST),
        .M_AXIMM_19_WVALID(M_AXIMM_19_WVALID),
        .M_AXIMM_19_WREADY(M_AXIMM_19_WREADY),
        .M_AXIMM_19_BRESP(M_AXIMM_19_BRESP),
        .M_AXIMM_19_BVALID(M_AXIMM_19_BVALID),
        .M_AXIMM_19_BREADY(M_AXIMM_19_BREADY),
        .M_AXIMM_19_ARADDR(M_AXIMM_19_ARADDR),
        .M_AXIMM_19_ARLEN(M_AXIMM_19_ARLEN),
        .M_AXIMM_19_ARSIZE(M_AXIMM_19_ARSIZE),
        .M_AXIMM_19_ARBURST(M_AXIMM_19_ARBURST),
        .M_AXIMM_19_ARLOCK(M_AXIMM_19_ARLOCK),
        .M_AXIMM_19_ARCACHE(M_AXIMM_19_ARCACHE),
        .M_AXIMM_19_ARPROT(M_AXIMM_19_ARPROT),
        .M_AXIMM_19_ARREGION(M_AXIMM_19_ARREGION),
        .M_AXIMM_19_ARQOS(M_AXIMM_19_ARQOS),
        .M_AXIMM_19_ARVALID(M_AXIMM_19_ARVALID),
        .M_AXIMM_19_ARREADY(M_AXIMM_19_ARREADY),
        .M_AXIMM_19_RDATA(M_AXIMM_19_RDATA),
        .M_AXIMM_19_RRESP(M_AXIMM_19_RRESP),
        .M_AXIMM_19_RLAST(M_AXIMM_19_RLAST),
        .M_AXIMM_19_RVALID(M_AXIMM_19_RVALID),
        .M_AXIMM_19_RREADY(M_AXIMM_19_RREADY),
        .AP_AXIMM_20_AWADDR(AP_AXIMM_20_AWADDR),
        .AP_AXIMM_20_AWLEN(AP_AXIMM_20_AWLEN),
        .AP_AXIMM_20_AWSIZE(AP_AXIMM_20_AWSIZE),
        .AP_AXIMM_20_AWBURST(AP_AXIMM_20_AWBURST),
        .AP_AXIMM_20_AWLOCK(AP_AXIMM_20_AWLOCK),
        .AP_AXIMM_20_AWCACHE(AP_AXIMM_20_AWCACHE),
        .AP_AXIMM_20_AWPROT(AP_AXIMM_20_AWPROT),
        .AP_AXIMM_20_AWREGION(AP_AXIMM_20_AWREGION),
        .AP_AXIMM_20_AWQOS(AP_AXIMM_20_AWQOS),
        .AP_AXIMM_20_AWVALID(AP_AXIMM_20_AWVALID),
        .AP_AXIMM_20_AWREADY(AP_AXIMM_20_AWREADY),
        .AP_AXIMM_20_WDATA(AP_AXIMM_20_WDATA),
        .AP_AXIMM_20_WSTRB(AP_AXIMM_20_WSTRB),
        .AP_AXIMM_20_WLAST(AP_AXIMM_20_WLAST),
        .AP_AXIMM_20_WVALID(AP_AXIMM_20_WVALID),
        .AP_AXIMM_20_WREADY(AP_AXIMM_20_WREADY),
        .AP_AXIMM_20_BRESP(AP_AXIMM_20_BRESP),
        .AP_AXIMM_20_BVALID(AP_AXIMM_20_BVALID),
        .AP_AXIMM_20_BREADY(AP_AXIMM_20_BREADY),
        .AP_AXIMM_20_ARADDR(AP_AXIMM_20_ARADDR),
        .AP_AXIMM_20_ARLEN(AP_AXIMM_20_ARLEN),
        .AP_AXIMM_20_ARSIZE(AP_AXIMM_20_ARSIZE),
        .AP_AXIMM_20_ARBURST(AP_AXIMM_20_ARBURST),
        .AP_AXIMM_20_ARLOCK(AP_AXIMM_20_ARLOCK),
        .AP_AXIMM_20_ARCACHE(AP_AXIMM_20_ARCACHE),
        .AP_AXIMM_20_ARPROT(AP_AXIMM_20_ARPROT),
        .AP_AXIMM_20_ARREGION(AP_AXIMM_20_ARREGION),
        .AP_AXIMM_20_ARQOS(AP_AXIMM_20_ARQOS),
        .AP_AXIMM_20_ARVALID(AP_AXIMM_20_ARVALID),
        .AP_AXIMM_20_ARREADY(AP_AXIMM_20_ARREADY),
        .AP_AXIMM_20_RDATA(AP_AXIMM_20_RDATA),
        .AP_AXIMM_20_RRESP(AP_AXIMM_20_RRESP),
        .AP_AXIMM_20_RLAST(AP_AXIMM_20_RLAST),
        .AP_AXIMM_20_RVALID(AP_AXIMM_20_RVALID),
        .AP_AXIMM_20_RREADY(AP_AXIMM_20_RREADY),
        .M_AXIMM_20_AWADDR(M_AXIMM_20_AWADDR),
        .M_AXIMM_20_AWLEN(M_AXIMM_20_AWLEN),
        .M_AXIMM_20_AWSIZE(M_AXIMM_20_AWSIZE),
        .M_AXIMM_20_AWBURST(M_AXIMM_20_AWBURST),
        .M_AXIMM_20_AWLOCK(M_AXIMM_20_AWLOCK),
        .M_AXIMM_20_AWCACHE(M_AXIMM_20_AWCACHE),
        .M_AXIMM_20_AWPROT(M_AXIMM_20_AWPROT),
        .M_AXIMM_20_AWREGION(M_AXIMM_20_AWREGION),
        .M_AXIMM_20_AWQOS(M_AXIMM_20_AWQOS),
        .M_AXIMM_20_AWVALID(M_AXIMM_20_AWVALID),
        .M_AXIMM_20_AWREADY(M_AXIMM_20_AWREADY),
        .M_AXIMM_20_WDATA(M_AXIMM_20_WDATA),
        .M_AXIMM_20_WSTRB(M_AXIMM_20_WSTRB),
        .M_AXIMM_20_WLAST(M_AXIMM_20_WLAST),
        .M_AXIMM_20_WVALID(M_AXIMM_20_WVALID),
        .M_AXIMM_20_WREADY(M_AXIMM_20_WREADY),
        .M_AXIMM_20_BRESP(M_AXIMM_20_BRESP),
        .M_AXIMM_20_BVALID(M_AXIMM_20_BVALID),
        .M_AXIMM_20_BREADY(M_AXIMM_20_BREADY),
        .M_AXIMM_20_ARADDR(M_AXIMM_20_ARADDR),
        .M_AXIMM_20_ARLEN(M_AXIMM_20_ARLEN),
        .M_AXIMM_20_ARSIZE(M_AXIMM_20_ARSIZE),
        .M_AXIMM_20_ARBURST(M_AXIMM_20_ARBURST),
        .M_AXIMM_20_ARLOCK(M_AXIMM_20_ARLOCK),
        .M_AXIMM_20_ARCACHE(M_AXIMM_20_ARCACHE),
        .M_AXIMM_20_ARPROT(M_AXIMM_20_ARPROT),
        .M_AXIMM_20_ARREGION(M_AXIMM_20_ARREGION),
        .M_AXIMM_20_ARQOS(M_AXIMM_20_ARQOS),
        .M_AXIMM_20_ARVALID(M_AXIMM_20_ARVALID),
        .M_AXIMM_20_ARREADY(M_AXIMM_20_ARREADY),
        .M_AXIMM_20_RDATA(M_AXIMM_20_RDATA),
        .M_AXIMM_20_RRESP(M_AXIMM_20_RRESP),
        .M_AXIMM_20_RLAST(M_AXIMM_20_RLAST),
        .M_AXIMM_20_RVALID(M_AXIMM_20_RVALID),
        .M_AXIMM_20_RREADY(M_AXIMM_20_RREADY),
        .AP_AXIMM_21_AWADDR(AP_AXIMM_21_AWADDR),
        .AP_AXIMM_21_AWLEN(AP_AXIMM_21_AWLEN),
        .AP_AXIMM_21_AWSIZE(AP_AXIMM_21_AWSIZE),
        .AP_AXIMM_21_AWBURST(AP_AXIMM_21_AWBURST),
        .AP_AXIMM_21_AWLOCK(AP_AXIMM_21_AWLOCK),
        .AP_AXIMM_21_AWCACHE(AP_AXIMM_21_AWCACHE),
        .AP_AXIMM_21_AWPROT(AP_AXIMM_21_AWPROT),
        .AP_AXIMM_21_AWREGION(AP_AXIMM_21_AWREGION),
        .AP_AXIMM_21_AWQOS(AP_AXIMM_21_AWQOS),
        .AP_AXIMM_21_AWVALID(AP_AXIMM_21_AWVALID),
        .AP_AXIMM_21_AWREADY(AP_AXIMM_21_AWREADY),
        .AP_AXIMM_21_WDATA(AP_AXIMM_21_WDATA),
        .AP_AXIMM_21_WSTRB(AP_AXIMM_21_WSTRB),
        .AP_AXIMM_21_WLAST(AP_AXIMM_21_WLAST),
        .AP_AXIMM_21_WVALID(AP_AXIMM_21_WVALID),
        .AP_AXIMM_21_WREADY(AP_AXIMM_21_WREADY),
        .AP_AXIMM_21_BRESP(AP_AXIMM_21_BRESP),
        .AP_AXIMM_21_BVALID(AP_AXIMM_21_BVALID),
        .AP_AXIMM_21_BREADY(AP_AXIMM_21_BREADY),
        .AP_AXIMM_21_ARADDR(AP_AXIMM_21_ARADDR),
        .AP_AXIMM_21_ARLEN(AP_AXIMM_21_ARLEN),
        .AP_AXIMM_21_ARSIZE(AP_AXIMM_21_ARSIZE),
        .AP_AXIMM_21_ARBURST(AP_AXIMM_21_ARBURST),
        .AP_AXIMM_21_ARLOCK(AP_AXIMM_21_ARLOCK),
        .AP_AXIMM_21_ARCACHE(AP_AXIMM_21_ARCACHE),
        .AP_AXIMM_21_ARPROT(AP_AXIMM_21_ARPROT),
        .AP_AXIMM_21_ARREGION(AP_AXIMM_21_ARREGION),
        .AP_AXIMM_21_ARQOS(AP_AXIMM_21_ARQOS),
        .AP_AXIMM_21_ARVALID(AP_AXIMM_21_ARVALID),
        .AP_AXIMM_21_ARREADY(AP_AXIMM_21_ARREADY),
        .AP_AXIMM_21_RDATA(AP_AXIMM_21_RDATA),
        .AP_AXIMM_21_RRESP(AP_AXIMM_21_RRESP),
        .AP_AXIMM_21_RLAST(AP_AXIMM_21_RLAST),
        .AP_AXIMM_21_RVALID(AP_AXIMM_21_RVALID),
        .AP_AXIMM_21_RREADY(AP_AXIMM_21_RREADY),
        .M_AXIMM_21_AWADDR(M_AXIMM_21_AWADDR),
        .M_AXIMM_21_AWLEN(M_AXIMM_21_AWLEN),
        .M_AXIMM_21_AWSIZE(M_AXIMM_21_AWSIZE),
        .M_AXIMM_21_AWBURST(M_AXIMM_21_AWBURST),
        .M_AXIMM_21_AWLOCK(M_AXIMM_21_AWLOCK),
        .M_AXIMM_21_AWCACHE(M_AXIMM_21_AWCACHE),
        .M_AXIMM_21_AWPROT(M_AXIMM_21_AWPROT),
        .M_AXIMM_21_AWREGION(M_AXIMM_21_AWREGION),
        .M_AXIMM_21_AWQOS(M_AXIMM_21_AWQOS),
        .M_AXIMM_21_AWVALID(M_AXIMM_21_AWVALID),
        .M_AXIMM_21_AWREADY(M_AXIMM_21_AWREADY),
        .M_AXIMM_21_WDATA(M_AXIMM_21_WDATA),
        .M_AXIMM_21_WSTRB(M_AXIMM_21_WSTRB),
        .M_AXIMM_21_WLAST(M_AXIMM_21_WLAST),
        .M_AXIMM_21_WVALID(M_AXIMM_21_WVALID),
        .M_AXIMM_21_WREADY(M_AXIMM_21_WREADY),
        .M_AXIMM_21_BRESP(M_AXIMM_21_BRESP),
        .M_AXIMM_21_BVALID(M_AXIMM_21_BVALID),
        .M_AXIMM_21_BREADY(M_AXIMM_21_BREADY),
        .M_AXIMM_21_ARADDR(M_AXIMM_21_ARADDR),
        .M_AXIMM_21_ARLEN(M_AXIMM_21_ARLEN),
        .M_AXIMM_21_ARSIZE(M_AXIMM_21_ARSIZE),
        .M_AXIMM_21_ARBURST(M_AXIMM_21_ARBURST),
        .M_AXIMM_21_ARLOCK(M_AXIMM_21_ARLOCK),
        .M_AXIMM_21_ARCACHE(M_AXIMM_21_ARCACHE),
        .M_AXIMM_21_ARPROT(M_AXIMM_21_ARPROT),
        .M_AXIMM_21_ARREGION(M_AXIMM_21_ARREGION),
        .M_AXIMM_21_ARQOS(M_AXIMM_21_ARQOS),
        .M_AXIMM_21_ARVALID(M_AXIMM_21_ARVALID),
        .M_AXIMM_21_ARREADY(M_AXIMM_21_ARREADY),
        .M_AXIMM_21_RDATA(M_AXIMM_21_RDATA),
        .M_AXIMM_21_RRESP(M_AXIMM_21_RRESP),
        .M_AXIMM_21_RLAST(M_AXIMM_21_RLAST),
        .M_AXIMM_21_RVALID(M_AXIMM_21_RVALID),
        .M_AXIMM_21_RREADY(M_AXIMM_21_RREADY),
        .AP_AXIMM_22_AWADDR(AP_AXIMM_22_AWADDR),
        .AP_AXIMM_22_AWLEN(AP_AXIMM_22_AWLEN),
        .AP_AXIMM_22_AWSIZE(AP_AXIMM_22_AWSIZE),
        .AP_AXIMM_22_AWBURST(AP_AXIMM_22_AWBURST),
        .AP_AXIMM_22_AWLOCK(AP_AXIMM_22_AWLOCK),
        .AP_AXIMM_22_AWCACHE(AP_AXIMM_22_AWCACHE),
        .AP_AXIMM_22_AWPROT(AP_AXIMM_22_AWPROT),
        .AP_AXIMM_22_AWREGION(AP_AXIMM_22_AWREGION),
        .AP_AXIMM_22_AWQOS(AP_AXIMM_22_AWQOS),
        .AP_AXIMM_22_AWVALID(AP_AXIMM_22_AWVALID),
        .AP_AXIMM_22_AWREADY(AP_AXIMM_22_AWREADY),
        .AP_AXIMM_22_WDATA(AP_AXIMM_22_WDATA),
        .AP_AXIMM_22_WSTRB(AP_AXIMM_22_WSTRB),
        .AP_AXIMM_22_WLAST(AP_AXIMM_22_WLAST),
        .AP_AXIMM_22_WVALID(AP_AXIMM_22_WVALID),
        .AP_AXIMM_22_WREADY(AP_AXIMM_22_WREADY),
        .AP_AXIMM_22_BRESP(AP_AXIMM_22_BRESP),
        .AP_AXIMM_22_BVALID(AP_AXIMM_22_BVALID),
        .AP_AXIMM_22_BREADY(AP_AXIMM_22_BREADY),
        .AP_AXIMM_22_ARADDR(AP_AXIMM_22_ARADDR),
        .AP_AXIMM_22_ARLEN(AP_AXIMM_22_ARLEN),
        .AP_AXIMM_22_ARSIZE(AP_AXIMM_22_ARSIZE),
        .AP_AXIMM_22_ARBURST(AP_AXIMM_22_ARBURST),
        .AP_AXIMM_22_ARLOCK(AP_AXIMM_22_ARLOCK),
        .AP_AXIMM_22_ARCACHE(AP_AXIMM_22_ARCACHE),
        .AP_AXIMM_22_ARPROT(AP_AXIMM_22_ARPROT),
        .AP_AXIMM_22_ARREGION(AP_AXIMM_22_ARREGION),
        .AP_AXIMM_22_ARQOS(AP_AXIMM_22_ARQOS),
        .AP_AXIMM_22_ARVALID(AP_AXIMM_22_ARVALID),
        .AP_AXIMM_22_ARREADY(AP_AXIMM_22_ARREADY),
        .AP_AXIMM_22_RDATA(AP_AXIMM_22_RDATA),
        .AP_AXIMM_22_RRESP(AP_AXIMM_22_RRESP),
        .AP_AXIMM_22_RLAST(AP_AXIMM_22_RLAST),
        .AP_AXIMM_22_RVALID(AP_AXIMM_22_RVALID),
        .AP_AXIMM_22_RREADY(AP_AXIMM_22_RREADY),
        .M_AXIMM_22_AWADDR(M_AXIMM_22_AWADDR),
        .M_AXIMM_22_AWLEN(M_AXIMM_22_AWLEN),
        .M_AXIMM_22_AWSIZE(M_AXIMM_22_AWSIZE),
        .M_AXIMM_22_AWBURST(M_AXIMM_22_AWBURST),
        .M_AXIMM_22_AWLOCK(M_AXIMM_22_AWLOCK),
        .M_AXIMM_22_AWCACHE(M_AXIMM_22_AWCACHE),
        .M_AXIMM_22_AWPROT(M_AXIMM_22_AWPROT),
        .M_AXIMM_22_AWREGION(M_AXIMM_22_AWREGION),
        .M_AXIMM_22_AWQOS(M_AXIMM_22_AWQOS),
        .M_AXIMM_22_AWVALID(M_AXIMM_22_AWVALID),
        .M_AXIMM_22_AWREADY(M_AXIMM_22_AWREADY),
        .M_AXIMM_22_WDATA(M_AXIMM_22_WDATA),
        .M_AXIMM_22_WSTRB(M_AXIMM_22_WSTRB),
        .M_AXIMM_22_WLAST(M_AXIMM_22_WLAST),
        .M_AXIMM_22_WVALID(M_AXIMM_22_WVALID),
        .M_AXIMM_22_WREADY(M_AXIMM_22_WREADY),
        .M_AXIMM_22_BRESP(M_AXIMM_22_BRESP),
        .M_AXIMM_22_BVALID(M_AXIMM_22_BVALID),
        .M_AXIMM_22_BREADY(M_AXIMM_22_BREADY),
        .M_AXIMM_22_ARADDR(M_AXIMM_22_ARADDR),
        .M_AXIMM_22_ARLEN(M_AXIMM_22_ARLEN),
        .M_AXIMM_22_ARSIZE(M_AXIMM_22_ARSIZE),
        .M_AXIMM_22_ARBURST(M_AXIMM_22_ARBURST),
        .M_AXIMM_22_ARLOCK(M_AXIMM_22_ARLOCK),
        .M_AXIMM_22_ARCACHE(M_AXIMM_22_ARCACHE),
        .M_AXIMM_22_ARPROT(M_AXIMM_22_ARPROT),
        .M_AXIMM_22_ARREGION(M_AXIMM_22_ARREGION),
        .M_AXIMM_22_ARQOS(M_AXIMM_22_ARQOS),
        .M_AXIMM_22_ARVALID(M_AXIMM_22_ARVALID),
        .M_AXIMM_22_ARREADY(M_AXIMM_22_ARREADY),
        .M_AXIMM_22_RDATA(M_AXIMM_22_RDATA),
        .M_AXIMM_22_RRESP(M_AXIMM_22_RRESP),
        .M_AXIMM_22_RLAST(M_AXIMM_22_RLAST),
        .M_AXIMM_22_RVALID(M_AXIMM_22_RVALID),
        .M_AXIMM_22_RREADY(M_AXIMM_22_RREADY),
        .AP_AXIMM_23_AWADDR(AP_AXIMM_23_AWADDR),
        .AP_AXIMM_23_AWLEN(AP_AXIMM_23_AWLEN),
        .AP_AXIMM_23_AWSIZE(AP_AXIMM_23_AWSIZE),
        .AP_AXIMM_23_AWBURST(AP_AXIMM_23_AWBURST),
        .AP_AXIMM_23_AWLOCK(AP_AXIMM_23_AWLOCK),
        .AP_AXIMM_23_AWCACHE(AP_AXIMM_23_AWCACHE),
        .AP_AXIMM_23_AWPROT(AP_AXIMM_23_AWPROT),
        .AP_AXIMM_23_AWREGION(AP_AXIMM_23_AWREGION),
        .AP_AXIMM_23_AWQOS(AP_AXIMM_23_AWQOS),
        .AP_AXIMM_23_AWVALID(AP_AXIMM_23_AWVALID),
        .AP_AXIMM_23_AWREADY(AP_AXIMM_23_AWREADY),
        .AP_AXIMM_23_WDATA(AP_AXIMM_23_WDATA),
        .AP_AXIMM_23_WSTRB(AP_AXIMM_23_WSTRB),
        .AP_AXIMM_23_WLAST(AP_AXIMM_23_WLAST),
        .AP_AXIMM_23_WVALID(AP_AXIMM_23_WVALID),
        .AP_AXIMM_23_WREADY(AP_AXIMM_23_WREADY),
        .AP_AXIMM_23_BRESP(AP_AXIMM_23_BRESP),
        .AP_AXIMM_23_BVALID(AP_AXIMM_23_BVALID),
        .AP_AXIMM_23_BREADY(AP_AXIMM_23_BREADY),
        .AP_AXIMM_23_ARADDR(AP_AXIMM_23_ARADDR),
        .AP_AXIMM_23_ARLEN(AP_AXIMM_23_ARLEN),
        .AP_AXIMM_23_ARSIZE(AP_AXIMM_23_ARSIZE),
        .AP_AXIMM_23_ARBURST(AP_AXIMM_23_ARBURST),
        .AP_AXIMM_23_ARLOCK(AP_AXIMM_23_ARLOCK),
        .AP_AXIMM_23_ARCACHE(AP_AXIMM_23_ARCACHE),
        .AP_AXIMM_23_ARPROT(AP_AXIMM_23_ARPROT),
        .AP_AXIMM_23_ARREGION(AP_AXIMM_23_ARREGION),
        .AP_AXIMM_23_ARQOS(AP_AXIMM_23_ARQOS),
        .AP_AXIMM_23_ARVALID(AP_AXIMM_23_ARVALID),
        .AP_AXIMM_23_ARREADY(AP_AXIMM_23_ARREADY),
        .AP_AXIMM_23_RDATA(AP_AXIMM_23_RDATA),
        .AP_AXIMM_23_RRESP(AP_AXIMM_23_RRESP),
        .AP_AXIMM_23_RLAST(AP_AXIMM_23_RLAST),
        .AP_AXIMM_23_RVALID(AP_AXIMM_23_RVALID),
        .AP_AXIMM_23_RREADY(AP_AXIMM_23_RREADY),
        .M_AXIMM_23_AWADDR(M_AXIMM_23_AWADDR),
        .M_AXIMM_23_AWLEN(M_AXIMM_23_AWLEN),
        .M_AXIMM_23_AWSIZE(M_AXIMM_23_AWSIZE),
        .M_AXIMM_23_AWBURST(M_AXIMM_23_AWBURST),
        .M_AXIMM_23_AWLOCK(M_AXIMM_23_AWLOCK),
        .M_AXIMM_23_AWCACHE(M_AXIMM_23_AWCACHE),
        .M_AXIMM_23_AWPROT(M_AXIMM_23_AWPROT),
        .M_AXIMM_23_AWREGION(M_AXIMM_23_AWREGION),
        .M_AXIMM_23_AWQOS(M_AXIMM_23_AWQOS),
        .M_AXIMM_23_AWVALID(M_AXIMM_23_AWVALID),
        .M_AXIMM_23_AWREADY(M_AXIMM_23_AWREADY),
        .M_AXIMM_23_WDATA(M_AXIMM_23_WDATA),
        .M_AXIMM_23_WSTRB(M_AXIMM_23_WSTRB),
        .M_AXIMM_23_WLAST(M_AXIMM_23_WLAST),
        .M_AXIMM_23_WVALID(M_AXIMM_23_WVALID),
        .M_AXIMM_23_WREADY(M_AXIMM_23_WREADY),
        .M_AXIMM_23_BRESP(M_AXIMM_23_BRESP),
        .M_AXIMM_23_BVALID(M_AXIMM_23_BVALID),
        .M_AXIMM_23_BREADY(M_AXIMM_23_BREADY),
        .M_AXIMM_23_ARADDR(M_AXIMM_23_ARADDR),
        .M_AXIMM_23_ARLEN(M_AXIMM_23_ARLEN),
        .M_AXIMM_23_ARSIZE(M_AXIMM_23_ARSIZE),
        .M_AXIMM_23_ARBURST(M_AXIMM_23_ARBURST),
        .M_AXIMM_23_ARLOCK(M_AXIMM_23_ARLOCK),
        .M_AXIMM_23_ARCACHE(M_AXIMM_23_ARCACHE),
        .M_AXIMM_23_ARPROT(M_AXIMM_23_ARPROT),
        .M_AXIMM_23_ARREGION(M_AXIMM_23_ARREGION),
        .M_AXIMM_23_ARQOS(M_AXIMM_23_ARQOS),
        .M_AXIMM_23_ARVALID(M_AXIMM_23_ARVALID),
        .M_AXIMM_23_ARREADY(M_AXIMM_23_ARREADY),
        .M_AXIMM_23_RDATA(M_AXIMM_23_RDATA),
        .M_AXIMM_23_RRESP(M_AXIMM_23_RRESP),
        .M_AXIMM_23_RLAST(M_AXIMM_23_RLAST),
        .M_AXIMM_23_RVALID(M_AXIMM_23_RVALID),
        .M_AXIMM_23_RREADY(M_AXIMM_23_RREADY),
        .AP_AXIMM_24_AWADDR(AP_AXIMM_24_AWADDR),
        .AP_AXIMM_24_AWLEN(AP_AXIMM_24_AWLEN),
        .AP_AXIMM_24_AWSIZE(AP_AXIMM_24_AWSIZE),
        .AP_AXIMM_24_AWBURST(AP_AXIMM_24_AWBURST),
        .AP_AXIMM_24_AWLOCK(AP_AXIMM_24_AWLOCK),
        .AP_AXIMM_24_AWCACHE(AP_AXIMM_24_AWCACHE),
        .AP_AXIMM_24_AWPROT(AP_AXIMM_24_AWPROT),
        .AP_AXIMM_24_AWREGION(AP_AXIMM_24_AWREGION),
        .AP_AXIMM_24_AWQOS(AP_AXIMM_24_AWQOS),
        .AP_AXIMM_24_AWVALID(AP_AXIMM_24_AWVALID),
        .AP_AXIMM_24_AWREADY(AP_AXIMM_24_AWREADY),
        .AP_AXIMM_24_WDATA(AP_AXIMM_24_WDATA),
        .AP_AXIMM_24_WSTRB(AP_AXIMM_24_WSTRB),
        .AP_AXIMM_24_WLAST(AP_AXIMM_24_WLAST),
        .AP_AXIMM_24_WVALID(AP_AXIMM_24_WVALID),
        .AP_AXIMM_24_WREADY(AP_AXIMM_24_WREADY),
        .AP_AXIMM_24_BRESP(AP_AXIMM_24_BRESP),
        .AP_AXIMM_24_BVALID(AP_AXIMM_24_BVALID),
        .AP_AXIMM_24_BREADY(AP_AXIMM_24_BREADY),
        .AP_AXIMM_24_ARADDR(AP_AXIMM_24_ARADDR),
        .AP_AXIMM_24_ARLEN(AP_AXIMM_24_ARLEN),
        .AP_AXIMM_24_ARSIZE(AP_AXIMM_24_ARSIZE),
        .AP_AXIMM_24_ARBURST(AP_AXIMM_24_ARBURST),
        .AP_AXIMM_24_ARLOCK(AP_AXIMM_24_ARLOCK),
        .AP_AXIMM_24_ARCACHE(AP_AXIMM_24_ARCACHE),
        .AP_AXIMM_24_ARPROT(AP_AXIMM_24_ARPROT),
        .AP_AXIMM_24_ARREGION(AP_AXIMM_24_ARREGION),
        .AP_AXIMM_24_ARQOS(AP_AXIMM_24_ARQOS),
        .AP_AXIMM_24_ARVALID(AP_AXIMM_24_ARVALID),
        .AP_AXIMM_24_ARREADY(AP_AXIMM_24_ARREADY),
        .AP_AXIMM_24_RDATA(AP_AXIMM_24_RDATA),
        .AP_AXIMM_24_RRESP(AP_AXIMM_24_RRESP),
        .AP_AXIMM_24_RLAST(AP_AXIMM_24_RLAST),
        .AP_AXIMM_24_RVALID(AP_AXIMM_24_RVALID),
        .AP_AXIMM_24_RREADY(AP_AXIMM_24_RREADY),
        .M_AXIMM_24_AWADDR(M_AXIMM_24_AWADDR),
        .M_AXIMM_24_AWLEN(M_AXIMM_24_AWLEN),
        .M_AXIMM_24_AWSIZE(M_AXIMM_24_AWSIZE),
        .M_AXIMM_24_AWBURST(M_AXIMM_24_AWBURST),
        .M_AXIMM_24_AWLOCK(M_AXIMM_24_AWLOCK),
        .M_AXIMM_24_AWCACHE(M_AXIMM_24_AWCACHE),
        .M_AXIMM_24_AWPROT(M_AXIMM_24_AWPROT),
        .M_AXIMM_24_AWREGION(M_AXIMM_24_AWREGION),
        .M_AXIMM_24_AWQOS(M_AXIMM_24_AWQOS),
        .M_AXIMM_24_AWVALID(M_AXIMM_24_AWVALID),
        .M_AXIMM_24_AWREADY(M_AXIMM_24_AWREADY),
        .M_AXIMM_24_WDATA(M_AXIMM_24_WDATA),
        .M_AXIMM_24_WSTRB(M_AXIMM_24_WSTRB),
        .M_AXIMM_24_WLAST(M_AXIMM_24_WLAST),
        .M_AXIMM_24_WVALID(M_AXIMM_24_WVALID),
        .M_AXIMM_24_WREADY(M_AXIMM_24_WREADY),
        .M_AXIMM_24_BRESP(M_AXIMM_24_BRESP),
        .M_AXIMM_24_BVALID(M_AXIMM_24_BVALID),
        .M_AXIMM_24_BREADY(M_AXIMM_24_BREADY),
        .M_AXIMM_24_ARADDR(M_AXIMM_24_ARADDR),
        .M_AXIMM_24_ARLEN(M_AXIMM_24_ARLEN),
        .M_AXIMM_24_ARSIZE(M_AXIMM_24_ARSIZE),
        .M_AXIMM_24_ARBURST(M_AXIMM_24_ARBURST),
        .M_AXIMM_24_ARLOCK(M_AXIMM_24_ARLOCK),
        .M_AXIMM_24_ARCACHE(M_AXIMM_24_ARCACHE),
        .M_AXIMM_24_ARPROT(M_AXIMM_24_ARPROT),
        .M_AXIMM_24_ARREGION(M_AXIMM_24_ARREGION),
        .M_AXIMM_24_ARQOS(M_AXIMM_24_ARQOS),
        .M_AXIMM_24_ARVALID(M_AXIMM_24_ARVALID),
        .M_AXIMM_24_ARREADY(M_AXIMM_24_ARREADY),
        .M_AXIMM_24_RDATA(M_AXIMM_24_RDATA),
        .M_AXIMM_24_RRESP(M_AXIMM_24_RRESP),
        .M_AXIMM_24_RLAST(M_AXIMM_24_RLAST),
        .M_AXIMM_24_RVALID(M_AXIMM_24_RVALID),
        .M_AXIMM_24_RREADY(M_AXIMM_24_RREADY),
        .AP_AXIMM_25_AWADDR(AP_AXIMM_25_AWADDR),
        .AP_AXIMM_25_AWLEN(AP_AXIMM_25_AWLEN),
        .AP_AXIMM_25_AWSIZE(AP_AXIMM_25_AWSIZE),
        .AP_AXIMM_25_AWBURST(AP_AXIMM_25_AWBURST),
        .AP_AXIMM_25_AWLOCK(AP_AXIMM_25_AWLOCK),
        .AP_AXIMM_25_AWCACHE(AP_AXIMM_25_AWCACHE),
        .AP_AXIMM_25_AWPROT(AP_AXIMM_25_AWPROT),
        .AP_AXIMM_25_AWREGION(AP_AXIMM_25_AWREGION),
        .AP_AXIMM_25_AWQOS(AP_AXIMM_25_AWQOS),
        .AP_AXIMM_25_AWVALID(AP_AXIMM_25_AWVALID),
        .AP_AXIMM_25_AWREADY(AP_AXIMM_25_AWREADY),
        .AP_AXIMM_25_WDATA(AP_AXIMM_25_WDATA),
        .AP_AXIMM_25_WSTRB(AP_AXIMM_25_WSTRB),
        .AP_AXIMM_25_WLAST(AP_AXIMM_25_WLAST),
        .AP_AXIMM_25_WVALID(AP_AXIMM_25_WVALID),
        .AP_AXIMM_25_WREADY(AP_AXIMM_25_WREADY),
        .AP_AXIMM_25_BRESP(AP_AXIMM_25_BRESP),
        .AP_AXIMM_25_BVALID(AP_AXIMM_25_BVALID),
        .AP_AXIMM_25_BREADY(AP_AXIMM_25_BREADY),
        .AP_AXIMM_25_ARADDR(AP_AXIMM_25_ARADDR),
        .AP_AXIMM_25_ARLEN(AP_AXIMM_25_ARLEN),
        .AP_AXIMM_25_ARSIZE(AP_AXIMM_25_ARSIZE),
        .AP_AXIMM_25_ARBURST(AP_AXIMM_25_ARBURST),
        .AP_AXIMM_25_ARLOCK(AP_AXIMM_25_ARLOCK),
        .AP_AXIMM_25_ARCACHE(AP_AXIMM_25_ARCACHE),
        .AP_AXIMM_25_ARPROT(AP_AXIMM_25_ARPROT),
        .AP_AXIMM_25_ARREGION(AP_AXIMM_25_ARREGION),
        .AP_AXIMM_25_ARQOS(AP_AXIMM_25_ARQOS),
        .AP_AXIMM_25_ARVALID(AP_AXIMM_25_ARVALID),
        .AP_AXIMM_25_ARREADY(AP_AXIMM_25_ARREADY),
        .AP_AXIMM_25_RDATA(AP_AXIMM_25_RDATA),
        .AP_AXIMM_25_RRESP(AP_AXIMM_25_RRESP),
        .AP_AXIMM_25_RLAST(AP_AXIMM_25_RLAST),
        .AP_AXIMM_25_RVALID(AP_AXIMM_25_RVALID),
        .AP_AXIMM_25_RREADY(AP_AXIMM_25_RREADY),
        .M_AXIMM_25_AWADDR(M_AXIMM_25_AWADDR),
        .M_AXIMM_25_AWLEN(M_AXIMM_25_AWLEN),
        .M_AXIMM_25_AWSIZE(M_AXIMM_25_AWSIZE),
        .M_AXIMM_25_AWBURST(M_AXIMM_25_AWBURST),
        .M_AXIMM_25_AWLOCK(M_AXIMM_25_AWLOCK),
        .M_AXIMM_25_AWCACHE(M_AXIMM_25_AWCACHE),
        .M_AXIMM_25_AWPROT(M_AXIMM_25_AWPROT),
        .M_AXIMM_25_AWREGION(M_AXIMM_25_AWREGION),
        .M_AXIMM_25_AWQOS(M_AXIMM_25_AWQOS),
        .M_AXIMM_25_AWVALID(M_AXIMM_25_AWVALID),
        .M_AXIMM_25_AWREADY(M_AXIMM_25_AWREADY),
        .M_AXIMM_25_WDATA(M_AXIMM_25_WDATA),
        .M_AXIMM_25_WSTRB(M_AXIMM_25_WSTRB),
        .M_AXIMM_25_WLAST(M_AXIMM_25_WLAST),
        .M_AXIMM_25_WVALID(M_AXIMM_25_WVALID),
        .M_AXIMM_25_WREADY(M_AXIMM_25_WREADY),
        .M_AXIMM_25_BRESP(M_AXIMM_25_BRESP),
        .M_AXIMM_25_BVALID(M_AXIMM_25_BVALID),
        .M_AXIMM_25_BREADY(M_AXIMM_25_BREADY),
        .M_AXIMM_25_ARADDR(M_AXIMM_25_ARADDR),
        .M_AXIMM_25_ARLEN(M_AXIMM_25_ARLEN),
        .M_AXIMM_25_ARSIZE(M_AXIMM_25_ARSIZE),
        .M_AXIMM_25_ARBURST(M_AXIMM_25_ARBURST),
        .M_AXIMM_25_ARLOCK(M_AXIMM_25_ARLOCK),
        .M_AXIMM_25_ARCACHE(M_AXIMM_25_ARCACHE),
        .M_AXIMM_25_ARPROT(M_AXIMM_25_ARPROT),
        .M_AXIMM_25_ARREGION(M_AXIMM_25_ARREGION),
        .M_AXIMM_25_ARQOS(M_AXIMM_25_ARQOS),
        .M_AXIMM_25_ARVALID(M_AXIMM_25_ARVALID),
        .M_AXIMM_25_ARREADY(M_AXIMM_25_ARREADY),
        .M_AXIMM_25_RDATA(M_AXIMM_25_RDATA),
        .M_AXIMM_25_RRESP(M_AXIMM_25_RRESP),
        .M_AXIMM_25_RLAST(M_AXIMM_25_RLAST),
        .M_AXIMM_25_RVALID(M_AXIMM_25_RVALID),
        .M_AXIMM_25_RREADY(M_AXIMM_25_RREADY),
        .AP_AXIMM_26_AWADDR(AP_AXIMM_26_AWADDR),
        .AP_AXIMM_26_AWLEN(AP_AXIMM_26_AWLEN),
        .AP_AXIMM_26_AWSIZE(AP_AXIMM_26_AWSIZE),
        .AP_AXIMM_26_AWBURST(AP_AXIMM_26_AWBURST),
        .AP_AXIMM_26_AWLOCK(AP_AXIMM_26_AWLOCK),
        .AP_AXIMM_26_AWCACHE(AP_AXIMM_26_AWCACHE),
        .AP_AXIMM_26_AWPROT(AP_AXIMM_26_AWPROT),
        .AP_AXIMM_26_AWREGION(AP_AXIMM_26_AWREGION),
        .AP_AXIMM_26_AWQOS(AP_AXIMM_26_AWQOS),
        .AP_AXIMM_26_AWVALID(AP_AXIMM_26_AWVALID),
        .AP_AXIMM_26_AWREADY(AP_AXIMM_26_AWREADY),
        .AP_AXIMM_26_WDATA(AP_AXIMM_26_WDATA),
        .AP_AXIMM_26_WSTRB(AP_AXIMM_26_WSTRB),
        .AP_AXIMM_26_WLAST(AP_AXIMM_26_WLAST),
        .AP_AXIMM_26_WVALID(AP_AXIMM_26_WVALID),
        .AP_AXIMM_26_WREADY(AP_AXIMM_26_WREADY),
        .AP_AXIMM_26_BRESP(AP_AXIMM_26_BRESP),
        .AP_AXIMM_26_BVALID(AP_AXIMM_26_BVALID),
        .AP_AXIMM_26_BREADY(AP_AXIMM_26_BREADY),
        .AP_AXIMM_26_ARADDR(AP_AXIMM_26_ARADDR),
        .AP_AXIMM_26_ARLEN(AP_AXIMM_26_ARLEN),
        .AP_AXIMM_26_ARSIZE(AP_AXIMM_26_ARSIZE),
        .AP_AXIMM_26_ARBURST(AP_AXIMM_26_ARBURST),
        .AP_AXIMM_26_ARLOCK(AP_AXIMM_26_ARLOCK),
        .AP_AXIMM_26_ARCACHE(AP_AXIMM_26_ARCACHE),
        .AP_AXIMM_26_ARPROT(AP_AXIMM_26_ARPROT),
        .AP_AXIMM_26_ARREGION(AP_AXIMM_26_ARREGION),
        .AP_AXIMM_26_ARQOS(AP_AXIMM_26_ARQOS),
        .AP_AXIMM_26_ARVALID(AP_AXIMM_26_ARVALID),
        .AP_AXIMM_26_ARREADY(AP_AXIMM_26_ARREADY),
        .AP_AXIMM_26_RDATA(AP_AXIMM_26_RDATA),
        .AP_AXIMM_26_RRESP(AP_AXIMM_26_RRESP),
        .AP_AXIMM_26_RLAST(AP_AXIMM_26_RLAST),
        .AP_AXIMM_26_RVALID(AP_AXIMM_26_RVALID),
        .AP_AXIMM_26_RREADY(AP_AXIMM_26_RREADY),
        .M_AXIMM_26_AWADDR(M_AXIMM_26_AWADDR),
        .M_AXIMM_26_AWLEN(M_AXIMM_26_AWLEN),
        .M_AXIMM_26_AWSIZE(M_AXIMM_26_AWSIZE),
        .M_AXIMM_26_AWBURST(M_AXIMM_26_AWBURST),
        .M_AXIMM_26_AWLOCK(M_AXIMM_26_AWLOCK),
        .M_AXIMM_26_AWCACHE(M_AXIMM_26_AWCACHE),
        .M_AXIMM_26_AWPROT(M_AXIMM_26_AWPROT),
        .M_AXIMM_26_AWREGION(M_AXIMM_26_AWREGION),
        .M_AXIMM_26_AWQOS(M_AXIMM_26_AWQOS),
        .M_AXIMM_26_AWVALID(M_AXIMM_26_AWVALID),
        .M_AXIMM_26_AWREADY(M_AXIMM_26_AWREADY),
        .M_AXIMM_26_WDATA(M_AXIMM_26_WDATA),
        .M_AXIMM_26_WSTRB(M_AXIMM_26_WSTRB),
        .M_AXIMM_26_WLAST(M_AXIMM_26_WLAST),
        .M_AXIMM_26_WVALID(M_AXIMM_26_WVALID),
        .M_AXIMM_26_WREADY(M_AXIMM_26_WREADY),
        .M_AXIMM_26_BRESP(M_AXIMM_26_BRESP),
        .M_AXIMM_26_BVALID(M_AXIMM_26_BVALID),
        .M_AXIMM_26_BREADY(M_AXIMM_26_BREADY),
        .M_AXIMM_26_ARADDR(M_AXIMM_26_ARADDR),
        .M_AXIMM_26_ARLEN(M_AXIMM_26_ARLEN),
        .M_AXIMM_26_ARSIZE(M_AXIMM_26_ARSIZE),
        .M_AXIMM_26_ARBURST(M_AXIMM_26_ARBURST),
        .M_AXIMM_26_ARLOCK(M_AXIMM_26_ARLOCK),
        .M_AXIMM_26_ARCACHE(M_AXIMM_26_ARCACHE),
        .M_AXIMM_26_ARPROT(M_AXIMM_26_ARPROT),
        .M_AXIMM_26_ARREGION(M_AXIMM_26_ARREGION),
        .M_AXIMM_26_ARQOS(M_AXIMM_26_ARQOS),
        .M_AXIMM_26_ARVALID(M_AXIMM_26_ARVALID),
        .M_AXIMM_26_ARREADY(M_AXIMM_26_ARREADY),
        .M_AXIMM_26_RDATA(M_AXIMM_26_RDATA),
        .M_AXIMM_26_RRESP(M_AXIMM_26_RRESP),
        .M_AXIMM_26_RLAST(M_AXIMM_26_RLAST),
        .M_AXIMM_26_RVALID(M_AXIMM_26_RVALID),
        .M_AXIMM_26_RREADY(M_AXIMM_26_RREADY),
        .AP_AXIMM_27_AWADDR(AP_AXIMM_27_AWADDR),
        .AP_AXIMM_27_AWLEN(AP_AXIMM_27_AWLEN),
        .AP_AXIMM_27_AWSIZE(AP_AXIMM_27_AWSIZE),
        .AP_AXIMM_27_AWBURST(AP_AXIMM_27_AWBURST),
        .AP_AXIMM_27_AWLOCK(AP_AXIMM_27_AWLOCK),
        .AP_AXIMM_27_AWCACHE(AP_AXIMM_27_AWCACHE),
        .AP_AXIMM_27_AWPROT(AP_AXIMM_27_AWPROT),
        .AP_AXIMM_27_AWREGION(AP_AXIMM_27_AWREGION),
        .AP_AXIMM_27_AWQOS(AP_AXIMM_27_AWQOS),
        .AP_AXIMM_27_AWVALID(AP_AXIMM_27_AWVALID),
        .AP_AXIMM_27_AWREADY(AP_AXIMM_27_AWREADY),
        .AP_AXIMM_27_WDATA(AP_AXIMM_27_WDATA),
        .AP_AXIMM_27_WSTRB(AP_AXIMM_27_WSTRB),
        .AP_AXIMM_27_WLAST(AP_AXIMM_27_WLAST),
        .AP_AXIMM_27_WVALID(AP_AXIMM_27_WVALID),
        .AP_AXIMM_27_WREADY(AP_AXIMM_27_WREADY),
        .AP_AXIMM_27_BRESP(AP_AXIMM_27_BRESP),
        .AP_AXIMM_27_BVALID(AP_AXIMM_27_BVALID),
        .AP_AXIMM_27_BREADY(AP_AXIMM_27_BREADY),
        .AP_AXIMM_27_ARADDR(AP_AXIMM_27_ARADDR),
        .AP_AXIMM_27_ARLEN(AP_AXIMM_27_ARLEN),
        .AP_AXIMM_27_ARSIZE(AP_AXIMM_27_ARSIZE),
        .AP_AXIMM_27_ARBURST(AP_AXIMM_27_ARBURST),
        .AP_AXIMM_27_ARLOCK(AP_AXIMM_27_ARLOCK),
        .AP_AXIMM_27_ARCACHE(AP_AXIMM_27_ARCACHE),
        .AP_AXIMM_27_ARPROT(AP_AXIMM_27_ARPROT),
        .AP_AXIMM_27_ARREGION(AP_AXIMM_27_ARREGION),
        .AP_AXIMM_27_ARQOS(AP_AXIMM_27_ARQOS),
        .AP_AXIMM_27_ARVALID(AP_AXIMM_27_ARVALID),
        .AP_AXIMM_27_ARREADY(AP_AXIMM_27_ARREADY),
        .AP_AXIMM_27_RDATA(AP_AXIMM_27_RDATA),
        .AP_AXIMM_27_RRESP(AP_AXIMM_27_RRESP),
        .AP_AXIMM_27_RLAST(AP_AXIMM_27_RLAST),
        .AP_AXIMM_27_RVALID(AP_AXIMM_27_RVALID),
        .AP_AXIMM_27_RREADY(AP_AXIMM_27_RREADY),
        .M_AXIMM_27_AWADDR(M_AXIMM_27_AWADDR),
        .M_AXIMM_27_AWLEN(M_AXIMM_27_AWLEN),
        .M_AXIMM_27_AWSIZE(M_AXIMM_27_AWSIZE),
        .M_AXIMM_27_AWBURST(M_AXIMM_27_AWBURST),
        .M_AXIMM_27_AWLOCK(M_AXIMM_27_AWLOCK),
        .M_AXIMM_27_AWCACHE(M_AXIMM_27_AWCACHE),
        .M_AXIMM_27_AWPROT(M_AXIMM_27_AWPROT),
        .M_AXIMM_27_AWREGION(M_AXIMM_27_AWREGION),
        .M_AXIMM_27_AWQOS(M_AXIMM_27_AWQOS),
        .M_AXIMM_27_AWVALID(M_AXIMM_27_AWVALID),
        .M_AXIMM_27_AWREADY(M_AXIMM_27_AWREADY),
        .M_AXIMM_27_WDATA(M_AXIMM_27_WDATA),
        .M_AXIMM_27_WSTRB(M_AXIMM_27_WSTRB),
        .M_AXIMM_27_WLAST(M_AXIMM_27_WLAST),
        .M_AXIMM_27_WVALID(M_AXIMM_27_WVALID),
        .M_AXIMM_27_WREADY(M_AXIMM_27_WREADY),
        .M_AXIMM_27_BRESP(M_AXIMM_27_BRESP),
        .M_AXIMM_27_BVALID(M_AXIMM_27_BVALID),
        .M_AXIMM_27_BREADY(M_AXIMM_27_BREADY),
        .M_AXIMM_27_ARADDR(M_AXIMM_27_ARADDR),
        .M_AXIMM_27_ARLEN(M_AXIMM_27_ARLEN),
        .M_AXIMM_27_ARSIZE(M_AXIMM_27_ARSIZE),
        .M_AXIMM_27_ARBURST(M_AXIMM_27_ARBURST),
        .M_AXIMM_27_ARLOCK(M_AXIMM_27_ARLOCK),
        .M_AXIMM_27_ARCACHE(M_AXIMM_27_ARCACHE),
        .M_AXIMM_27_ARPROT(M_AXIMM_27_ARPROT),
        .M_AXIMM_27_ARREGION(M_AXIMM_27_ARREGION),
        .M_AXIMM_27_ARQOS(M_AXIMM_27_ARQOS),
        .M_AXIMM_27_ARVALID(M_AXIMM_27_ARVALID),
        .M_AXIMM_27_ARREADY(M_AXIMM_27_ARREADY),
        .M_AXIMM_27_RDATA(M_AXIMM_27_RDATA),
        .M_AXIMM_27_RRESP(M_AXIMM_27_RRESP),
        .M_AXIMM_27_RLAST(M_AXIMM_27_RLAST),
        .M_AXIMM_27_RVALID(M_AXIMM_27_RVALID),
        .M_AXIMM_27_RREADY(M_AXIMM_27_RREADY),
        .AP_AXIMM_28_AWADDR(AP_AXIMM_28_AWADDR),
        .AP_AXIMM_28_AWLEN(AP_AXIMM_28_AWLEN),
        .AP_AXIMM_28_AWSIZE(AP_AXIMM_28_AWSIZE),
        .AP_AXIMM_28_AWBURST(AP_AXIMM_28_AWBURST),
        .AP_AXIMM_28_AWLOCK(AP_AXIMM_28_AWLOCK),
        .AP_AXIMM_28_AWCACHE(AP_AXIMM_28_AWCACHE),
        .AP_AXIMM_28_AWPROT(AP_AXIMM_28_AWPROT),
        .AP_AXIMM_28_AWREGION(AP_AXIMM_28_AWREGION),
        .AP_AXIMM_28_AWQOS(AP_AXIMM_28_AWQOS),
        .AP_AXIMM_28_AWVALID(AP_AXIMM_28_AWVALID),
        .AP_AXIMM_28_AWREADY(AP_AXIMM_28_AWREADY),
        .AP_AXIMM_28_WDATA(AP_AXIMM_28_WDATA),
        .AP_AXIMM_28_WSTRB(AP_AXIMM_28_WSTRB),
        .AP_AXIMM_28_WLAST(AP_AXIMM_28_WLAST),
        .AP_AXIMM_28_WVALID(AP_AXIMM_28_WVALID),
        .AP_AXIMM_28_WREADY(AP_AXIMM_28_WREADY),
        .AP_AXIMM_28_BRESP(AP_AXIMM_28_BRESP),
        .AP_AXIMM_28_BVALID(AP_AXIMM_28_BVALID),
        .AP_AXIMM_28_BREADY(AP_AXIMM_28_BREADY),
        .AP_AXIMM_28_ARADDR(AP_AXIMM_28_ARADDR),
        .AP_AXIMM_28_ARLEN(AP_AXIMM_28_ARLEN),
        .AP_AXIMM_28_ARSIZE(AP_AXIMM_28_ARSIZE),
        .AP_AXIMM_28_ARBURST(AP_AXIMM_28_ARBURST),
        .AP_AXIMM_28_ARLOCK(AP_AXIMM_28_ARLOCK),
        .AP_AXIMM_28_ARCACHE(AP_AXIMM_28_ARCACHE),
        .AP_AXIMM_28_ARPROT(AP_AXIMM_28_ARPROT),
        .AP_AXIMM_28_ARREGION(AP_AXIMM_28_ARREGION),
        .AP_AXIMM_28_ARQOS(AP_AXIMM_28_ARQOS),
        .AP_AXIMM_28_ARVALID(AP_AXIMM_28_ARVALID),
        .AP_AXIMM_28_ARREADY(AP_AXIMM_28_ARREADY),
        .AP_AXIMM_28_RDATA(AP_AXIMM_28_RDATA),
        .AP_AXIMM_28_RRESP(AP_AXIMM_28_RRESP),
        .AP_AXIMM_28_RLAST(AP_AXIMM_28_RLAST),
        .AP_AXIMM_28_RVALID(AP_AXIMM_28_RVALID),
        .AP_AXIMM_28_RREADY(AP_AXIMM_28_RREADY),
        .M_AXIMM_28_AWADDR(M_AXIMM_28_AWADDR),
        .M_AXIMM_28_AWLEN(M_AXIMM_28_AWLEN),
        .M_AXIMM_28_AWSIZE(M_AXIMM_28_AWSIZE),
        .M_AXIMM_28_AWBURST(M_AXIMM_28_AWBURST),
        .M_AXIMM_28_AWLOCK(M_AXIMM_28_AWLOCK),
        .M_AXIMM_28_AWCACHE(M_AXIMM_28_AWCACHE),
        .M_AXIMM_28_AWPROT(M_AXIMM_28_AWPROT),
        .M_AXIMM_28_AWREGION(M_AXIMM_28_AWREGION),
        .M_AXIMM_28_AWQOS(M_AXIMM_28_AWQOS),
        .M_AXIMM_28_AWVALID(M_AXIMM_28_AWVALID),
        .M_AXIMM_28_AWREADY(M_AXIMM_28_AWREADY),
        .M_AXIMM_28_WDATA(M_AXIMM_28_WDATA),
        .M_AXIMM_28_WSTRB(M_AXIMM_28_WSTRB),
        .M_AXIMM_28_WLAST(M_AXIMM_28_WLAST),
        .M_AXIMM_28_WVALID(M_AXIMM_28_WVALID),
        .M_AXIMM_28_WREADY(M_AXIMM_28_WREADY),
        .M_AXIMM_28_BRESP(M_AXIMM_28_BRESP),
        .M_AXIMM_28_BVALID(M_AXIMM_28_BVALID),
        .M_AXIMM_28_BREADY(M_AXIMM_28_BREADY),
        .M_AXIMM_28_ARADDR(M_AXIMM_28_ARADDR),
        .M_AXIMM_28_ARLEN(M_AXIMM_28_ARLEN),
        .M_AXIMM_28_ARSIZE(M_AXIMM_28_ARSIZE),
        .M_AXIMM_28_ARBURST(M_AXIMM_28_ARBURST),
        .M_AXIMM_28_ARLOCK(M_AXIMM_28_ARLOCK),
        .M_AXIMM_28_ARCACHE(M_AXIMM_28_ARCACHE),
        .M_AXIMM_28_ARPROT(M_AXIMM_28_ARPROT),
        .M_AXIMM_28_ARREGION(M_AXIMM_28_ARREGION),
        .M_AXIMM_28_ARQOS(M_AXIMM_28_ARQOS),
        .M_AXIMM_28_ARVALID(M_AXIMM_28_ARVALID),
        .M_AXIMM_28_ARREADY(M_AXIMM_28_ARREADY),
        .M_AXIMM_28_RDATA(M_AXIMM_28_RDATA),
        .M_AXIMM_28_RRESP(M_AXIMM_28_RRESP),
        .M_AXIMM_28_RLAST(M_AXIMM_28_RLAST),
        .M_AXIMM_28_RVALID(M_AXIMM_28_RVALID),
        .M_AXIMM_28_RREADY(M_AXIMM_28_RREADY),
        .AP_AXIMM_29_AWADDR(AP_AXIMM_29_AWADDR),
        .AP_AXIMM_29_AWLEN(AP_AXIMM_29_AWLEN),
        .AP_AXIMM_29_AWSIZE(AP_AXIMM_29_AWSIZE),
        .AP_AXIMM_29_AWBURST(AP_AXIMM_29_AWBURST),
        .AP_AXIMM_29_AWLOCK(AP_AXIMM_29_AWLOCK),
        .AP_AXIMM_29_AWCACHE(AP_AXIMM_29_AWCACHE),
        .AP_AXIMM_29_AWPROT(AP_AXIMM_29_AWPROT),
        .AP_AXIMM_29_AWREGION(AP_AXIMM_29_AWREGION),
        .AP_AXIMM_29_AWQOS(AP_AXIMM_29_AWQOS),
        .AP_AXIMM_29_AWVALID(AP_AXIMM_29_AWVALID),
        .AP_AXIMM_29_AWREADY(AP_AXIMM_29_AWREADY),
        .AP_AXIMM_29_WDATA(AP_AXIMM_29_WDATA),
        .AP_AXIMM_29_WSTRB(AP_AXIMM_29_WSTRB),
        .AP_AXIMM_29_WLAST(AP_AXIMM_29_WLAST),
        .AP_AXIMM_29_WVALID(AP_AXIMM_29_WVALID),
        .AP_AXIMM_29_WREADY(AP_AXIMM_29_WREADY),
        .AP_AXIMM_29_BRESP(AP_AXIMM_29_BRESP),
        .AP_AXIMM_29_BVALID(AP_AXIMM_29_BVALID),
        .AP_AXIMM_29_BREADY(AP_AXIMM_29_BREADY),
        .AP_AXIMM_29_ARADDR(AP_AXIMM_29_ARADDR),
        .AP_AXIMM_29_ARLEN(AP_AXIMM_29_ARLEN),
        .AP_AXIMM_29_ARSIZE(AP_AXIMM_29_ARSIZE),
        .AP_AXIMM_29_ARBURST(AP_AXIMM_29_ARBURST),
        .AP_AXIMM_29_ARLOCK(AP_AXIMM_29_ARLOCK),
        .AP_AXIMM_29_ARCACHE(AP_AXIMM_29_ARCACHE),
        .AP_AXIMM_29_ARPROT(AP_AXIMM_29_ARPROT),
        .AP_AXIMM_29_ARREGION(AP_AXIMM_29_ARREGION),
        .AP_AXIMM_29_ARQOS(AP_AXIMM_29_ARQOS),
        .AP_AXIMM_29_ARVALID(AP_AXIMM_29_ARVALID),
        .AP_AXIMM_29_ARREADY(AP_AXIMM_29_ARREADY),
        .AP_AXIMM_29_RDATA(AP_AXIMM_29_RDATA),
        .AP_AXIMM_29_RRESP(AP_AXIMM_29_RRESP),
        .AP_AXIMM_29_RLAST(AP_AXIMM_29_RLAST),
        .AP_AXIMM_29_RVALID(AP_AXIMM_29_RVALID),
        .AP_AXIMM_29_RREADY(AP_AXIMM_29_RREADY),
        .M_AXIMM_29_AWADDR(M_AXIMM_29_AWADDR),
        .M_AXIMM_29_AWLEN(M_AXIMM_29_AWLEN),
        .M_AXIMM_29_AWSIZE(M_AXIMM_29_AWSIZE),
        .M_AXIMM_29_AWBURST(M_AXIMM_29_AWBURST),
        .M_AXIMM_29_AWLOCK(M_AXIMM_29_AWLOCK),
        .M_AXIMM_29_AWCACHE(M_AXIMM_29_AWCACHE),
        .M_AXIMM_29_AWPROT(M_AXIMM_29_AWPROT),
        .M_AXIMM_29_AWREGION(M_AXIMM_29_AWREGION),
        .M_AXIMM_29_AWQOS(M_AXIMM_29_AWQOS),
        .M_AXIMM_29_AWVALID(M_AXIMM_29_AWVALID),
        .M_AXIMM_29_AWREADY(M_AXIMM_29_AWREADY),
        .M_AXIMM_29_WDATA(M_AXIMM_29_WDATA),
        .M_AXIMM_29_WSTRB(M_AXIMM_29_WSTRB),
        .M_AXIMM_29_WLAST(M_AXIMM_29_WLAST),
        .M_AXIMM_29_WVALID(M_AXIMM_29_WVALID),
        .M_AXIMM_29_WREADY(M_AXIMM_29_WREADY),
        .M_AXIMM_29_BRESP(M_AXIMM_29_BRESP),
        .M_AXIMM_29_BVALID(M_AXIMM_29_BVALID),
        .M_AXIMM_29_BREADY(M_AXIMM_29_BREADY),
        .M_AXIMM_29_ARADDR(M_AXIMM_29_ARADDR),
        .M_AXIMM_29_ARLEN(M_AXIMM_29_ARLEN),
        .M_AXIMM_29_ARSIZE(M_AXIMM_29_ARSIZE),
        .M_AXIMM_29_ARBURST(M_AXIMM_29_ARBURST),
        .M_AXIMM_29_ARLOCK(M_AXIMM_29_ARLOCK),
        .M_AXIMM_29_ARCACHE(M_AXIMM_29_ARCACHE),
        .M_AXIMM_29_ARPROT(M_AXIMM_29_ARPROT),
        .M_AXIMM_29_ARREGION(M_AXIMM_29_ARREGION),
        .M_AXIMM_29_ARQOS(M_AXIMM_29_ARQOS),
        .M_AXIMM_29_ARVALID(M_AXIMM_29_ARVALID),
        .M_AXIMM_29_ARREADY(M_AXIMM_29_ARREADY),
        .M_AXIMM_29_RDATA(M_AXIMM_29_RDATA),
        .M_AXIMM_29_RRESP(M_AXIMM_29_RRESP),
        .M_AXIMM_29_RLAST(M_AXIMM_29_RLAST),
        .M_AXIMM_29_RVALID(M_AXIMM_29_RVALID),
        .M_AXIMM_29_RREADY(M_AXIMM_29_RREADY),
        .AP_AXIMM_30_AWADDR(AP_AXIMM_30_AWADDR),
        .AP_AXIMM_30_AWLEN(AP_AXIMM_30_AWLEN),
        .AP_AXIMM_30_AWSIZE(AP_AXIMM_30_AWSIZE),
        .AP_AXIMM_30_AWBURST(AP_AXIMM_30_AWBURST),
        .AP_AXIMM_30_AWLOCK(AP_AXIMM_30_AWLOCK),
        .AP_AXIMM_30_AWCACHE(AP_AXIMM_30_AWCACHE),
        .AP_AXIMM_30_AWPROT(AP_AXIMM_30_AWPROT),
        .AP_AXIMM_30_AWREGION(AP_AXIMM_30_AWREGION),
        .AP_AXIMM_30_AWQOS(AP_AXIMM_30_AWQOS),
        .AP_AXIMM_30_AWVALID(AP_AXIMM_30_AWVALID),
        .AP_AXIMM_30_AWREADY(AP_AXIMM_30_AWREADY),
        .AP_AXIMM_30_WDATA(AP_AXIMM_30_WDATA),
        .AP_AXIMM_30_WSTRB(AP_AXIMM_30_WSTRB),
        .AP_AXIMM_30_WLAST(AP_AXIMM_30_WLAST),
        .AP_AXIMM_30_WVALID(AP_AXIMM_30_WVALID),
        .AP_AXIMM_30_WREADY(AP_AXIMM_30_WREADY),
        .AP_AXIMM_30_BRESP(AP_AXIMM_30_BRESP),
        .AP_AXIMM_30_BVALID(AP_AXIMM_30_BVALID),
        .AP_AXIMM_30_BREADY(AP_AXIMM_30_BREADY),
        .AP_AXIMM_30_ARADDR(AP_AXIMM_30_ARADDR),
        .AP_AXIMM_30_ARLEN(AP_AXIMM_30_ARLEN),
        .AP_AXIMM_30_ARSIZE(AP_AXIMM_30_ARSIZE),
        .AP_AXIMM_30_ARBURST(AP_AXIMM_30_ARBURST),
        .AP_AXIMM_30_ARLOCK(AP_AXIMM_30_ARLOCK),
        .AP_AXIMM_30_ARCACHE(AP_AXIMM_30_ARCACHE),
        .AP_AXIMM_30_ARPROT(AP_AXIMM_30_ARPROT),
        .AP_AXIMM_30_ARREGION(AP_AXIMM_30_ARREGION),
        .AP_AXIMM_30_ARQOS(AP_AXIMM_30_ARQOS),
        .AP_AXIMM_30_ARVALID(AP_AXIMM_30_ARVALID),
        .AP_AXIMM_30_ARREADY(AP_AXIMM_30_ARREADY),
        .AP_AXIMM_30_RDATA(AP_AXIMM_30_RDATA),
        .AP_AXIMM_30_RRESP(AP_AXIMM_30_RRESP),
        .AP_AXIMM_30_RLAST(AP_AXIMM_30_RLAST),
        .AP_AXIMM_30_RVALID(AP_AXIMM_30_RVALID),
        .AP_AXIMM_30_RREADY(AP_AXIMM_30_RREADY),
        .M_AXIMM_30_AWADDR(M_AXIMM_30_AWADDR),
        .M_AXIMM_30_AWLEN(M_AXIMM_30_AWLEN),
        .M_AXIMM_30_AWSIZE(M_AXIMM_30_AWSIZE),
        .M_AXIMM_30_AWBURST(M_AXIMM_30_AWBURST),
        .M_AXIMM_30_AWLOCK(M_AXIMM_30_AWLOCK),
        .M_AXIMM_30_AWCACHE(M_AXIMM_30_AWCACHE),
        .M_AXIMM_30_AWPROT(M_AXIMM_30_AWPROT),
        .M_AXIMM_30_AWREGION(M_AXIMM_30_AWREGION),
        .M_AXIMM_30_AWQOS(M_AXIMM_30_AWQOS),
        .M_AXIMM_30_AWVALID(M_AXIMM_30_AWVALID),
        .M_AXIMM_30_AWREADY(M_AXIMM_30_AWREADY),
        .M_AXIMM_30_WDATA(M_AXIMM_30_WDATA),
        .M_AXIMM_30_WSTRB(M_AXIMM_30_WSTRB),
        .M_AXIMM_30_WLAST(M_AXIMM_30_WLAST),
        .M_AXIMM_30_WVALID(M_AXIMM_30_WVALID),
        .M_AXIMM_30_WREADY(M_AXIMM_30_WREADY),
        .M_AXIMM_30_BRESP(M_AXIMM_30_BRESP),
        .M_AXIMM_30_BVALID(M_AXIMM_30_BVALID),
        .M_AXIMM_30_BREADY(M_AXIMM_30_BREADY),
        .M_AXIMM_30_ARADDR(M_AXIMM_30_ARADDR),
        .M_AXIMM_30_ARLEN(M_AXIMM_30_ARLEN),
        .M_AXIMM_30_ARSIZE(M_AXIMM_30_ARSIZE),
        .M_AXIMM_30_ARBURST(M_AXIMM_30_ARBURST),
        .M_AXIMM_30_ARLOCK(M_AXIMM_30_ARLOCK),
        .M_AXIMM_30_ARCACHE(M_AXIMM_30_ARCACHE),
        .M_AXIMM_30_ARPROT(M_AXIMM_30_ARPROT),
        .M_AXIMM_30_ARREGION(M_AXIMM_30_ARREGION),
        .M_AXIMM_30_ARQOS(M_AXIMM_30_ARQOS),
        .M_AXIMM_30_ARVALID(M_AXIMM_30_ARVALID),
        .M_AXIMM_30_ARREADY(M_AXIMM_30_ARREADY),
        .M_AXIMM_30_RDATA(M_AXIMM_30_RDATA),
        .M_AXIMM_30_RRESP(M_AXIMM_30_RRESP),
        .M_AXIMM_30_RLAST(M_AXIMM_30_RLAST),
        .M_AXIMM_30_RVALID(M_AXIMM_30_RVALID),
        .M_AXIMM_30_RREADY(M_AXIMM_30_RREADY),
        .AP_AXIMM_31_AWADDR(AP_AXIMM_31_AWADDR),
        .AP_AXIMM_31_AWLEN(AP_AXIMM_31_AWLEN),
        .AP_AXIMM_31_AWSIZE(AP_AXIMM_31_AWSIZE),
        .AP_AXIMM_31_AWBURST(AP_AXIMM_31_AWBURST),
        .AP_AXIMM_31_AWLOCK(AP_AXIMM_31_AWLOCK),
        .AP_AXIMM_31_AWCACHE(AP_AXIMM_31_AWCACHE),
        .AP_AXIMM_31_AWPROT(AP_AXIMM_31_AWPROT),
        .AP_AXIMM_31_AWREGION(AP_AXIMM_31_AWREGION),
        .AP_AXIMM_31_AWQOS(AP_AXIMM_31_AWQOS),
        .AP_AXIMM_31_AWVALID(AP_AXIMM_31_AWVALID),
        .AP_AXIMM_31_AWREADY(AP_AXIMM_31_AWREADY),
        .AP_AXIMM_31_WDATA(AP_AXIMM_31_WDATA),
        .AP_AXIMM_31_WSTRB(AP_AXIMM_31_WSTRB),
        .AP_AXIMM_31_WLAST(AP_AXIMM_31_WLAST),
        .AP_AXIMM_31_WVALID(AP_AXIMM_31_WVALID),
        .AP_AXIMM_31_WREADY(AP_AXIMM_31_WREADY),
        .AP_AXIMM_31_BRESP(AP_AXIMM_31_BRESP),
        .AP_AXIMM_31_BVALID(AP_AXIMM_31_BVALID),
        .AP_AXIMM_31_BREADY(AP_AXIMM_31_BREADY),
        .AP_AXIMM_31_ARADDR(AP_AXIMM_31_ARADDR),
        .AP_AXIMM_31_ARLEN(AP_AXIMM_31_ARLEN),
        .AP_AXIMM_31_ARSIZE(AP_AXIMM_31_ARSIZE),
        .AP_AXIMM_31_ARBURST(AP_AXIMM_31_ARBURST),
        .AP_AXIMM_31_ARLOCK(AP_AXIMM_31_ARLOCK),
        .AP_AXIMM_31_ARCACHE(AP_AXIMM_31_ARCACHE),
        .AP_AXIMM_31_ARPROT(AP_AXIMM_31_ARPROT),
        .AP_AXIMM_31_ARREGION(AP_AXIMM_31_ARREGION),
        .AP_AXIMM_31_ARQOS(AP_AXIMM_31_ARQOS),
        .AP_AXIMM_31_ARVALID(AP_AXIMM_31_ARVALID),
        .AP_AXIMM_31_ARREADY(AP_AXIMM_31_ARREADY),
        .AP_AXIMM_31_RDATA(AP_AXIMM_31_RDATA),
        .AP_AXIMM_31_RRESP(AP_AXIMM_31_RRESP),
        .AP_AXIMM_31_RLAST(AP_AXIMM_31_RLAST),
        .AP_AXIMM_31_RVALID(AP_AXIMM_31_RVALID),
        .AP_AXIMM_31_RREADY(AP_AXIMM_31_RREADY),
        .M_AXIMM_31_AWADDR(M_AXIMM_31_AWADDR),
        .M_AXIMM_31_AWLEN(M_AXIMM_31_AWLEN),
        .M_AXIMM_31_AWSIZE(M_AXIMM_31_AWSIZE),
        .M_AXIMM_31_AWBURST(M_AXIMM_31_AWBURST),
        .M_AXIMM_31_AWLOCK(M_AXIMM_31_AWLOCK),
        .M_AXIMM_31_AWCACHE(M_AXIMM_31_AWCACHE),
        .M_AXIMM_31_AWPROT(M_AXIMM_31_AWPROT),
        .M_AXIMM_31_AWREGION(M_AXIMM_31_AWREGION),
        .M_AXIMM_31_AWQOS(M_AXIMM_31_AWQOS),
        .M_AXIMM_31_AWVALID(M_AXIMM_31_AWVALID),
        .M_AXIMM_31_AWREADY(M_AXIMM_31_AWREADY),
        .M_AXIMM_31_WDATA(M_AXIMM_31_WDATA),
        .M_AXIMM_31_WSTRB(M_AXIMM_31_WSTRB),
        .M_AXIMM_31_WLAST(M_AXIMM_31_WLAST),
        .M_AXIMM_31_WVALID(M_AXIMM_31_WVALID),
        .M_AXIMM_31_WREADY(M_AXIMM_31_WREADY),
        .M_AXIMM_31_BRESP(M_AXIMM_31_BRESP),
        .M_AXIMM_31_BVALID(M_AXIMM_31_BVALID),
        .M_AXIMM_31_BREADY(M_AXIMM_31_BREADY),
        .M_AXIMM_31_ARADDR(M_AXIMM_31_ARADDR),
        .M_AXIMM_31_ARLEN(M_AXIMM_31_ARLEN),
        .M_AXIMM_31_ARSIZE(M_AXIMM_31_ARSIZE),
        .M_AXIMM_31_ARBURST(M_AXIMM_31_ARBURST),
        .M_AXIMM_31_ARLOCK(M_AXIMM_31_ARLOCK),
        .M_AXIMM_31_ARCACHE(M_AXIMM_31_ARCACHE),
        .M_AXIMM_31_ARPROT(M_AXIMM_31_ARPROT),
        .M_AXIMM_31_ARREGION(M_AXIMM_31_ARREGION),
        .M_AXIMM_31_ARQOS(M_AXIMM_31_ARQOS),
        .M_AXIMM_31_ARVALID(M_AXIMM_31_ARVALID),
        .M_AXIMM_31_ARREADY(M_AXIMM_31_ARREADY),
        .M_AXIMM_31_RDATA(M_AXIMM_31_RDATA),
        .M_AXIMM_31_RRESP(M_AXIMM_31_RRESP),
        .M_AXIMM_31_RLAST(M_AXIMM_31_RLAST),
        .M_AXIMM_31_RVALID(M_AXIMM_31_RVALID),
        .M_AXIMM_31_RREADY(M_AXIMM_31_RREADY),
        .AP_AXIMM_32_AWADDR(AP_AXIMM_32_AWADDR),
        .AP_AXIMM_32_AWLEN(AP_AXIMM_32_AWLEN),
        .AP_AXIMM_32_AWSIZE(AP_AXIMM_32_AWSIZE),
        .AP_AXIMM_32_AWBURST(AP_AXIMM_32_AWBURST),
        .AP_AXIMM_32_AWLOCK(AP_AXIMM_32_AWLOCK),
        .AP_AXIMM_32_AWCACHE(AP_AXIMM_32_AWCACHE),
        .AP_AXIMM_32_AWPROT(AP_AXIMM_32_AWPROT),
        .AP_AXIMM_32_AWREGION(AP_AXIMM_32_AWREGION),
        .AP_AXIMM_32_AWQOS(AP_AXIMM_32_AWQOS),
        .AP_AXIMM_32_AWVALID(AP_AXIMM_32_AWVALID),
        .AP_AXIMM_32_AWREADY(AP_AXIMM_32_AWREADY),
        .AP_AXIMM_32_WDATA(AP_AXIMM_32_WDATA),
        .AP_AXIMM_32_WSTRB(AP_AXIMM_32_WSTRB),
        .AP_AXIMM_32_WLAST(AP_AXIMM_32_WLAST),
        .AP_AXIMM_32_WVALID(AP_AXIMM_32_WVALID),
        .AP_AXIMM_32_WREADY(AP_AXIMM_32_WREADY),
        .AP_AXIMM_32_BRESP(AP_AXIMM_32_BRESP),
        .AP_AXIMM_32_BVALID(AP_AXIMM_32_BVALID),
        .AP_AXIMM_32_BREADY(AP_AXIMM_32_BREADY),
        .AP_AXIMM_32_ARADDR(AP_AXIMM_32_ARADDR),
        .AP_AXIMM_32_ARLEN(AP_AXIMM_32_ARLEN),
        .AP_AXIMM_32_ARSIZE(AP_AXIMM_32_ARSIZE),
        .AP_AXIMM_32_ARBURST(AP_AXIMM_32_ARBURST),
        .AP_AXIMM_32_ARLOCK(AP_AXIMM_32_ARLOCK),
        .AP_AXIMM_32_ARCACHE(AP_AXIMM_32_ARCACHE),
        .AP_AXIMM_32_ARPROT(AP_AXIMM_32_ARPROT),
        .AP_AXIMM_32_ARREGION(AP_AXIMM_32_ARREGION),
        .AP_AXIMM_32_ARQOS(AP_AXIMM_32_ARQOS),
        .AP_AXIMM_32_ARVALID(AP_AXIMM_32_ARVALID),
        .AP_AXIMM_32_ARREADY(AP_AXIMM_32_ARREADY),
        .AP_AXIMM_32_RDATA(AP_AXIMM_32_RDATA),
        .AP_AXIMM_32_RRESP(AP_AXIMM_32_RRESP),
        .AP_AXIMM_32_RLAST(AP_AXIMM_32_RLAST),
        .AP_AXIMM_32_RVALID(AP_AXIMM_32_RVALID),
        .AP_AXIMM_32_RREADY(AP_AXIMM_32_RREADY),
        .M_AXIMM_32_AWADDR(M_AXIMM_32_AWADDR),
        .M_AXIMM_32_AWLEN(M_AXIMM_32_AWLEN),
        .M_AXIMM_32_AWSIZE(M_AXIMM_32_AWSIZE),
        .M_AXIMM_32_AWBURST(M_AXIMM_32_AWBURST),
        .M_AXIMM_32_AWLOCK(M_AXIMM_32_AWLOCK),
        .M_AXIMM_32_AWCACHE(M_AXIMM_32_AWCACHE),
        .M_AXIMM_32_AWPROT(M_AXIMM_32_AWPROT),
        .M_AXIMM_32_AWREGION(M_AXIMM_32_AWREGION),
        .M_AXIMM_32_AWQOS(M_AXIMM_32_AWQOS),
        .M_AXIMM_32_AWVALID(M_AXIMM_32_AWVALID),
        .M_AXIMM_32_AWREADY(M_AXIMM_32_AWREADY),
        .M_AXIMM_32_WDATA(M_AXIMM_32_WDATA),
        .M_AXIMM_32_WSTRB(M_AXIMM_32_WSTRB),
        .M_AXIMM_32_WLAST(M_AXIMM_32_WLAST),
        .M_AXIMM_32_WVALID(M_AXIMM_32_WVALID),
        .M_AXIMM_32_WREADY(M_AXIMM_32_WREADY),
        .M_AXIMM_32_BRESP(M_AXIMM_32_BRESP),
        .M_AXIMM_32_BVALID(M_AXIMM_32_BVALID),
        .M_AXIMM_32_BREADY(M_AXIMM_32_BREADY),
        .M_AXIMM_32_ARADDR(M_AXIMM_32_ARADDR),
        .M_AXIMM_32_ARLEN(M_AXIMM_32_ARLEN),
        .M_AXIMM_32_ARSIZE(M_AXIMM_32_ARSIZE),
        .M_AXIMM_32_ARBURST(M_AXIMM_32_ARBURST),
        .M_AXIMM_32_ARLOCK(M_AXIMM_32_ARLOCK),
        .M_AXIMM_32_ARCACHE(M_AXIMM_32_ARCACHE),
        .M_AXIMM_32_ARPROT(M_AXIMM_32_ARPROT),
        .M_AXIMM_32_ARREGION(M_AXIMM_32_ARREGION),
        .M_AXIMM_32_ARQOS(M_AXIMM_32_ARQOS),
        .M_AXIMM_32_ARVALID(M_AXIMM_32_ARVALID),
        .M_AXIMM_32_ARREADY(M_AXIMM_32_ARREADY),
        .M_AXIMM_32_RDATA(M_AXIMM_32_RDATA),
        .M_AXIMM_32_RRESP(M_AXIMM_32_RRESP),
        .M_AXIMM_32_RLAST(M_AXIMM_32_RLAST),
        .M_AXIMM_32_RVALID(M_AXIMM_32_RVALID),
        .M_AXIMM_32_RREADY(M_AXIMM_32_RREADY),
        .AP_AXIMM_33_AWADDR(AP_AXIMM_33_AWADDR),
        .AP_AXIMM_33_AWLEN(AP_AXIMM_33_AWLEN),
        .AP_AXIMM_33_AWSIZE(AP_AXIMM_33_AWSIZE),
        .AP_AXIMM_33_AWBURST(AP_AXIMM_33_AWBURST),
        .AP_AXIMM_33_AWLOCK(AP_AXIMM_33_AWLOCK),
        .AP_AXIMM_33_AWCACHE(AP_AXIMM_33_AWCACHE),
        .AP_AXIMM_33_AWPROT(AP_AXIMM_33_AWPROT),
        .AP_AXIMM_33_AWREGION(AP_AXIMM_33_AWREGION),
        .AP_AXIMM_33_AWQOS(AP_AXIMM_33_AWQOS),
        .AP_AXIMM_33_AWVALID(AP_AXIMM_33_AWVALID),
        .AP_AXIMM_33_AWREADY(AP_AXIMM_33_AWREADY),
        .AP_AXIMM_33_WDATA(AP_AXIMM_33_WDATA),
        .AP_AXIMM_33_WSTRB(AP_AXIMM_33_WSTRB),
        .AP_AXIMM_33_WLAST(AP_AXIMM_33_WLAST),
        .AP_AXIMM_33_WVALID(AP_AXIMM_33_WVALID),
        .AP_AXIMM_33_WREADY(AP_AXIMM_33_WREADY),
        .AP_AXIMM_33_BRESP(AP_AXIMM_33_BRESP),
        .AP_AXIMM_33_BVALID(AP_AXIMM_33_BVALID),
        .AP_AXIMM_33_BREADY(AP_AXIMM_33_BREADY),
        .AP_AXIMM_33_ARADDR(AP_AXIMM_33_ARADDR),
        .AP_AXIMM_33_ARLEN(AP_AXIMM_33_ARLEN),
        .AP_AXIMM_33_ARSIZE(AP_AXIMM_33_ARSIZE),
        .AP_AXIMM_33_ARBURST(AP_AXIMM_33_ARBURST),
        .AP_AXIMM_33_ARLOCK(AP_AXIMM_33_ARLOCK),
        .AP_AXIMM_33_ARCACHE(AP_AXIMM_33_ARCACHE),
        .AP_AXIMM_33_ARPROT(AP_AXIMM_33_ARPROT),
        .AP_AXIMM_33_ARREGION(AP_AXIMM_33_ARREGION),
        .AP_AXIMM_33_ARQOS(AP_AXIMM_33_ARQOS),
        .AP_AXIMM_33_ARVALID(AP_AXIMM_33_ARVALID),
        .AP_AXIMM_33_ARREADY(AP_AXIMM_33_ARREADY),
        .AP_AXIMM_33_RDATA(AP_AXIMM_33_RDATA),
        .AP_AXIMM_33_RRESP(AP_AXIMM_33_RRESP),
        .AP_AXIMM_33_RLAST(AP_AXIMM_33_RLAST),
        .AP_AXIMM_33_RVALID(AP_AXIMM_33_RVALID),
        .AP_AXIMM_33_RREADY(AP_AXIMM_33_RREADY),
        .M_AXIMM_33_AWADDR(M_AXIMM_33_AWADDR),
        .M_AXIMM_33_AWLEN(M_AXIMM_33_AWLEN),
        .M_AXIMM_33_AWSIZE(M_AXIMM_33_AWSIZE),
        .M_AXIMM_33_AWBURST(M_AXIMM_33_AWBURST),
        .M_AXIMM_33_AWLOCK(M_AXIMM_33_AWLOCK),
        .M_AXIMM_33_AWCACHE(M_AXIMM_33_AWCACHE),
        .M_AXIMM_33_AWPROT(M_AXIMM_33_AWPROT),
        .M_AXIMM_33_AWREGION(M_AXIMM_33_AWREGION),
        .M_AXIMM_33_AWQOS(M_AXIMM_33_AWQOS),
        .M_AXIMM_33_AWVALID(M_AXIMM_33_AWVALID),
        .M_AXIMM_33_AWREADY(M_AXIMM_33_AWREADY),
        .M_AXIMM_33_WDATA(M_AXIMM_33_WDATA),
        .M_AXIMM_33_WSTRB(M_AXIMM_33_WSTRB),
        .M_AXIMM_33_WLAST(M_AXIMM_33_WLAST),
        .M_AXIMM_33_WVALID(M_AXIMM_33_WVALID),
        .M_AXIMM_33_WREADY(M_AXIMM_33_WREADY),
        .M_AXIMM_33_BRESP(M_AXIMM_33_BRESP),
        .M_AXIMM_33_BVALID(M_AXIMM_33_BVALID),
        .M_AXIMM_33_BREADY(M_AXIMM_33_BREADY),
        .M_AXIMM_33_ARADDR(M_AXIMM_33_ARADDR),
        .M_AXIMM_33_ARLEN(M_AXIMM_33_ARLEN),
        .M_AXIMM_33_ARSIZE(M_AXIMM_33_ARSIZE),
        .M_AXIMM_33_ARBURST(M_AXIMM_33_ARBURST),
        .M_AXIMM_33_ARLOCK(M_AXIMM_33_ARLOCK),
        .M_AXIMM_33_ARCACHE(M_AXIMM_33_ARCACHE),
        .M_AXIMM_33_ARPROT(M_AXIMM_33_ARPROT),
        .M_AXIMM_33_ARREGION(M_AXIMM_33_ARREGION),
        .M_AXIMM_33_ARQOS(M_AXIMM_33_ARQOS),
        .M_AXIMM_33_ARVALID(M_AXIMM_33_ARVALID),
        .M_AXIMM_33_ARREADY(M_AXIMM_33_ARREADY),
        .M_AXIMM_33_RDATA(M_AXIMM_33_RDATA),
        .M_AXIMM_33_RRESP(M_AXIMM_33_RRESP),
        .M_AXIMM_33_RLAST(M_AXIMM_33_RLAST),
        .M_AXIMM_33_RVALID(M_AXIMM_33_RVALID),
        .M_AXIMM_33_RREADY(M_AXIMM_33_RREADY),
        .AP_AXIMM_34_AWADDR(AP_AXIMM_34_AWADDR),
        .AP_AXIMM_34_AWLEN(AP_AXIMM_34_AWLEN),
        .AP_AXIMM_34_AWSIZE(AP_AXIMM_34_AWSIZE),
        .AP_AXIMM_34_AWBURST(AP_AXIMM_34_AWBURST),
        .AP_AXIMM_34_AWLOCK(AP_AXIMM_34_AWLOCK),
        .AP_AXIMM_34_AWCACHE(AP_AXIMM_34_AWCACHE),
        .AP_AXIMM_34_AWPROT(AP_AXIMM_34_AWPROT),
        .AP_AXIMM_34_AWREGION(AP_AXIMM_34_AWREGION),
        .AP_AXIMM_34_AWQOS(AP_AXIMM_34_AWQOS),
        .AP_AXIMM_34_AWVALID(AP_AXIMM_34_AWVALID),
        .AP_AXIMM_34_AWREADY(AP_AXIMM_34_AWREADY),
        .AP_AXIMM_34_WDATA(AP_AXIMM_34_WDATA),
        .AP_AXIMM_34_WSTRB(AP_AXIMM_34_WSTRB),
        .AP_AXIMM_34_WLAST(AP_AXIMM_34_WLAST),
        .AP_AXIMM_34_WVALID(AP_AXIMM_34_WVALID),
        .AP_AXIMM_34_WREADY(AP_AXIMM_34_WREADY),
        .AP_AXIMM_34_BRESP(AP_AXIMM_34_BRESP),
        .AP_AXIMM_34_BVALID(AP_AXIMM_34_BVALID),
        .AP_AXIMM_34_BREADY(AP_AXIMM_34_BREADY),
        .AP_AXIMM_34_ARADDR(AP_AXIMM_34_ARADDR),
        .AP_AXIMM_34_ARLEN(AP_AXIMM_34_ARLEN),
        .AP_AXIMM_34_ARSIZE(AP_AXIMM_34_ARSIZE),
        .AP_AXIMM_34_ARBURST(AP_AXIMM_34_ARBURST),
        .AP_AXIMM_34_ARLOCK(AP_AXIMM_34_ARLOCK),
        .AP_AXIMM_34_ARCACHE(AP_AXIMM_34_ARCACHE),
        .AP_AXIMM_34_ARPROT(AP_AXIMM_34_ARPROT),
        .AP_AXIMM_34_ARREGION(AP_AXIMM_34_ARREGION),
        .AP_AXIMM_34_ARQOS(AP_AXIMM_34_ARQOS),
        .AP_AXIMM_34_ARVALID(AP_AXIMM_34_ARVALID),
        .AP_AXIMM_34_ARREADY(AP_AXIMM_34_ARREADY),
        .AP_AXIMM_34_RDATA(AP_AXIMM_34_RDATA),
        .AP_AXIMM_34_RRESP(AP_AXIMM_34_RRESP),
        .AP_AXIMM_34_RLAST(AP_AXIMM_34_RLAST),
        .AP_AXIMM_34_RVALID(AP_AXIMM_34_RVALID),
        .AP_AXIMM_34_RREADY(AP_AXIMM_34_RREADY),
        .M_AXIMM_34_AWADDR(M_AXIMM_34_AWADDR),
        .M_AXIMM_34_AWLEN(M_AXIMM_34_AWLEN),
        .M_AXIMM_34_AWSIZE(M_AXIMM_34_AWSIZE),
        .M_AXIMM_34_AWBURST(M_AXIMM_34_AWBURST),
        .M_AXIMM_34_AWLOCK(M_AXIMM_34_AWLOCK),
        .M_AXIMM_34_AWCACHE(M_AXIMM_34_AWCACHE),
        .M_AXIMM_34_AWPROT(M_AXIMM_34_AWPROT),
        .M_AXIMM_34_AWREGION(M_AXIMM_34_AWREGION),
        .M_AXIMM_34_AWQOS(M_AXIMM_34_AWQOS),
        .M_AXIMM_34_AWVALID(M_AXIMM_34_AWVALID),
        .M_AXIMM_34_AWREADY(M_AXIMM_34_AWREADY),
        .M_AXIMM_34_WDATA(M_AXIMM_34_WDATA),
        .M_AXIMM_34_WSTRB(M_AXIMM_34_WSTRB),
        .M_AXIMM_34_WLAST(M_AXIMM_34_WLAST),
        .M_AXIMM_34_WVALID(M_AXIMM_34_WVALID),
        .M_AXIMM_34_WREADY(M_AXIMM_34_WREADY),
        .M_AXIMM_34_BRESP(M_AXIMM_34_BRESP),
        .M_AXIMM_34_BVALID(M_AXIMM_34_BVALID),
        .M_AXIMM_34_BREADY(M_AXIMM_34_BREADY),
        .M_AXIMM_34_ARADDR(M_AXIMM_34_ARADDR),
        .M_AXIMM_34_ARLEN(M_AXIMM_34_ARLEN),
        .M_AXIMM_34_ARSIZE(M_AXIMM_34_ARSIZE),
        .M_AXIMM_34_ARBURST(M_AXIMM_34_ARBURST),
        .M_AXIMM_34_ARLOCK(M_AXIMM_34_ARLOCK),
        .M_AXIMM_34_ARCACHE(M_AXIMM_34_ARCACHE),
        .M_AXIMM_34_ARPROT(M_AXIMM_34_ARPROT),
        .M_AXIMM_34_ARREGION(M_AXIMM_34_ARREGION),
        .M_AXIMM_34_ARQOS(M_AXIMM_34_ARQOS),
        .M_AXIMM_34_ARVALID(M_AXIMM_34_ARVALID),
        .M_AXIMM_34_ARREADY(M_AXIMM_34_ARREADY),
        .M_AXIMM_34_RDATA(M_AXIMM_34_RDATA),
        .M_AXIMM_34_RRESP(M_AXIMM_34_RRESP),
        .M_AXIMM_34_RLAST(M_AXIMM_34_RLAST),
        .M_AXIMM_34_RVALID(M_AXIMM_34_RVALID),
        .M_AXIMM_34_RREADY(M_AXIMM_34_RREADY),
        .AP_AXIMM_35_AWADDR(AP_AXIMM_35_AWADDR),
        .AP_AXIMM_35_AWLEN(AP_AXIMM_35_AWLEN),
        .AP_AXIMM_35_AWSIZE(AP_AXIMM_35_AWSIZE),
        .AP_AXIMM_35_AWBURST(AP_AXIMM_35_AWBURST),
        .AP_AXIMM_35_AWLOCK(AP_AXIMM_35_AWLOCK),
        .AP_AXIMM_35_AWCACHE(AP_AXIMM_35_AWCACHE),
        .AP_AXIMM_35_AWPROT(AP_AXIMM_35_AWPROT),
        .AP_AXIMM_35_AWREGION(AP_AXIMM_35_AWREGION),
        .AP_AXIMM_35_AWQOS(AP_AXIMM_35_AWQOS),
        .AP_AXIMM_35_AWVALID(AP_AXIMM_35_AWVALID),
        .AP_AXIMM_35_AWREADY(AP_AXIMM_35_AWREADY),
        .AP_AXIMM_35_WDATA(AP_AXIMM_35_WDATA),
        .AP_AXIMM_35_WSTRB(AP_AXIMM_35_WSTRB),
        .AP_AXIMM_35_WLAST(AP_AXIMM_35_WLAST),
        .AP_AXIMM_35_WVALID(AP_AXIMM_35_WVALID),
        .AP_AXIMM_35_WREADY(AP_AXIMM_35_WREADY),
        .AP_AXIMM_35_BRESP(AP_AXIMM_35_BRESP),
        .AP_AXIMM_35_BVALID(AP_AXIMM_35_BVALID),
        .AP_AXIMM_35_BREADY(AP_AXIMM_35_BREADY),
        .AP_AXIMM_35_ARADDR(AP_AXIMM_35_ARADDR),
        .AP_AXIMM_35_ARLEN(AP_AXIMM_35_ARLEN),
        .AP_AXIMM_35_ARSIZE(AP_AXIMM_35_ARSIZE),
        .AP_AXIMM_35_ARBURST(AP_AXIMM_35_ARBURST),
        .AP_AXIMM_35_ARLOCK(AP_AXIMM_35_ARLOCK),
        .AP_AXIMM_35_ARCACHE(AP_AXIMM_35_ARCACHE),
        .AP_AXIMM_35_ARPROT(AP_AXIMM_35_ARPROT),
        .AP_AXIMM_35_ARREGION(AP_AXIMM_35_ARREGION),
        .AP_AXIMM_35_ARQOS(AP_AXIMM_35_ARQOS),
        .AP_AXIMM_35_ARVALID(AP_AXIMM_35_ARVALID),
        .AP_AXIMM_35_ARREADY(AP_AXIMM_35_ARREADY),
        .AP_AXIMM_35_RDATA(AP_AXIMM_35_RDATA),
        .AP_AXIMM_35_RRESP(AP_AXIMM_35_RRESP),
        .AP_AXIMM_35_RLAST(AP_AXIMM_35_RLAST),
        .AP_AXIMM_35_RVALID(AP_AXIMM_35_RVALID),
        .AP_AXIMM_35_RREADY(AP_AXIMM_35_RREADY),
        .M_AXIMM_35_AWADDR(M_AXIMM_35_AWADDR),
        .M_AXIMM_35_AWLEN(M_AXIMM_35_AWLEN),
        .M_AXIMM_35_AWSIZE(M_AXIMM_35_AWSIZE),
        .M_AXIMM_35_AWBURST(M_AXIMM_35_AWBURST),
        .M_AXIMM_35_AWLOCK(M_AXIMM_35_AWLOCK),
        .M_AXIMM_35_AWCACHE(M_AXIMM_35_AWCACHE),
        .M_AXIMM_35_AWPROT(M_AXIMM_35_AWPROT),
        .M_AXIMM_35_AWREGION(M_AXIMM_35_AWREGION),
        .M_AXIMM_35_AWQOS(M_AXIMM_35_AWQOS),
        .M_AXIMM_35_AWVALID(M_AXIMM_35_AWVALID),
        .M_AXIMM_35_AWREADY(M_AXIMM_35_AWREADY),
        .M_AXIMM_35_WDATA(M_AXIMM_35_WDATA),
        .M_AXIMM_35_WSTRB(M_AXIMM_35_WSTRB),
        .M_AXIMM_35_WLAST(M_AXIMM_35_WLAST),
        .M_AXIMM_35_WVALID(M_AXIMM_35_WVALID),
        .M_AXIMM_35_WREADY(M_AXIMM_35_WREADY),
        .M_AXIMM_35_BRESP(M_AXIMM_35_BRESP),
        .M_AXIMM_35_BVALID(M_AXIMM_35_BVALID),
        .M_AXIMM_35_BREADY(M_AXIMM_35_BREADY),
        .M_AXIMM_35_ARADDR(M_AXIMM_35_ARADDR),
        .M_AXIMM_35_ARLEN(M_AXIMM_35_ARLEN),
        .M_AXIMM_35_ARSIZE(M_AXIMM_35_ARSIZE),
        .M_AXIMM_35_ARBURST(M_AXIMM_35_ARBURST),
        .M_AXIMM_35_ARLOCK(M_AXIMM_35_ARLOCK),
        .M_AXIMM_35_ARCACHE(M_AXIMM_35_ARCACHE),
        .M_AXIMM_35_ARPROT(M_AXIMM_35_ARPROT),
        .M_AXIMM_35_ARREGION(M_AXIMM_35_ARREGION),
        .M_AXIMM_35_ARQOS(M_AXIMM_35_ARQOS),
        .M_AXIMM_35_ARVALID(M_AXIMM_35_ARVALID),
        .M_AXIMM_35_ARREADY(M_AXIMM_35_ARREADY),
        .M_AXIMM_35_RDATA(M_AXIMM_35_RDATA),
        .M_AXIMM_35_RRESP(M_AXIMM_35_RRESP),
        .M_AXIMM_35_RLAST(M_AXIMM_35_RLAST),
        .M_AXIMM_35_RVALID(M_AXIMM_35_RVALID),
        .M_AXIMM_35_RREADY(M_AXIMM_35_RREADY),
        .AP_AXIMM_36_AWADDR(AP_AXIMM_36_AWADDR),
        .AP_AXIMM_36_AWLEN(AP_AXIMM_36_AWLEN),
        .AP_AXIMM_36_AWSIZE(AP_AXIMM_36_AWSIZE),
        .AP_AXIMM_36_AWBURST(AP_AXIMM_36_AWBURST),
        .AP_AXIMM_36_AWLOCK(AP_AXIMM_36_AWLOCK),
        .AP_AXIMM_36_AWCACHE(AP_AXIMM_36_AWCACHE),
        .AP_AXIMM_36_AWPROT(AP_AXIMM_36_AWPROT),
        .AP_AXIMM_36_AWREGION(AP_AXIMM_36_AWREGION),
        .AP_AXIMM_36_AWQOS(AP_AXIMM_36_AWQOS),
        .AP_AXIMM_36_AWVALID(AP_AXIMM_36_AWVALID),
        .AP_AXIMM_36_AWREADY(AP_AXIMM_36_AWREADY),
        .AP_AXIMM_36_WDATA(AP_AXIMM_36_WDATA),
        .AP_AXIMM_36_WSTRB(AP_AXIMM_36_WSTRB),
        .AP_AXIMM_36_WLAST(AP_AXIMM_36_WLAST),
        .AP_AXIMM_36_WVALID(AP_AXIMM_36_WVALID),
        .AP_AXIMM_36_WREADY(AP_AXIMM_36_WREADY),
        .AP_AXIMM_36_BRESP(AP_AXIMM_36_BRESP),
        .AP_AXIMM_36_BVALID(AP_AXIMM_36_BVALID),
        .AP_AXIMM_36_BREADY(AP_AXIMM_36_BREADY),
        .AP_AXIMM_36_ARADDR(AP_AXIMM_36_ARADDR),
        .AP_AXIMM_36_ARLEN(AP_AXIMM_36_ARLEN),
        .AP_AXIMM_36_ARSIZE(AP_AXIMM_36_ARSIZE),
        .AP_AXIMM_36_ARBURST(AP_AXIMM_36_ARBURST),
        .AP_AXIMM_36_ARLOCK(AP_AXIMM_36_ARLOCK),
        .AP_AXIMM_36_ARCACHE(AP_AXIMM_36_ARCACHE),
        .AP_AXIMM_36_ARPROT(AP_AXIMM_36_ARPROT),
        .AP_AXIMM_36_ARREGION(AP_AXIMM_36_ARREGION),
        .AP_AXIMM_36_ARQOS(AP_AXIMM_36_ARQOS),
        .AP_AXIMM_36_ARVALID(AP_AXIMM_36_ARVALID),
        .AP_AXIMM_36_ARREADY(AP_AXIMM_36_ARREADY),
        .AP_AXIMM_36_RDATA(AP_AXIMM_36_RDATA),
        .AP_AXIMM_36_RRESP(AP_AXIMM_36_RRESP),
        .AP_AXIMM_36_RLAST(AP_AXIMM_36_RLAST),
        .AP_AXIMM_36_RVALID(AP_AXIMM_36_RVALID),
        .AP_AXIMM_36_RREADY(AP_AXIMM_36_RREADY),
        .M_AXIMM_36_AWADDR(M_AXIMM_36_AWADDR),
        .M_AXIMM_36_AWLEN(M_AXIMM_36_AWLEN),
        .M_AXIMM_36_AWSIZE(M_AXIMM_36_AWSIZE),
        .M_AXIMM_36_AWBURST(M_AXIMM_36_AWBURST),
        .M_AXIMM_36_AWLOCK(M_AXIMM_36_AWLOCK),
        .M_AXIMM_36_AWCACHE(M_AXIMM_36_AWCACHE),
        .M_AXIMM_36_AWPROT(M_AXIMM_36_AWPROT),
        .M_AXIMM_36_AWREGION(M_AXIMM_36_AWREGION),
        .M_AXIMM_36_AWQOS(M_AXIMM_36_AWQOS),
        .M_AXIMM_36_AWVALID(M_AXIMM_36_AWVALID),
        .M_AXIMM_36_AWREADY(M_AXIMM_36_AWREADY),
        .M_AXIMM_36_WDATA(M_AXIMM_36_WDATA),
        .M_AXIMM_36_WSTRB(M_AXIMM_36_WSTRB),
        .M_AXIMM_36_WLAST(M_AXIMM_36_WLAST),
        .M_AXIMM_36_WVALID(M_AXIMM_36_WVALID),
        .M_AXIMM_36_WREADY(M_AXIMM_36_WREADY),
        .M_AXIMM_36_BRESP(M_AXIMM_36_BRESP),
        .M_AXIMM_36_BVALID(M_AXIMM_36_BVALID),
        .M_AXIMM_36_BREADY(M_AXIMM_36_BREADY),
        .M_AXIMM_36_ARADDR(M_AXIMM_36_ARADDR),
        .M_AXIMM_36_ARLEN(M_AXIMM_36_ARLEN),
        .M_AXIMM_36_ARSIZE(M_AXIMM_36_ARSIZE),
        .M_AXIMM_36_ARBURST(M_AXIMM_36_ARBURST),
        .M_AXIMM_36_ARLOCK(M_AXIMM_36_ARLOCK),
        .M_AXIMM_36_ARCACHE(M_AXIMM_36_ARCACHE),
        .M_AXIMM_36_ARPROT(M_AXIMM_36_ARPROT),
        .M_AXIMM_36_ARREGION(M_AXIMM_36_ARREGION),
        .M_AXIMM_36_ARQOS(M_AXIMM_36_ARQOS),
        .M_AXIMM_36_ARVALID(M_AXIMM_36_ARVALID),
        .M_AXIMM_36_ARREADY(M_AXIMM_36_ARREADY),
        .M_AXIMM_36_RDATA(M_AXIMM_36_RDATA),
        .M_AXIMM_36_RRESP(M_AXIMM_36_RRESP),
        .M_AXIMM_36_RLAST(M_AXIMM_36_RLAST),
        .M_AXIMM_36_RVALID(M_AXIMM_36_RVALID),
        .M_AXIMM_36_RREADY(M_AXIMM_36_RREADY),
        .AP_AXIMM_37_AWADDR(AP_AXIMM_37_AWADDR),
        .AP_AXIMM_37_AWLEN(AP_AXIMM_37_AWLEN),
        .AP_AXIMM_37_AWSIZE(AP_AXIMM_37_AWSIZE),
        .AP_AXIMM_37_AWBURST(AP_AXIMM_37_AWBURST),
        .AP_AXIMM_37_AWLOCK(AP_AXIMM_37_AWLOCK),
        .AP_AXIMM_37_AWCACHE(AP_AXIMM_37_AWCACHE),
        .AP_AXIMM_37_AWPROT(AP_AXIMM_37_AWPROT),
        .AP_AXIMM_37_AWREGION(AP_AXIMM_37_AWREGION),
        .AP_AXIMM_37_AWQOS(AP_AXIMM_37_AWQOS),
        .AP_AXIMM_37_AWVALID(AP_AXIMM_37_AWVALID),
        .AP_AXIMM_37_AWREADY(AP_AXIMM_37_AWREADY),
        .AP_AXIMM_37_WDATA(AP_AXIMM_37_WDATA),
        .AP_AXIMM_37_WSTRB(AP_AXIMM_37_WSTRB),
        .AP_AXIMM_37_WLAST(AP_AXIMM_37_WLAST),
        .AP_AXIMM_37_WVALID(AP_AXIMM_37_WVALID),
        .AP_AXIMM_37_WREADY(AP_AXIMM_37_WREADY),
        .AP_AXIMM_37_BRESP(AP_AXIMM_37_BRESP),
        .AP_AXIMM_37_BVALID(AP_AXIMM_37_BVALID),
        .AP_AXIMM_37_BREADY(AP_AXIMM_37_BREADY),
        .AP_AXIMM_37_ARADDR(AP_AXIMM_37_ARADDR),
        .AP_AXIMM_37_ARLEN(AP_AXIMM_37_ARLEN),
        .AP_AXIMM_37_ARSIZE(AP_AXIMM_37_ARSIZE),
        .AP_AXIMM_37_ARBURST(AP_AXIMM_37_ARBURST),
        .AP_AXIMM_37_ARLOCK(AP_AXIMM_37_ARLOCK),
        .AP_AXIMM_37_ARCACHE(AP_AXIMM_37_ARCACHE),
        .AP_AXIMM_37_ARPROT(AP_AXIMM_37_ARPROT),
        .AP_AXIMM_37_ARREGION(AP_AXIMM_37_ARREGION),
        .AP_AXIMM_37_ARQOS(AP_AXIMM_37_ARQOS),
        .AP_AXIMM_37_ARVALID(AP_AXIMM_37_ARVALID),
        .AP_AXIMM_37_ARREADY(AP_AXIMM_37_ARREADY),
        .AP_AXIMM_37_RDATA(AP_AXIMM_37_RDATA),
        .AP_AXIMM_37_RRESP(AP_AXIMM_37_RRESP),
        .AP_AXIMM_37_RLAST(AP_AXIMM_37_RLAST),
        .AP_AXIMM_37_RVALID(AP_AXIMM_37_RVALID),
        .AP_AXIMM_37_RREADY(AP_AXIMM_37_RREADY),
        .M_AXIMM_37_AWADDR(M_AXIMM_37_AWADDR),
        .M_AXIMM_37_AWLEN(M_AXIMM_37_AWLEN),
        .M_AXIMM_37_AWSIZE(M_AXIMM_37_AWSIZE),
        .M_AXIMM_37_AWBURST(M_AXIMM_37_AWBURST),
        .M_AXIMM_37_AWLOCK(M_AXIMM_37_AWLOCK),
        .M_AXIMM_37_AWCACHE(M_AXIMM_37_AWCACHE),
        .M_AXIMM_37_AWPROT(M_AXIMM_37_AWPROT),
        .M_AXIMM_37_AWREGION(M_AXIMM_37_AWREGION),
        .M_AXIMM_37_AWQOS(M_AXIMM_37_AWQOS),
        .M_AXIMM_37_AWVALID(M_AXIMM_37_AWVALID),
        .M_AXIMM_37_AWREADY(M_AXIMM_37_AWREADY),
        .M_AXIMM_37_WDATA(M_AXIMM_37_WDATA),
        .M_AXIMM_37_WSTRB(M_AXIMM_37_WSTRB),
        .M_AXIMM_37_WLAST(M_AXIMM_37_WLAST),
        .M_AXIMM_37_WVALID(M_AXIMM_37_WVALID),
        .M_AXIMM_37_WREADY(M_AXIMM_37_WREADY),
        .M_AXIMM_37_BRESP(M_AXIMM_37_BRESP),
        .M_AXIMM_37_BVALID(M_AXIMM_37_BVALID),
        .M_AXIMM_37_BREADY(M_AXIMM_37_BREADY),
        .M_AXIMM_37_ARADDR(M_AXIMM_37_ARADDR),
        .M_AXIMM_37_ARLEN(M_AXIMM_37_ARLEN),
        .M_AXIMM_37_ARSIZE(M_AXIMM_37_ARSIZE),
        .M_AXIMM_37_ARBURST(M_AXIMM_37_ARBURST),
        .M_AXIMM_37_ARLOCK(M_AXIMM_37_ARLOCK),
        .M_AXIMM_37_ARCACHE(M_AXIMM_37_ARCACHE),
        .M_AXIMM_37_ARPROT(M_AXIMM_37_ARPROT),
        .M_AXIMM_37_ARREGION(M_AXIMM_37_ARREGION),
        .M_AXIMM_37_ARQOS(M_AXIMM_37_ARQOS),
        .M_AXIMM_37_ARVALID(M_AXIMM_37_ARVALID),
        .M_AXIMM_37_ARREADY(M_AXIMM_37_ARREADY),
        .M_AXIMM_37_RDATA(M_AXIMM_37_RDATA),
        .M_AXIMM_37_RRESP(M_AXIMM_37_RRESP),
        .M_AXIMM_37_RLAST(M_AXIMM_37_RLAST),
        .M_AXIMM_37_RVALID(M_AXIMM_37_RVALID),
        .M_AXIMM_37_RREADY(M_AXIMM_37_RREADY),
        .AP_AXIMM_38_AWADDR(AP_AXIMM_38_AWADDR),
        .AP_AXIMM_38_AWLEN(AP_AXIMM_38_AWLEN),
        .AP_AXIMM_38_AWSIZE(AP_AXIMM_38_AWSIZE),
        .AP_AXIMM_38_AWBURST(AP_AXIMM_38_AWBURST),
        .AP_AXIMM_38_AWLOCK(AP_AXIMM_38_AWLOCK),
        .AP_AXIMM_38_AWCACHE(AP_AXIMM_38_AWCACHE),
        .AP_AXIMM_38_AWPROT(AP_AXIMM_38_AWPROT),
        .AP_AXIMM_38_AWREGION(AP_AXIMM_38_AWREGION),
        .AP_AXIMM_38_AWQOS(AP_AXIMM_38_AWQOS),
        .AP_AXIMM_38_AWVALID(AP_AXIMM_38_AWVALID),
        .AP_AXIMM_38_AWREADY(AP_AXIMM_38_AWREADY),
        .AP_AXIMM_38_WDATA(AP_AXIMM_38_WDATA),
        .AP_AXIMM_38_WSTRB(AP_AXIMM_38_WSTRB),
        .AP_AXIMM_38_WLAST(AP_AXIMM_38_WLAST),
        .AP_AXIMM_38_WVALID(AP_AXIMM_38_WVALID),
        .AP_AXIMM_38_WREADY(AP_AXIMM_38_WREADY),
        .AP_AXIMM_38_BRESP(AP_AXIMM_38_BRESP),
        .AP_AXIMM_38_BVALID(AP_AXIMM_38_BVALID),
        .AP_AXIMM_38_BREADY(AP_AXIMM_38_BREADY),
        .AP_AXIMM_38_ARADDR(AP_AXIMM_38_ARADDR),
        .AP_AXIMM_38_ARLEN(AP_AXIMM_38_ARLEN),
        .AP_AXIMM_38_ARSIZE(AP_AXIMM_38_ARSIZE),
        .AP_AXIMM_38_ARBURST(AP_AXIMM_38_ARBURST),
        .AP_AXIMM_38_ARLOCK(AP_AXIMM_38_ARLOCK),
        .AP_AXIMM_38_ARCACHE(AP_AXIMM_38_ARCACHE),
        .AP_AXIMM_38_ARPROT(AP_AXIMM_38_ARPROT),
        .AP_AXIMM_38_ARREGION(AP_AXIMM_38_ARREGION),
        .AP_AXIMM_38_ARQOS(AP_AXIMM_38_ARQOS),
        .AP_AXIMM_38_ARVALID(AP_AXIMM_38_ARVALID),
        .AP_AXIMM_38_ARREADY(AP_AXIMM_38_ARREADY),
        .AP_AXIMM_38_RDATA(AP_AXIMM_38_RDATA),
        .AP_AXIMM_38_RRESP(AP_AXIMM_38_RRESP),
        .AP_AXIMM_38_RLAST(AP_AXIMM_38_RLAST),
        .AP_AXIMM_38_RVALID(AP_AXIMM_38_RVALID),
        .AP_AXIMM_38_RREADY(AP_AXIMM_38_RREADY),
        .M_AXIMM_38_AWADDR(M_AXIMM_38_AWADDR),
        .M_AXIMM_38_AWLEN(M_AXIMM_38_AWLEN),
        .M_AXIMM_38_AWSIZE(M_AXIMM_38_AWSIZE),
        .M_AXIMM_38_AWBURST(M_AXIMM_38_AWBURST),
        .M_AXIMM_38_AWLOCK(M_AXIMM_38_AWLOCK),
        .M_AXIMM_38_AWCACHE(M_AXIMM_38_AWCACHE),
        .M_AXIMM_38_AWPROT(M_AXIMM_38_AWPROT),
        .M_AXIMM_38_AWREGION(M_AXIMM_38_AWREGION),
        .M_AXIMM_38_AWQOS(M_AXIMM_38_AWQOS),
        .M_AXIMM_38_AWVALID(M_AXIMM_38_AWVALID),
        .M_AXIMM_38_AWREADY(M_AXIMM_38_AWREADY),
        .M_AXIMM_38_WDATA(M_AXIMM_38_WDATA),
        .M_AXIMM_38_WSTRB(M_AXIMM_38_WSTRB),
        .M_AXIMM_38_WLAST(M_AXIMM_38_WLAST),
        .M_AXIMM_38_WVALID(M_AXIMM_38_WVALID),
        .M_AXIMM_38_WREADY(M_AXIMM_38_WREADY),
        .M_AXIMM_38_BRESP(M_AXIMM_38_BRESP),
        .M_AXIMM_38_BVALID(M_AXIMM_38_BVALID),
        .M_AXIMM_38_BREADY(M_AXIMM_38_BREADY),
        .M_AXIMM_38_ARADDR(M_AXIMM_38_ARADDR),
        .M_AXIMM_38_ARLEN(M_AXIMM_38_ARLEN),
        .M_AXIMM_38_ARSIZE(M_AXIMM_38_ARSIZE),
        .M_AXIMM_38_ARBURST(M_AXIMM_38_ARBURST),
        .M_AXIMM_38_ARLOCK(M_AXIMM_38_ARLOCK),
        .M_AXIMM_38_ARCACHE(M_AXIMM_38_ARCACHE),
        .M_AXIMM_38_ARPROT(M_AXIMM_38_ARPROT),
        .M_AXIMM_38_ARREGION(M_AXIMM_38_ARREGION),
        .M_AXIMM_38_ARQOS(M_AXIMM_38_ARQOS),
        .M_AXIMM_38_ARVALID(M_AXIMM_38_ARVALID),
        .M_AXIMM_38_ARREADY(M_AXIMM_38_ARREADY),
        .M_AXIMM_38_RDATA(M_AXIMM_38_RDATA),
        .M_AXIMM_38_RRESP(M_AXIMM_38_RRESP),
        .M_AXIMM_38_RLAST(M_AXIMM_38_RLAST),
        .M_AXIMM_38_RVALID(M_AXIMM_38_RVALID),
        .M_AXIMM_38_RREADY(M_AXIMM_38_RREADY),
        .AP_AXIMM_39_AWADDR(AP_AXIMM_39_AWADDR),
        .AP_AXIMM_39_AWLEN(AP_AXIMM_39_AWLEN),
        .AP_AXIMM_39_AWSIZE(AP_AXIMM_39_AWSIZE),
        .AP_AXIMM_39_AWBURST(AP_AXIMM_39_AWBURST),
        .AP_AXIMM_39_AWLOCK(AP_AXIMM_39_AWLOCK),
        .AP_AXIMM_39_AWCACHE(AP_AXIMM_39_AWCACHE),
        .AP_AXIMM_39_AWPROT(AP_AXIMM_39_AWPROT),
        .AP_AXIMM_39_AWREGION(AP_AXIMM_39_AWREGION),
        .AP_AXIMM_39_AWQOS(AP_AXIMM_39_AWQOS),
        .AP_AXIMM_39_AWVALID(AP_AXIMM_39_AWVALID),
        .AP_AXIMM_39_AWREADY(AP_AXIMM_39_AWREADY),
        .AP_AXIMM_39_WDATA(AP_AXIMM_39_WDATA),
        .AP_AXIMM_39_WSTRB(AP_AXIMM_39_WSTRB),
        .AP_AXIMM_39_WLAST(AP_AXIMM_39_WLAST),
        .AP_AXIMM_39_WVALID(AP_AXIMM_39_WVALID),
        .AP_AXIMM_39_WREADY(AP_AXIMM_39_WREADY),
        .AP_AXIMM_39_BRESP(AP_AXIMM_39_BRESP),
        .AP_AXIMM_39_BVALID(AP_AXIMM_39_BVALID),
        .AP_AXIMM_39_BREADY(AP_AXIMM_39_BREADY),
        .AP_AXIMM_39_ARADDR(AP_AXIMM_39_ARADDR),
        .AP_AXIMM_39_ARLEN(AP_AXIMM_39_ARLEN),
        .AP_AXIMM_39_ARSIZE(AP_AXIMM_39_ARSIZE),
        .AP_AXIMM_39_ARBURST(AP_AXIMM_39_ARBURST),
        .AP_AXIMM_39_ARLOCK(AP_AXIMM_39_ARLOCK),
        .AP_AXIMM_39_ARCACHE(AP_AXIMM_39_ARCACHE),
        .AP_AXIMM_39_ARPROT(AP_AXIMM_39_ARPROT),
        .AP_AXIMM_39_ARREGION(AP_AXIMM_39_ARREGION),
        .AP_AXIMM_39_ARQOS(AP_AXIMM_39_ARQOS),
        .AP_AXIMM_39_ARVALID(AP_AXIMM_39_ARVALID),
        .AP_AXIMM_39_ARREADY(AP_AXIMM_39_ARREADY),
        .AP_AXIMM_39_RDATA(AP_AXIMM_39_RDATA),
        .AP_AXIMM_39_RRESP(AP_AXIMM_39_RRESP),
        .AP_AXIMM_39_RLAST(AP_AXIMM_39_RLAST),
        .AP_AXIMM_39_RVALID(AP_AXIMM_39_RVALID),
        .AP_AXIMM_39_RREADY(AP_AXIMM_39_RREADY),
        .M_AXIMM_39_AWADDR(M_AXIMM_39_AWADDR),
        .M_AXIMM_39_AWLEN(M_AXIMM_39_AWLEN),
        .M_AXIMM_39_AWSIZE(M_AXIMM_39_AWSIZE),
        .M_AXIMM_39_AWBURST(M_AXIMM_39_AWBURST),
        .M_AXIMM_39_AWLOCK(M_AXIMM_39_AWLOCK),
        .M_AXIMM_39_AWCACHE(M_AXIMM_39_AWCACHE),
        .M_AXIMM_39_AWPROT(M_AXIMM_39_AWPROT),
        .M_AXIMM_39_AWREGION(M_AXIMM_39_AWREGION),
        .M_AXIMM_39_AWQOS(M_AXIMM_39_AWQOS),
        .M_AXIMM_39_AWVALID(M_AXIMM_39_AWVALID),
        .M_AXIMM_39_AWREADY(M_AXIMM_39_AWREADY),
        .M_AXIMM_39_WDATA(M_AXIMM_39_WDATA),
        .M_AXIMM_39_WSTRB(M_AXIMM_39_WSTRB),
        .M_AXIMM_39_WLAST(M_AXIMM_39_WLAST),
        .M_AXIMM_39_WVALID(M_AXIMM_39_WVALID),
        .M_AXIMM_39_WREADY(M_AXIMM_39_WREADY),
        .M_AXIMM_39_BRESP(M_AXIMM_39_BRESP),
        .M_AXIMM_39_BVALID(M_AXIMM_39_BVALID),
        .M_AXIMM_39_BREADY(M_AXIMM_39_BREADY),
        .M_AXIMM_39_ARADDR(M_AXIMM_39_ARADDR),
        .M_AXIMM_39_ARLEN(M_AXIMM_39_ARLEN),
        .M_AXIMM_39_ARSIZE(M_AXIMM_39_ARSIZE),
        .M_AXIMM_39_ARBURST(M_AXIMM_39_ARBURST),
        .M_AXIMM_39_ARLOCK(M_AXIMM_39_ARLOCK),
        .M_AXIMM_39_ARCACHE(M_AXIMM_39_ARCACHE),
        .M_AXIMM_39_ARPROT(M_AXIMM_39_ARPROT),
        .M_AXIMM_39_ARREGION(M_AXIMM_39_ARREGION),
        .M_AXIMM_39_ARQOS(M_AXIMM_39_ARQOS),
        .M_AXIMM_39_ARVALID(M_AXIMM_39_ARVALID),
        .M_AXIMM_39_ARREADY(M_AXIMM_39_ARREADY),
        .M_AXIMM_39_RDATA(M_AXIMM_39_RDATA),
        .M_AXIMM_39_RRESP(M_AXIMM_39_RRESP),
        .M_AXIMM_39_RLAST(M_AXIMM_39_RLAST),
        .M_AXIMM_39_RVALID(M_AXIMM_39_RVALID),
        .M_AXIMM_39_RREADY(M_AXIMM_39_RREADY),
        .AP_AXIMM_40_AWADDR(AP_AXIMM_40_AWADDR),
        .AP_AXIMM_40_AWLEN(AP_AXIMM_40_AWLEN),
        .AP_AXIMM_40_AWSIZE(AP_AXIMM_40_AWSIZE),
        .AP_AXIMM_40_AWBURST(AP_AXIMM_40_AWBURST),
        .AP_AXIMM_40_AWLOCK(AP_AXIMM_40_AWLOCK),
        .AP_AXIMM_40_AWCACHE(AP_AXIMM_40_AWCACHE),
        .AP_AXIMM_40_AWPROT(AP_AXIMM_40_AWPROT),
        .AP_AXIMM_40_AWREGION(AP_AXIMM_40_AWREGION),
        .AP_AXIMM_40_AWQOS(AP_AXIMM_40_AWQOS),
        .AP_AXIMM_40_AWVALID(AP_AXIMM_40_AWVALID),
        .AP_AXIMM_40_AWREADY(AP_AXIMM_40_AWREADY),
        .AP_AXIMM_40_WDATA(AP_AXIMM_40_WDATA),
        .AP_AXIMM_40_WSTRB(AP_AXIMM_40_WSTRB),
        .AP_AXIMM_40_WLAST(AP_AXIMM_40_WLAST),
        .AP_AXIMM_40_WVALID(AP_AXIMM_40_WVALID),
        .AP_AXIMM_40_WREADY(AP_AXIMM_40_WREADY),
        .AP_AXIMM_40_BRESP(AP_AXIMM_40_BRESP),
        .AP_AXIMM_40_BVALID(AP_AXIMM_40_BVALID),
        .AP_AXIMM_40_BREADY(AP_AXIMM_40_BREADY),
        .AP_AXIMM_40_ARADDR(AP_AXIMM_40_ARADDR),
        .AP_AXIMM_40_ARLEN(AP_AXIMM_40_ARLEN),
        .AP_AXIMM_40_ARSIZE(AP_AXIMM_40_ARSIZE),
        .AP_AXIMM_40_ARBURST(AP_AXIMM_40_ARBURST),
        .AP_AXIMM_40_ARLOCK(AP_AXIMM_40_ARLOCK),
        .AP_AXIMM_40_ARCACHE(AP_AXIMM_40_ARCACHE),
        .AP_AXIMM_40_ARPROT(AP_AXIMM_40_ARPROT),
        .AP_AXIMM_40_ARREGION(AP_AXIMM_40_ARREGION),
        .AP_AXIMM_40_ARQOS(AP_AXIMM_40_ARQOS),
        .AP_AXIMM_40_ARVALID(AP_AXIMM_40_ARVALID),
        .AP_AXIMM_40_ARREADY(AP_AXIMM_40_ARREADY),
        .AP_AXIMM_40_RDATA(AP_AXIMM_40_RDATA),
        .AP_AXIMM_40_RRESP(AP_AXIMM_40_RRESP),
        .AP_AXIMM_40_RLAST(AP_AXIMM_40_RLAST),
        .AP_AXIMM_40_RVALID(AP_AXIMM_40_RVALID),
        .AP_AXIMM_40_RREADY(AP_AXIMM_40_RREADY),
        .M_AXIMM_40_AWADDR(M_AXIMM_40_AWADDR),
        .M_AXIMM_40_AWLEN(M_AXIMM_40_AWLEN),
        .M_AXIMM_40_AWSIZE(M_AXIMM_40_AWSIZE),
        .M_AXIMM_40_AWBURST(M_AXIMM_40_AWBURST),
        .M_AXIMM_40_AWLOCK(M_AXIMM_40_AWLOCK),
        .M_AXIMM_40_AWCACHE(M_AXIMM_40_AWCACHE),
        .M_AXIMM_40_AWPROT(M_AXIMM_40_AWPROT),
        .M_AXIMM_40_AWREGION(M_AXIMM_40_AWREGION),
        .M_AXIMM_40_AWQOS(M_AXIMM_40_AWQOS),
        .M_AXIMM_40_AWVALID(M_AXIMM_40_AWVALID),
        .M_AXIMM_40_AWREADY(M_AXIMM_40_AWREADY),
        .M_AXIMM_40_WDATA(M_AXIMM_40_WDATA),
        .M_AXIMM_40_WSTRB(M_AXIMM_40_WSTRB),
        .M_AXIMM_40_WLAST(M_AXIMM_40_WLAST),
        .M_AXIMM_40_WVALID(M_AXIMM_40_WVALID),
        .M_AXIMM_40_WREADY(M_AXIMM_40_WREADY),
        .M_AXIMM_40_BRESP(M_AXIMM_40_BRESP),
        .M_AXIMM_40_BVALID(M_AXIMM_40_BVALID),
        .M_AXIMM_40_BREADY(M_AXIMM_40_BREADY),
        .M_AXIMM_40_ARADDR(M_AXIMM_40_ARADDR),
        .M_AXIMM_40_ARLEN(M_AXIMM_40_ARLEN),
        .M_AXIMM_40_ARSIZE(M_AXIMM_40_ARSIZE),
        .M_AXIMM_40_ARBURST(M_AXIMM_40_ARBURST),
        .M_AXIMM_40_ARLOCK(M_AXIMM_40_ARLOCK),
        .M_AXIMM_40_ARCACHE(M_AXIMM_40_ARCACHE),
        .M_AXIMM_40_ARPROT(M_AXIMM_40_ARPROT),
        .M_AXIMM_40_ARREGION(M_AXIMM_40_ARREGION),
        .M_AXIMM_40_ARQOS(M_AXIMM_40_ARQOS),
        .M_AXIMM_40_ARVALID(M_AXIMM_40_ARVALID),
        .M_AXIMM_40_ARREADY(M_AXIMM_40_ARREADY),
        .M_AXIMM_40_RDATA(M_AXIMM_40_RDATA),
        .M_AXIMM_40_RRESP(M_AXIMM_40_RRESP),
        .M_AXIMM_40_RLAST(M_AXIMM_40_RLAST),
        .M_AXIMM_40_RVALID(M_AXIMM_40_RVALID),
        .M_AXIMM_40_RREADY(M_AXIMM_40_RREADY),
        .AP_AXIMM_41_AWADDR(AP_AXIMM_41_AWADDR),
        .AP_AXIMM_41_AWLEN(AP_AXIMM_41_AWLEN),
        .AP_AXIMM_41_AWSIZE(AP_AXIMM_41_AWSIZE),
        .AP_AXIMM_41_AWBURST(AP_AXIMM_41_AWBURST),
        .AP_AXIMM_41_AWLOCK(AP_AXIMM_41_AWLOCK),
        .AP_AXIMM_41_AWCACHE(AP_AXIMM_41_AWCACHE),
        .AP_AXIMM_41_AWPROT(AP_AXIMM_41_AWPROT),
        .AP_AXIMM_41_AWREGION(AP_AXIMM_41_AWREGION),
        .AP_AXIMM_41_AWQOS(AP_AXIMM_41_AWQOS),
        .AP_AXIMM_41_AWVALID(AP_AXIMM_41_AWVALID),
        .AP_AXIMM_41_AWREADY(AP_AXIMM_41_AWREADY),
        .AP_AXIMM_41_WDATA(AP_AXIMM_41_WDATA),
        .AP_AXIMM_41_WSTRB(AP_AXIMM_41_WSTRB),
        .AP_AXIMM_41_WLAST(AP_AXIMM_41_WLAST),
        .AP_AXIMM_41_WVALID(AP_AXIMM_41_WVALID),
        .AP_AXIMM_41_WREADY(AP_AXIMM_41_WREADY),
        .AP_AXIMM_41_BRESP(AP_AXIMM_41_BRESP),
        .AP_AXIMM_41_BVALID(AP_AXIMM_41_BVALID),
        .AP_AXIMM_41_BREADY(AP_AXIMM_41_BREADY),
        .AP_AXIMM_41_ARADDR(AP_AXIMM_41_ARADDR),
        .AP_AXIMM_41_ARLEN(AP_AXIMM_41_ARLEN),
        .AP_AXIMM_41_ARSIZE(AP_AXIMM_41_ARSIZE),
        .AP_AXIMM_41_ARBURST(AP_AXIMM_41_ARBURST),
        .AP_AXIMM_41_ARLOCK(AP_AXIMM_41_ARLOCK),
        .AP_AXIMM_41_ARCACHE(AP_AXIMM_41_ARCACHE),
        .AP_AXIMM_41_ARPROT(AP_AXIMM_41_ARPROT),
        .AP_AXIMM_41_ARREGION(AP_AXIMM_41_ARREGION),
        .AP_AXIMM_41_ARQOS(AP_AXIMM_41_ARQOS),
        .AP_AXIMM_41_ARVALID(AP_AXIMM_41_ARVALID),
        .AP_AXIMM_41_ARREADY(AP_AXIMM_41_ARREADY),
        .AP_AXIMM_41_RDATA(AP_AXIMM_41_RDATA),
        .AP_AXIMM_41_RRESP(AP_AXIMM_41_RRESP),
        .AP_AXIMM_41_RLAST(AP_AXIMM_41_RLAST),
        .AP_AXIMM_41_RVALID(AP_AXIMM_41_RVALID),
        .AP_AXIMM_41_RREADY(AP_AXIMM_41_RREADY),
        .M_AXIMM_41_AWADDR(M_AXIMM_41_AWADDR),
        .M_AXIMM_41_AWLEN(M_AXIMM_41_AWLEN),
        .M_AXIMM_41_AWSIZE(M_AXIMM_41_AWSIZE),
        .M_AXIMM_41_AWBURST(M_AXIMM_41_AWBURST),
        .M_AXIMM_41_AWLOCK(M_AXIMM_41_AWLOCK),
        .M_AXIMM_41_AWCACHE(M_AXIMM_41_AWCACHE),
        .M_AXIMM_41_AWPROT(M_AXIMM_41_AWPROT),
        .M_AXIMM_41_AWREGION(M_AXIMM_41_AWREGION),
        .M_AXIMM_41_AWQOS(M_AXIMM_41_AWQOS),
        .M_AXIMM_41_AWVALID(M_AXIMM_41_AWVALID),
        .M_AXIMM_41_AWREADY(M_AXIMM_41_AWREADY),
        .M_AXIMM_41_WDATA(M_AXIMM_41_WDATA),
        .M_AXIMM_41_WSTRB(M_AXIMM_41_WSTRB),
        .M_AXIMM_41_WLAST(M_AXIMM_41_WLAST),
        .M_AXIMM_41_WVALID(M_AXIMM_41_WVALID),
        .M_AXIMM_41_WREADY(M_AXIMM_41_WREADY),
        .M_AXIMM_41_BRESP(M_AXIMM_41_BRESP),
        .M_AXIMM_41_BVALID(M_AXIMM_41_BVALID),
        .M_AXIMM_41_BREADY(M_AXIMM_41_BREADY),
        .M_AXIMM_41_ARADDR(M_AXIMM_41_ARADDR),
        .M_AXIMM_41_ARLEN(M_AXIMM_41_ARLEN),
        .M_AXIMM_41_ARSIZE(M_AXIMM_41_ARSIZE),
        .M_AXIMM_41_ARBURST(M_AXIMM_41_ARBURST),
        .M_AXIMM_41_ARLOCK(M_AXIMM_41_ARLOCK),
        .M_AXIMM_41_ARCACHE(M_AXIMM_41_ARCACHE),
        .M_AXIMM_41_ARPROT(M_AXIMM_41_ARPROT),
        .M_AXIMM_41_ARREGION(M_AXIMM_41_ARREGION),
        .M_AXIMM_41_ARQOS(M_AXIMM_41_ARQOS),
        .M_AXIMM_41_ARVALID(M_AXIMM_41_ARVALID),
        .M_AXIMM_41_ARREADY(M_AXIMM_41_ARREADY),
        .M_AXIMM_41_RDATA(M_AXIMM_41_RDATA),
        .M_AXIMM_41_RRESP(M_AXIMM_41_RRESP),
        .M_AXIMM_41_RLAST(M_AXIMM_41_RLAST),
        .M_AXIMM_41_RVALID(M_AXIMM_41_RVALID),
        .M_AXIMM_41_RREADY(M_AXIMM_41_RREADY),
        .AP_AXIMM_42_AWADDR(AP_AXIMM_42_AWADDR),
        .AP_AXIMM_42_AWLEN(AP_AXIMM_42_AWLEN),
        .AP_AXIMM_42_AWSIZE(AP_AXIMM_42_AWSIZE),
        .AP_AXIMM_42_AWBURST(AP_AXIMM_42_AWBURST),
        .AP_AXIMM_42_AWLOCK(AP_AXIMM_42_AWLOCK),
        .AP_AXIMM_42_AWCACHE(AP_AXIMM_42_AWCACHE),
        .AP_AXIMM_42_AWPROT(AP_AXIMM_42_AWPROT),
        .AP_AXIMM_42_AWREGION(AP_AXIMM_42_AWREGION),
        .AP_AXIMM_42_AWQOS(AP_AXIMM_42_AWQOS),
        .AP_AXIMM_42_AWVALID(AP_AXIMM_42_AWVALID),
        .AP_AXIMM_42_AWREADY(AP_AXIMM_42_AWREADY),
        .AP_AXIMM_42_WDATA(AP_AXIMM_42_WDATA),
        .AP_AXIMM_42_WSTRB(AP_AXIMM_42_WSTRB),
        .AP_AXIMM_42_WLAST(AP_AXIMM_42_WLAST),
        .AP_AXIMM_42_WVALID(AP_AXIMM_42_WVALID),
        .AP_AXIMM_42_WREADY(AP_AXIMM_42_WREADY),
        .AP_AXIMM_42_BRESP(AP_AXIMM_42_BRESP),
        .AP_AXIMM_42_BVALID(AP_AXIMM_42_BVALID),
        .AP_AXIMM_42_BREADY(AP_AXIMM_42_BREADY),
        .AP_AXIMM_42_ARADDR(AP_AXIMM_42_ARADDR),
        .AP_AXIMM_42_ARLEN(AP_AXIMM_42_ARLEN),
        .AP_AXIMM_42_ARSIZE(AP_AXIMM_42_ARSIZE),
        .AP_AXIMM_42_ARBURST(AP_AXIMM_42_ARBURST),
        .AP_AXIMM_42_ARLOCK(AP_AXIMM_42_ARLOCK),
        .AP_AXIMM_42_ARCACHE(AP_AXIMM_42_ARCACHE),
        .AP_AXIMM_42_ARPROT(AP_AXIMM_42_ARPROT),
        .AP_AXIMM_42_ARREGION(AP_AXIMM_42_ARREGION),
        .AP_AXIMM_42_ARQOS(AP_AXIMM_42_ARQOS),
        .AP_AXIMM_42_ARVALID(AP_AXIMM_42_ARVALID),
        .AP_AXIMM_42_ARREADY(AP_AXIMM_42_ARREADY),
        .AP_AXIMM_42_RDATA(AP_AXIMM_42_RDATA),
        .AP_AXIMM_42_RRESP(AP_AXIMM_42_RRESP),
        .AP_AXIMM_42_RLAST(AP_AXIMM_42_RLAST),
        .AP_AXIMM_42_RVALID(AP_AXIMM_42_RVALID),
        .AP_AXIMM_42_RREADY(AP_AXIMM_42_RREADY),
        .M_AXIMM_42_AWADDR(M_AXIMM_42_AWADDR),
        .M_AXIMM_42_AWLEN(M_AXIMM_42_AWLEN),
        .M_AXIMM_42_AWSIZE(M_AXIMM_42_AWSIZE),
        .M_AXIMM_42_AWBURST(M_AXIMM_42_AWBURST),
        .M_AXIMM_42_AWLOCK(M_AXIMM_42_AWLOCK),
        .M_AXIMM_42_AWCACHE(M_AXIMM_42_AWCACHE),
        .M_AXIMM_42_AWPROT(M_AXIMM_42_AWPROT),
        .M_AXIMM_42_AWREGION(M_AXIMM_42_AWREGION),
        .M_AXIMM_42_AWQOS(M_AXIMM_42_AWQOS),
        .M_AXIMM_42_AWVALID(M_AXIMM_42_AWVALID),
        .M_AXIMM_42_AWREADY(M_AXIMM_42_AWREADY),
        .M_AXIMM_42_WDATA(M_AXIMM_42_WDATA),
        .M_AXIMM_42_WSTRB(M_AXIMM_42_WSTRB),
        .M_AXIMM_42_WLAST(M_AXIMM_42_WLAST),
        .M_AXIMM_42_WVALID(M_AXIMM_42_WVALID),
        .M_AXIMM_42_WREADY(M_AXIMM_42_WREADY),
        .M_AXIMM_42_BRESP(M_AXIMM_42_BRESP),
        .M_AXIMM_42_BVALID(M_AXIMM_42_BVALID),
        .M_AXIMM_42_BREADY(M_AXIMM_42_BREADY),
        .M_AXIMM_42_ARADDR(M_AXIMM_42_ARADDR),
        .M_AXIMM_42_ARLEN(M_AXIMM_42_ARLEN),
        .M_AXIMM_42_ARSIZE(M_AXIMM_42_ARSIZE),
        .M_AXIMM_42_ARBURST(M_AXIMM_42_ARBURST),
        .M_AXIMM_42_ARLOCK(M_AXIMM_42_ARLOCK),
        .M_AXIMM_42_ARCACHE(M_AXIMM_42_ARCACHE),
        .M_AXIMM_42_ARPROT(M_AXIMM_42_ARPROT),
        .M_AXIMM_42_ARREGION(M_AXIMM_42_ARREGION),
        .M_AXIMM_42_ARQOS(M_AXIMM_42_ARQOS),
        .M_AXIMM_42_ARVALID(M_AXIMM_42_ARVALID),
        .M_AXIMM_42_ARREADY(M_AXIMM_42_ARREADY),
        .M_AXIMM_42_RDATA(M_AXIMM_42_RDATA),
        .M_AXIMM_42_RRESP(M_AXIMM_42_RRESP),
        .M_AXIMM_42_RLAST(M_AXIMM_42_RLAST),
        .M_AXIMM_42_RVALID(M_AXIMM_42_RVALID),
        .M_AXIMM_42_RREADY(M_AXIMM_42_RREADY),
        .AP_AXIMM_43_AWADDR(AP_AXIMM_43_AWADDR),
        .AP_AXIMM_43_AWLEN(AP_AXIMM_43_AWLEN),
        .AP_AXIMM_43_AWSIZE(AP_AXIMM_43_AWSIZE),
        .AP_AXIMM_43_AWBURST(AP_AXIMM_43_AWBURST),
        .AP_AXIMM_43_AWLOCK(AP_AXIMM_43_AWLOCK),
        .AP_AXIMM_43_AWCACHE(AP_AXIMM_43_AWCACHE),
        .AP_AXIMM_43_AWPROT(AP_AXIMM_43_AWPROT),
        .AP_AXIMM_43_AWREGION(AP_AXIMM_43_AWREGION),
        .AP_AXIMM_43_AWQOS(AP_AXIMM_43_AWQOS),
        .AP_AXIMM_43_AWVALID(AP_AXIMM_43_AWVALID),
        .AP_AXIMM_43_AWREADY(AP_AXIMM_43_AWREADY),
        .AP_AXIMM_43_WDATA(AP_AXIMM_43_WDATA),
        .AP_AXIMM_43_WSTRB(AP_AXIMM_43_WSTRB),
        .AP_AXIMM_43_WLAST(AP_AXIMM_43_WLAST),
        .AP_AXIMM_43_WVALID(AP_AXIMM_43_WVALID),
        .AP_AXIMM_43_WREADY(AP_AXIMM_43_WREADY),
        .AP_AXIMM_43_BRESP(AP_AXIMM_43_BRESP),
        .AP_AXIMM_43_BVALID(AP_AXIMM_43_BVALID),
        .AP_AXIMM_43_BREADY(AP_AXIMM_43_BREADY),
        .AP_AXIMM_43_ARADDR(AP_AXIMM_43_ARADDR),
        .AP_AXIMM_43_ARLEN(AP_AXIMM_43_ARLEN),
        .AP_AXIMM_43_ARSIZE(AP_AXIMM_43_ARSIZE),
        .AP_AXIMM_43_ARBURST(AP_AXIMM_43_ARBURST),
        .AP_AXIMM_43_ARLOCK(AP_AXIMM_43_ARLOCK),
        .AP_AXIMM_43_ARCACHE(AP_AXIMM_43_ARCACHE),
        .AP_AXIMM_43_ARPROT(AP_AXIMM_43_ARPROT),
        .AP_AXIMM_43_ARREGION(AP_AXIMM_43_ARREGION),
        .AP_AXIMM_43_ARQOS(AP_AXIMM_43_ARQOS),
        .AP_AXIMM_43_ARVALID(AP_AXIMM_43_ARVALID),
        .AP_AXIMM_43_ARREADY(AP_AXIMM_43_ARREADY),
        .AP_AXIMM_43_RDATA(AP_AXIMM_43_RDATA),
        .AP_AXIMM_43_RRESP(AP_AXIMM_43_RRESP),
        .AP_AXIMM_43_RLAST(AP_AXIMM_43_RLAST),
        .AP_AXIMM_43_RVALID(AP_AXIMM_43_RVALID),
        .AP_AXIMM_43_RREADY(AP_AXIMM_43_RREADY),
        .M_AXIMM_43_AWADDR(M_AXIMM_43_AWADDR),
        .M_AXIMM_43_AWLEN(M_AXIMM_43_AWLEN),
        .M_AXIMM_43_AWSIZE(M_AXIMM_43_AWSIZE),
        .M_AXIMM_43_AWBURST(M_AXIMM_43_AWBURST),
        .M_AXIMM_43_AWLOCK(M_AXIMM_43_AWLOCK),
        .M_AXIMM_43_AWCACHE(M_AXIMM_43_AWCACHE),
        .M_AXIMM_43_AWPROT(M_AXIMM_43_AWPROT),
        .M_AXIMM_43_AWREGION(M_AXIMM_43_AWREGION),
        .M_AXIMM_43_AWQOS(M_AXIMM_43_AWQOS),
        .M_AXIMM_43_AWVALID(M_AXIMM_43_AWVALID),
        .M_AXIMM_43_AWREADY(M_AXIMM_43_AWREADY),
        .M_AXIMM_43_WDATA(M_AXIMM_43_WDATA),
        .M_AXIMM_43_WSTRB(M_AXIMM_43_WSTRB),
        .M_AXIMM_43_WLAST(M_AXIMM_43_WLAST),
        .M_AXIMM_43_WVALID(M_AXIMM_43_WVALID),
        .M_AXIMM_43_WREADY(M_AXIMM_43_WREADY),
        .M_AXIMM_43_BRESP(M_AXIMM_43_BRESP),
        .M_AXIMM_43_BVALID(M_AXIMM_43_BVALID),
        .M_AXIMM_43_BREADY(M_AXIMM_43_BREADY),
        .M_AXIMM_43_ARADDR(M_AXIMM_43_ARADDR),
        .M_AXIMM_43_ARLEN(M_AXIMM_43_ARLEN),
        .M_AXIMM_43_ARSIZE(M_AXIMM_43_ARSIZE),
        .M_AXIMM_43_ARBURST(M_AXIMM_43_ARBURST),
        .M_AXIMM_43_ARLOCK(M_AXIMM_43_ARLOCK),
        .M_AXIMM_43_ARCACHE(M_AXIMM_43_ARCACHE),
        .M_AXIMM_43_ARPROT(M_AXIMM_43_ARPROT),
        .M_AXIMM_43_ARREGION(M_AXIMM_43_ARREGION),
        .M_AXIMM_43_ARQOS(M_AXIMM_43_ARQOS),
        .M_AXIMM_43_ARVALID(M_AXIMM_43_ARVALID),
        .M_AXIMM_43_ARREADY(M_AXIMM_43_ARREADY),
        .M_AXIMM_43_RDATA(M_AXIMM_43_RDATA),
        .M_AXIMM_43_RRESP(M_AXIMM_43_RRESP),
        .M_AXIMM_43_RLAST(M_AXIMM_43_RLAST),
        .M_AXIMM_43_RVALID(M_AXIMM_43_RVALID),
        .M_AXIMM_43_RREADY(M_AXIMM_43_RREADY),
        .AP_AXIMM_44_AWADDR(AP_AXIMM_44_AWADDR),
        .AP_AXIMM_44_AWLEN(AP_AXIMM_44_AWLEN),
        .AP_AXIMM_44_AWSIZE(AP_AXIMM_44_AWSIZE),
        .AP_AXIMM_44_AWBURST(AP_AXIMM_44_AWBURST),
        .AP_AXIMM_44_AWLOCK(AP_AXIMM_44_AWLOCK),
        .AP_AXIMM_44_AWCACHE(AP_AXIMM_44_AWCACHE),
        .AP_AXIMM_44_AWPROT(AP_AXIMM_44_AWPROT),
        .AP_AXIMM_44_AWREGION(AP_AXIMM_44_AWREGION),
        .AP_AXIMM_44_AWQOS(AP_AXIMM_44_AWQOS),
        .AP_AXIMM_44_AWVALID(AP_AXIMM_44_AWVALID),
        .AP_AXIMM_44_AWREADY(AP_AXIMM_44_AWREADY),
        .AP_AXIMM_44_WDATA(AP_AXIMM_44_WDATA),
        .AP_AXIMM_44_WSTRB(AP_AXIMM_44_WSTRB),
        .AP_AXIMM_44_WLAST(AP_AXIMM_44_WLAST),
        .AP_AXIMM_44_WVALID(AP_AXIMM_44_WVALID),
        .AP_AXIMM_44_WREADY(AP_AXIMM_44_WREADY),
        .AP_AXIMM_44_BRESP(AP_AXIMM_44_BRESP),
        .AP_AXIMM_44_BVALID(AP_AXIMM_44_BVALID),
        .AP_AXIMM_44_BREADY(AP_AXIMM_44_BREADY),
        .AP_AXIMM_44_ARADDR(AP_AXIMM_44_ARADDR),
        .AP_AXIMM_44_ARLEN(AP_AXIMM_44_ARLEN),
        .AP_AXIMM_44_ARSIZE(AP_AXIMM_44_ARSIZE),
        .AP_AXIMM_44_ARBURST(AP_AXIMM_44_ARBURST),
        .AP_AXIMM_44_ARLOCK(AP_AXIMM_44_ARLOCK),
        .AP_AXIMM_44_ARCACHE(AP_AXIMM_44_ARCACHE),
        .AP_AXIMM_44_ARPROT(AP_AXIMM_44_ARPROT),
        .AP_AXIMM_44_ARREGION(AP_AXIMM_44_ARREGION),
        .AP_AXIMM_44_ARQOS(AP_AXIMM_44_ARQOS),
        .AP_AXIMM_44_ARVALID(AP_AXIMM_44_ARVALID),
        .AP_AXIMM_44_ARREADY(AP_AXIMM_44_ARREADY),
        .AP_AXIMM_44_RDATA(AP_AXIMM_44_RDATA),
        .AP_AXIMM_44_RRESP(AP_AXIMM_44_RRESP),
        .AP_AXIMM_44_RLAST(AP_AXIMM_44_RLAST),
        .AP_AXIMM_44_RVALID(AP_AXIMM_44_RVALID),
        .AP_AXIMM_44_RREADY(AP_AXIMM_44_RREADY),
        .M_AXIMM_44_AWADDR(M_AXIMM_44_AWADDR),
        .M_AXIMM_44_AWLEN(M_AXIMM_44_AWLEN),
        .M_AXIMM_44_AWSIZE(M_AXIMM_44_AWSIZE),
        .M_AXIMM_44_AWBURST(M_AXIMM_44_AWBURST),
        .M_AXIMM_44_AWLOCK(M_AXIMM_44_AWLOCK),
        .M_AXIMM_44_AWCACHE(M_AXIMM_44_AWCACHE),
        .M_AXIMM_44_AWPROT(M_AXIMM_44_AWPROT),
        .M_AXIMM_44_AWREGION(M_AXIMM_44_AWREGION),
        .M_AXIMM_44_AWQOS(M_AXIMM_44_AWQOS),
        .M_AXIMM_44_AWVALID(M_AXIMM_44_AWVALID),
        .M_AXIMM_44_AWREADY(M_AXIMM_44_AWREADY),
        .M_AXIMM_44_WDATA(M_AXIMM_44_WDATA),
        .M_AXIMM_44_WSTRB(M_AXIMM_44_WSTRB),
        .M_AXIMM_44_WLAST(M_AXIMM_44_WLAST),
        .M_AXIMM_44_WVALID(M_AXIMM_44_WVALID),
        .M_AXIMM_44_WREADY(M_AXIMM_44_WREADY),
        .M_AXIMM_44_BRESP(M_AXIMM_44_BRESP),
        .M_AXIMM_44_BVALID(M_AXIMM_44_BVALID),
        .M_AXIMM_44_BREADY(M_AXIMM_44_BREADY),
        .M_AXIMM_44_ARADDR(M_AXIMM_44_ARADDR),
        .M_AXIMM_44_ARLEN(M_AXIMM_44_ARLEN),
        .M_AXIMM_44_ARSIZE(M_AXIMM_44_ARSIZE),
        .M_AXIMM_44_ARBURST(M_AXIMM_44_ARBURST),
        .M_AXIMM_44_ARLOCK(M_AXIMM_44_ARLOCK),
        .M_AXIMM_44_ARCACHE(M_AXIMM_44_ARCACHE),
        .M_AXIMM_44_ARPROT(M_AXIMM_44_ARPROT),
        .M_AXIMM_44_ARREGION(M_AXIMM_44_ARREGION),
        .M_AXIMM_44_ARQOS(M_AXIMM_44_ARQOS),
        .M_AXIMM_44_ARVALID(M_AXIMM_44_ARVALID),
        .M_AXIMM_44_ARREADY(M_AXIMM_44_ARREADY),
        .M_AXIMM_44_RDATA(M_AXIMM_44_RDATA),
        .M_AXIMM_44_RRESP(M_AXIMM_44_RRESP),
        .M_AXIMM_44_RLAST(M_AXIMM_44_RLAST),
        .M_AXIMM_44_RVALID(M_AXIMM_44_RVALID),
        .M_AXIMM_44_RREADY(M_AXIMM_44_RREADY),
        .AP_AXIMM_45_AWADDR(AP_AXIMM_45_AWADDR),
        .AP_AXIMM_45_AWLEN(AP_AXIMM_45_AWLEN),
        .AP_AXIMM_45_AWSIZE(AP_AXIMM_45_AWSIZE),
        .AP_AXIMM_45_AWBURST(AP_AXIMM_45_AWBURST),
        .AP_AXIMM_45_AWLOCK(AP_AXIMM_45_AWLOCK),
        .AP_AXIMM_45_AWCACHE(AP_AXIMM_45_AWCACHE),
        .AP_AXIMM_45_AWPROT(AP_AXIMM_45_AWPROT),
        .AP_AXIMM_45_AWREGION(AP_AXIMM_45_AWREGION),
        .AP_AXIMM_45_AWQOS(AP_AXIMM_45_AWQOS),
        .AP_AXIMM_45_AWVALID(AP_AXIMM_45_AWVALID),
        .AP_AXIMM_45_AWREADY(AP_AXIMM_45_AWREADY),
        .AP_AXIMM_45_WDATA(AP_AXIMM_45_WDATA),
        .AP_AXIMM_45_WSTRB(AP_AXIMM_45_WSTRB),
        .AP_AXIMM_45_WLAST(AP_AXIMM_45_WLAST),
        .AP_AXIMM_45_WVALID(AP_AXIMM_45_WVALID),
        .AP_AXIMM_45_WREADY(AP_AXIMM_45_WREADY),
        .AP_AXIMM_45_BRESP(AP_AXIMM_45_BRESP),
        .AP_AXIMM_45_BVALID(AP_AXIMM_45_BVALID),
        .AP_AXIMM_45_BREADY(AP_AXIMM_45_BREADY),
        .AP_AXIMM_45_ARADDR(AP_AXIMM_45_ARADDR),
        .AP_AXIMM_45_ARLEN(AP_AXIMM_45_ARLEN),
        .AP_AXIMM_45_ARSIZE(AP_AXIMM_45_ARSIZE),
        .AP_AXIMM_45_ARBURST(AP_AXIMM_45_ARBURST),
        .AP_AXIMM_45_ARLOCK(AP_AXIMM_45_ARLOCK),
        .AP_AXIMM_45_ARCACHE(AP_AXIMM_45_ARCACHE),
        .AP_AXIMM_45_ARPROT(AP_AXIMM_45_ARPROT),
        .AP_AXIMM_45_ARREGION(AP_AXIMM_45_ARREGION),
        .AP_AXIMM_45_ARQOS(AP_AXIMM_45_ARQOS),
        .AP_AXIMM_45_ARVALID(AP_AXIMM_45_ARVALID),
        .AP_AXIMM_45_ARREADY(AP_AXIMM_45_ARREADY),
        .AP_AXIMM_45_RDATA(AP_AXIMM_45_RDATA),
        .AP_AXIMM_45_RRESP(AP_AXIMM_45_RRESP),
        .AP_AXIMM_45_RLAST(AP_AXIMM_45_RLAST),
        .AP_AXIMM_45_RVALID(AP_AXIMM_45_RVALID),
        .AP_AXIMM_45_RREADY(AP_AXIMM_45_RREADY),
        .M_AXIMM_45_AWADDR(M_AXIMM_45_AWADDR),
        .M_AXIMM_45_AWLEN(M_AXIMM_45_AWLEN),
        .M_AXIMM_45_AWSIZE(M_AXIMM_45_AWSIZE),
        .M_AXIMM_45_AWBURST(M_AXIMM_45_AWBURST),
        .M_AXIMM_45_AWLOCK(M_AXIMM_45_AWLOCK),
        .M_AXIMM_45_AWCACHE(M_AXIMM_45_AWCACHE),
        .M_AXIMM_45_AWPROT(M_AXIMM_45_AWPROT),
        .M_AXIMM_45_AWREGION(M_AXIMM_45_AWREGION),
        .M_AXIMM_45_AWQOS(M_AXIMM_45_AWQOS),
        .M_AXIMM_45_AWVALID(M_AXIMM_45_AWVALID),
        .M_AXIMM_45_AWREADY(M_AXIMM_45_AWREADY),
        .M_AXIMM_45_WDATA(M_AXIMM_45_WDATA),
        .M_AXIMM_45_WSTRB(M_AXIMM_45_WSTRB),
        .M_AXIMM_45_WLAST(M_AXIMM_45_WLAST),
        .M_AXIMM_45_WVALID(M_AXIMM_45_WVALID),
        .M_AXIMM_45_WREADY(M_AXIMM_45_WREADY),
        .M_AXIMM_45_BRESP(M_AXIMM_45_BRESP),
        .M_AXIMM_45_BVALID(M_AXIMM_45_BVALID),
        .M_AXIMM_45_BREADY(M_AXIMM_45_BREADY),
        .M_AXIMM_45_ARADDR(M_AXIMM_45_ARADDR),
        .M_AXIMM_45_ARLEN(M_AXIMM_45_ARLEN),
        .M_AXIMM_45_ARSIZE(M_AXIMM_45_ARSIZE),
        .M_AXIMM_45_ARBURST(M_AXIMM_45_ARBURST),
        .M_AXIMM_45_ARLOCK(M_AXIMM_45_ARLOCK),
        .M_AXIMM_45_ARCACHE(M_AXIMM_45_ARCACHE),
        .M_AXIMM_45_ARPROT(M_AXIMM_45_ARPROT),
        .M_AXIMM_45_ARREGION(M_AXIMM_45_ARREGION),
        .M_AXIMM_45_ARQOS(M_AXIMM_45_ARQOS),
        .M_AXIMM_45_ARVALID(M_AXIMM_45_ARVALID),
        .M_AXIMM_45_ARREADY(M_AXIMM_45_ARREADY),
        .M_AXIMM_45_RDATA(M_AXIMM_45_RDATA),
        .M_AXIMM_45_RRESP(M_AXIMM_45_RRESP),
        .M_AXIMM_45_RLAST(M_AXIMM_45_RLAST),
        .M_AXIMM_45_RVALID(M_AXIMM_45_RVALID),
        .M_AXIMM_45_RREADY(M_AXIMM_45_RREADY),
        .AP_AXIMM_46_AWADDR(AP_AXIMM_46_AWADDR),
        .AP_AXIMM_46_AWLEN(AP_AXIMM_46_AWLEN),
        .AP_AXIMM_46_AWSIZE(AP_AXIMM_46_AWSIZE),
        .AP_AXIMM_46_AWBURST(AP_AXIMM_46_AWBURST),
        .AP_AXIMM_46_AWLOCK(AP_AXIMM_46_AWLOCK),
        .AP_AXIMM_46_AWCACHE(AP_AXIMM_46_AWCACHE),
        .AP_AXIMM_46_AWPROT(AP_AXIMM_46_AWPROT),
        .AP_AXIMM_46_AWREGION(AP_AXIMM_46_AWREGION),
        .AP_AXIMM_46_AWQOS(AP_AXIMM_46_AWQOS),
        .AP_AXIMM_46_AWVALID(AP_AXIMM_46_AWVALID),
        .AP_AXIMM_46_AWREADY(AP_AXIMM_46_AWREADY),
        .AP_AXIMM_46_WDATA(AP_AXIMM_46_WDATA),
        .AP_AXIMM_46_WSTRB(AP_AXIMM_46_WSTRB),
        .AP_AXIMM_46_WLAST(AP_AXIMM_46_WLAST),
        .AP_AXIMM_46_WVALID(AP_AXIMM_46_WVALID),
        .AP_AXIMM_46_WREADY(AP_AXIMM_46_WREADY),
        .AP_AXIMM_46_BRESP(AP_AXIMM_46_BRESP),
        .AP_AXIMM_46_BVALID(AP_AXIMM_46_BVALID),
        .AP_AXIMM_46_BREADY(AP_AXIMM_46_BREADY),
        .AP_AXIMM_46_ARADDR(AP_AXIMM_46_ARADDR),
        .AP_AXIMM_46_ARLEN(AP_AXIMM_46_ARLEN),
        .AP_AXIMM_46_ARSIZE(AP_AXIMM_46_ARSIZE),
        .AP_AXIMM_46_ARBURST(AP_AXIMM_46_ARBURST),
        .AP_AXIMM_46_ARLOCK(AP_AXIMM_46_ARLOCK),
        .AP_AXIMM_46_ARCACHE(AP_AXIMM_46_ARCACHE),
        .AP_AXIMM_46_ARPROT(AP_AXIMM_46_ARPROT),
        .AP_AXIMM_46_ARREGION(AP_AXIMM_46_ARREGION),
        .AP_AXIMM_46_ARQOS(AP_AXIMM_46_ARQOS),
        .AP_AXIMM_46_ARVALID(AP_AXIMM_46_ARVALID),
        .AP_AXIMM_46_ARREADY(AP_AXIMM_46_ARREADY),
        .AP_AXIMM_46_RDATA(AP_AXIMM_46_RDATA),
        .AP_AXIMM_46_RRESP(AP_AXIMM_46_RRESP),
        .AP_AXIMM_46_RLAST(AP_AXIMM_46_RLAST),
        .AP_AXIMM_46_RVALID(AP_AXIMM_46_RVALID),
        .AP_AXIMM_46_RREADY(AP_AXIMM_46_RREADY),
        .M_AXIMM_46_AWADDR(M_AXIMM_46_AWADDR),
        .M_AXIMM_46_AWLEN(M_AXIMM_46_AWLEN),
        .M_AXIMM_46_AWSIZE(M_AXIMM_46_AWSIZE),
        .M_AXIMM_46_AWBURST(M_AXIMM_46_AWBURST),
        .M_AXIMM_46_AWLOCK(M_AXIMM_46_AWLOCK),
        .M_AXIMM_46_AWCACHE(M_AXIMM_46_AWCACHE),
        .M_AXIMM_46_AWPROT(M_AXIMM_46_AWPROT),
        .M_AXIMM_46_AWREGION(M_AXIMM_46_AWREGION),
        .M_AXIMM_46_AWQOS(M_AXIMM_46_AWQOS),
        .M_AXIMM_46_AWVALID(M_AXIMM_46_AWVALID),
        .M_AXIMM_46_AWREADY(M_AXIMM_46_AWREADY),
        .M_AXIMM_46_WDATA(M_AXIMM_46_WDATA),
        .M_AXIMM_46_WSTRB(M_AXIMM_46_WSTRB),
        .M_AXIMM_46_WLAST(M_AXIMM_46_WLAST),
        .M_AXIMM_46_WVALID(M_AXIMM_46_WVALID),
        .M_AXIMM_46_WREADY(M_AXIMM_46_WREADY),
        .M_AXIMM_46_BRESP(M_AXIMM_46_BRESP),
        .M_AXIMM_46_BVALID(M_AXIMM_46_BVALID),
        .M_AXIMM_46_BREADY(M_AXIMM_46_BREADY),
        .M_AXIMM_46_ARADDR(M_AXIMM_46_ARADDR),
        .M_AXIMM_46_ARLEN(M_AXIMM_46_ARLEN),
        .M_AXIMM_46_ARSIZE(M_AXIMM_46_ARSIZE),
        .M_AXIMM_46_ARBURST(M_AXIMM_46_ARBURST),
        .M_AXIMM_46_ARLOCK(M_AXIMM_46_ARLOCK),
        .M_AXIMM_46_ARCACHE(M_AXIMM_46_ARCACHE),
        .M_AXIMM_46_ARPROT(M_AXIMM_46_ARPROT),
        .M_AXIMM_46_ARREGION(M_AXIMM_46_ARREGION),
        .M_AXIMM_46_ARQOS(M_AXIMM_46_ARQOS),
        .M_AXIMM_46_ARVALID(M_AXIMM_46_ARVALID),
        .M_AXIMM_46_ARREADY(M_AXIMM_46_ARREADY),
        .M_AXIMM_46_RDATA(M_AXIMM_46_RDATA),
        .M_AXIMM_46_RRESP(M_AXIMM_46_RRESP),
        .M_AXIMM_46_RLAST(M_AXIMM_46_RLAST),
        .M_AXIMM_46_RVALID(M_AXIMM_46_RVALID),
        .M_AXIMM_46_RREADY(M_AXIMM_46_RREADY),
        .AP_AXIMM_47_AWADDR(AP_AXIMM_47_AWADDR),
        .AP_AXIMM_47_AWLEN(AP_AXIMM_47_AWLEN),
        .AP_AXIMM_47_AWSIZE(AP_AXIMM_47_AWSIZE),
        .AP_AXIMM_47_AWBURST(AP_AXIMM_47_AWBURST),
        .AP_AXIMM_47_AWLOCK(AP_AXIMM_47_AWLOCK),
        .AP_AXIMM_47_AWCACHE(AP_AXIMM_47_AWCACHE),
        .AP_AXIMM_47_AWPROT(AP_AXIMM_47_AWPROT),
        .AP_AXIMM_47_AWREGION(AP_AXIMM_47_AWREGION),
        .AP_AXIMM_47_AWQOS(AP_AXIMM_47_AWQOS),
        .AP_AXIMM_47_AWVALID(AP_AXIMM_47_AWVALID),
        .AP_AXIMM_47_AWREADY(AP_AXIMM_47_AWREADY),
        .AP_AXIMM_47_WDATA(AP_AXIMM_47_WDATA),
        .AP_AXIMM_47_WSTRB(AP_AXIMM_47_WSTRB),
        .AP_AXIMM_47_WLAST(AP_AXIMM_47_WLAST),
        .AP_AXIMM_47_WVALID(AP_AXIMM_47_WVALID),
        .AP_AXIMM_47_WREADY(AP_AXIMM_47_WREADY),
        .AP_AXIMM_47_BRESP(AP_AXIMM_47_BRESP),
        .AP_AXIMM_47_BVALID(AP_AXIMM_47_BVALID),
        .AP_AXIMM_47_BREADY(AP_AXIMM_47_BREADY),
        .AP_AXIMM_47_ARADDR(AP_AXIMM_47_ARADDR),
        .AP_AXIMM_47_ARLEN(AP_AXIMM_47_ARLEN),
        .AP_AXIMM_47_ARSIZE(AP_AXIMM_47_ARSIZE),
        .AP_AXIMM_47_ARBURST(AP_AXIMM_47_ARBURST),
        .AP_AXIMM_47_ARLOCK(AP_AXIMM_47_ARLOCK),
        .AP_AXIMM_47_ARCACHE(AP_AXIMM_47_ARCACHE),
        .AP_AXIMM_47_ARPROT(AP_AXIMM_47_ARPROT),
        .AP_AXIMM_47_ARREGION(AP_AXIMM_47_ARREGION),
        .AP_AXIMM_47_ARQOS(AP_AXIMM_47_ARQOS),
        .AP_AXIMM_47_ARVALID(AP_AXIMM_47_ARVALID),
        .AP_AXIMM_47_ARREADY(AP_AXIMM_47_ARREADY),
        .AP_AXIMM_47_RDATA(AP_AXIMM_47_RDATA),
        .AP_AXIMM_47_RRESP(AP_AXIMM_47_RRESP),
        .AP_AXIMM_47_RLAST(AP_AXIMM_47_RLAST),
        .AP_AXIMM_47_RVALID(AP_AXIMM_47_RVALID),
        .AP_AXIMM_47_RREADY(AP_AXIMM_47_RREADY),
        .M_AXIMM_47_AWADDR(M_AXIMM_47_AWADDR),
        .M_AXIMM_47_AWLEN(M_AXIMM_47_AWLEN),
        .M_AXIMM_47_AWSIZE(M_AXIMM_47_AWSIZE),
        .M_AXIMM_47_AWBURST(M_AXIMM_47_AWBURST),
        .M_AXIMM_47_AWLOCK(M_AXIMM_47_AWLOCK),
        .M_AXIMM_47_AWCACHE(M_AXIMM_47_AWCACHE),
        .M_AXIMM_47_AWPROT(M_AXIMM_47_AWPROT),
        .M_AXIMM_47_AWREGION(M_AXIMM_47_AWREGION),
        .M_AXIMM_47_AWQOS(M_AXIMM_47_AWQOS),
        .M_AXIMM_47_AWVALID(M_AXIMM_47_AWVALID),
        .M_AXIMM_47_AWREADY(M_AXIMM_47_AWREADY),
        .M_AXIMM_47_WDATA(M_AXIMM_47_WDATA),
        .M_AXIMM_47_WSTRB(M_AXIMM_47_WSTRB),
        .M_AXIMM_47_WLAST(M_AXIMM_47_WLAST),
        .M_AXIMM_47_WVALID(M_AXIMM_47_WVALID),
        .M_AXIMM_47_WREADY(M_AXIMM_47_WREADY),
        .M_AXIMM_47_BRESP(M_AXIMM_47_BRESP),
        .M_AXIMM_47_BVALID(M_AXIMM_47_BVALID),
        .M_AXIMM_47_BREADY(M_AXIMM_47_BREADY),
        .M_AXIMM_47_ARADDR(M_AXIMM_47_ARADDR),
        .M_AXIMM_47_ARLEN(M_AXIMM_47_ARLEN),
        .M_AXIMM_47_ARSIZE(M_AXIMM_47_ARSIZE),
        .M_AXIMM_47_ARBURST(M_AXIMM_47_ARBURST),
        .M_AXIMM_47_ARLOCK(M_AXIMM_47_ARLOCK),
        .M_AXIMM_47_ARCACHE(M_AXIMM_47_ARCACHE),
        .M_AXIMM_47_ARPROT(M_AXIMM_47_ARPROT),
        .M_AXIMM_47_ARREGION(M_AXIMM_47_ARREGION),
        .M_AXIMM_47_ARQOS(M_AXIMM_47_ARQOS),
        .M_AXIMM_47_ARVALID(M_AXIMM_47_ARVALID),
        .M_AXIMM_47_ARREADY(M_AXIMM_47_ARREADY),
        .M_AXIMM_47_RDATA(M_AXIMM_47_RDATA),
        .M_AXIMM_47_RRESP(M_AXIMM_47_RRESP),
        .M_AXIMM_47_RLAST(M_AXIMM_47_RLAST),
        .M_AXIMM_47_RVALID(M_AXIMM_47_RVALID),
        .M_AXIMM_47_RREADY(M_AXIMM_47_RREADY),
        .AP_AXIMM_48_AWADDR(AP_AXIMM_48_AWADDR),
        .AP_AXIMM_48_AWLEN(AP_AXIMM_48_AWLEN),
        .AP_AXIMM_48_AWSIZE(AP_AXIMM_48_AWSIZE),
        .AP_AXIMM_48_AWBURST(AP_AXIMM_48_AWBURST),
        .AP_AXIMM_48_AWLOCK(AP_AXIMM_48_AWLOCK),
        .AP_AXIMM_48_AWCACHE(AP_AXIMM_48_AWCACHE),
        .AP_AXIMM_48_AWPROT(AP_AXIMM_48_AWPROT),
        .AP_AXIMM_48_AWREGION(AP_AXIMM_48_AWREGION),
        .AP_AXIMM_48_AWQOS(AP_AXIMM_48_AWQOS),
        .AP_AXIMM_48_AWVALID(AP_AXIMM_48_AWVALID),
        .AP_AXIMM_48_AWREADY(AP_AXIMM_48_AWREADY),
        .AP_AXIMM_48_WDATA(AP_AXIMM_48_WDATA),
        .AP_AXIMM_48_WSTRB(AP_AXIMM_48_WSTRB),
        .AP_AXIMM_48_WLAST(AP_AXIMM_48_WLAST),
        .AP_AXIMM_48_WVALID(AP_AXIMM_48_WVALID),
        .AP_AXIMM_48_WREADY(AP_AXIMM_48_WREADY),
        .AP_AXIMM_48_BRESP(AP_AXIMM_48_BRESP),
        .AP_AXIMM_48_BVALID(AP_AXIMM_48_BVALID),
        .AP_AXIMM_48_BREADY(AP_AXIMM_48_BREADY),
        .AP_AXIMM_48_ARADDR(AP_AXIMM_48_ARADDR),
        .AP_AXIMM_48_ARLEN(AP_AXIMM_48_ARLEN),
        .AP_AXIMM_48_ARSIZE(AP_AXIMM_48_ARSIZE),
        .AP_AXIMM_48_ARBURST(AP_AXIMM_48_ARBURST),
        .AP_AXIMM_48_ARLOCK(AP_AXIMM_48_ARLOCK),
        .AP_AXIMM_48_ARCACHE(AP_AXIMM_48_ARCACHE),
        .AP_AXIMM_48_ARPROT(AP_AXIMM_48_ARPROT),
        .AP_AXIMM_48_ARREGION(AP_AXIMM_48_ARREGION),
        .AP_AXIMM_48_ARQOS(AP_AXIMM_48_ARQOS),
        .AP_AXIMM_48_ARVALID(AP_AXIMM_48_ARVALID),
        .AP_AXIMM_48_ARREADY(AP_AXIMM_48_ARREADY),
        .AP_AXIMM_48_RDATA(AP_AXIMM_48_RDATA),
        .AP_AXIMM_48_RRESP(AP_AXIMM_48_RRESP),
        .AP_AXIMM_48_RLAST(AP_AXIMM_48_RLAST),
        .AP_AXIMM_48_RVALID(AP_AXIMM_48_RVALID),
        .AP_AXIMM_48_RREADY(AP_AXIMM_48_RREADY),
        .M_AXIMM_48_AWADDR(M_AXIMM_48_AWADDR),
        .M_AXIMM_48_AWLEN(M_AXIMM_48_AWLEN),
        .M_AXIMM_48_AWSIZE(M_AXIMM_48_AWSIZE),
        .M_AXIMM_48_AWBURST(M_AXIMM_48_AWBURST),
        .M_AXIMM_48_AWLOCK(M_AXIMM_48_AWLOCK),
        .M_AXIMM_48_AWCACHE(M_AXIMM_48_AWCACHE),
        .M_AXIMM_48_AWPROT(M_AXIMM_48_AWPROT),
        .M_AXIMM_48_AWREGION(M_AXIMM_48_AWREGION),
        .M_AXIMM_48_AWQOS(M_AXIMM_48_AWQOS),
        .M_AXIMM_48_AWVALID(M_AXIMM_48_AWVALID),
        .M_AXIMM_48_AWREADY(M_AXIMM_48_AWREADY),
        .M_AXIMM_48_WDATA(M_AXIMM_48_WDATA),
        .M_AXIMM_48_WSTRB(M_AXIMM_48_WSTRB),
        .M_AXIMM_48_WLAST(M_AXIMM_48_WLAST),
        .M_AXIMM_48_WVALID(M_AXIMM_48_WVALID),
        .M_AXIMM_48_WREADY(M_AXIMM_48_WREADY),
        .M_AXIMM_48_BRESP(M_AXIMM_48_BRESP),
        .M_AXIMM_48_BVALID(M_AXIMM_48_BVALID),
        .M_AXIMM_48_BREADY(M_AXIMM_48_BREADY),
        .M_AXIMM_48_ARADDR(M_AXIMM_48_ARADDR),
        .M_AXIMM_48_ARLEN(M_AXIMM_48_ARLEN),
        .M_AXIMM_48_ARSIZE(M_AXIMM_48_ARSIZE),
        .M_AXIMM_48_ARBURST(M_AXIMM_48_ARBURST),
        .M_AXIMM_48_ARLOCK(M_AXIMM_48_ARLOCK),
        .M_AXIMM_48_ARCACHE(M_AXIMM_48_ARCACHE),
        .M_AXIMM_48_ARPROT(M_AXIMM_48_ARPROT),
        .M_AXIMM_48_ARREGION(M_AXIMM_48_ARREGION),
        .M_AXIMM_48_ARQOS(M_AXIMM_48_ARQOS),
        .M_AXIMM_48_ARVALID(M_AXIMM_48_ARVALID),
        .M_AXIMM_48_ARREADY(M_AXIMM_48_ARREADY),
        .M_AXIMM_48_RDATA(M_AXIMM_48_RDATA),
        .M_AXIMM_48_RRESP(M_AXIMM_48_RRESP),
        .M_AXIMM_48_RLAST(M_AXIMM_48_RLAST),
        .M_AXIMM_48_RVALID(M_AXIMM_48_RVALID),
        .M_AXIMM_48_RREADY(M_AXIMM_48_RREADY),
        .AP_AXIMM_49_AWADDR(AP_AXIMM_49_AWADDR),
        .AP_AXIMM_49_AWLEN(AP_AXIMM_49_AWLEN),
        .AP_AXIMM_49_AWSIZE(AP_AXIMM_49_AWSIZE),
        .AP_AXIMM_49_AWBURST(AP_AXIMM_49_AWBURST),
        .AP_AXIMM_49_AWLOCK(AP_AXIMM_49_AWLOCK),
        .AP_AXIMM_49_AWCACHE(AP_AXIMM_49_AWCACHE),
        .AP_AXIMM_49_AWPROT(AP_AXIMM_49_AWPROT),
        .AP_AXIMM_49_AWREGION(AP_AXIMM_49_AWREGION),
        .AP_AXIMM_49_AWQOS(AP_AXIMM_49_AWQOS),
        .AP_AXIMM_49_AWVALID(AP_AXIMM_49_AWVALID),
        .AP_AXIMM_49_AWREADY(AP_AXIMM_49_AWREADY),
        .AP_AXIMM_49_WDATA(AP_AXIMM_49_WDATA),
        .AP_AXIMM_49_WSTRB(AP_AXIMM_49_WSTRB),
        .AP_AXIMM_49_WLAST(AP_AXIMM_49_WLAST),
        .AP_AXIMM_49_WVALID(AP_AXIMM_49_WVALID),
        .AP_AXIMM_49_WREADY(AP_AXIMM_49_WREADY),
        .AP_AXIMM_49_BRESP(AP_AXIMM_49_BRESP),
        .AP_AXIMM_49_BVALID(AP_AXIMM_49_BVALID),
        .AP_AXIMM_49_BREADY(AP_AXIMM_49_BREADY),
        .AP_AXIMM_49_ARADDR(AP_AXIMM_49_ARADDR),
        .AP_AXIMM_49_ARLEN(AP_AXIMM_49_ARLEN),
        .AP_AXIMM_49_ARSIZE(AP_AXIMM_49_ARSIZE),
        .AP_AXIMM_49_ARBURST(AP_AXIMM_49_ARBURST),
        .AP_AXIMM_49_ARLOCK(AP_AXIMM_49_ARLOCK),
        .AP_AXIMM_49_ARCACHE(AP_AXIMM_49_ARCACHE),
        .AP_AXIMM_49_ARPROT(AP_AXIMM_49_ARPROT),
        .AP_AXIMM_49_ARREGION(AP_AXIMM_49_ARREGION),
        .AP_AXIMM_49_ARQOS(AP_AXIMM_49_ARQOS),
        .AP_AXIMM_49_ARVALID(AP_AXIMM_49_ARVALID),
        .AP_AXIMM_49_ARREADY(AP_AXIMM_49_ARREADY),
        .AP_AXIMM_49_RDATA(AP_AXIMM_49_RDATA),
        .AP_AXIMM_49_RRESP(AP_AXIMM_49_RRESP),
        .AP_AXIMM_49_RLAST(AP_AXIMM_49_RLAST),
        .AP_AXIMM_49_RVALID(AP_AXIMM_49_RVALID),
        .AP_AXIMM_49_RREADY(AP_AXIMM_49_RREADY),
        .M_AXIMM_49_AWADDR(M_AXIMM_49_AWADDR),
        .M_AXIMM_49_AWLEN(M_AXIMM_49_AWLEN),
        .M_AXIMM_49_AWSIZE(M_AXIMM_49_AWSIZE),
        .M_AXIMM_49_AWBURST(M_AXIMM_49_AWBURST),
        .M_AXIMM_49_AWLOCK(M_AXIMM_49_AWLOCK),
        .M_AXIMM_49_AWCACHE(M_AXIMM_49_AWCACHE),
        .M_AXIMM_49_AWPROT(M_AXIMM_49_AWPROT),
        .M_AXIMM_49_AWREGION(M_AXIMM_49_AWREGION),
        .M_AXIMM_49_AWQOS(M_AXIMM_49_AWQOS),
        .M_AXIMM_49_AWVALID(M_AXIMM_49_AWVALID),
        .M_AXIMM_49_AWREADY(M_AXIMM_49_AWREADY),
        .M_AXIMM_49_WDATA(M_AXIMM_49_WDATA),
        .M_AXIMM_49_WSTRB(M_AXIMM_49_WSTRB),
        .M_AXIMM_49_WLAST(M_AXIMM_49_WLAST),
        .M_AXIMM_49_WVALID(M_AXIMM_49_WVALID),
        .M_AXIMM_49_WREADY(M_AXIMM_49_WREADY),
        .M_AXIMM_49_BRESP(M_AXIMM_49_BRESP),
        .M_AXIMM_49_BVALID(M_AXIMM_49_BVALID),
        .M_AXIMM_49_BREADY(M_AXIMM_49_BREADY),
        .M_AXIMM_49_ARADDR(M_AXIMM_49_ARADDR),
        .M_AXIMM_49_ARLEN(M_AXIMM_49_ARLEN),
        .M_AXIMM_49_ARSIZE(M_AXIMM_49_ARSIZE),
        .M_AXIMM_49_ARBURST(M_AXIMM_49_ARBURST),
        .M_AXIMM_49_ARLOCK(M_AXIMM_49_ARLOCK),
        .M_AXIMM_49_ARCACHE(M_AXIMM_49_ARCACHE),
        .M_AXIMM_49_ARPROT(M_AXIMM_49_ARPROT),
        .M_AXIMM_49_ARREGION(M_AXIMM_49_ARREGION),
        .M_AXIMM_49_ARQOS(M_AXIMM_49_ARQOS),
        .M_AXIMM_49_ARVALID(M_AXIMM_49_ARVALID),
        .M_AXIMM_49_ARREADY(M_AXIMM_49_ARREADY),
        .M_AXIMM_49_RDATA(M_AXIMM_49_RDATA),
        .M_AXIMM_49_RRESP(M_AXIMM_49_RRESP),
        .M_AXIMM_49_RLAST(M_AXIMM_49_RLAST),
        .M_AXIMM_49_RVALID(M_AXIMM_49_RVALID),
        .M_AXIMM_49_RREADY(M_AXIMM_49_RREADY),
        .AP_AXIMM_50_AWADDR(AP_AXIMM_50_AWADDR),
        .AP_AXIMM_50_AWLEN(AP_AXIMM_50_AWLEN),
        .AP_AXIMM_50_AWSIZE(AP_AXIMM_50_AWSIZE),
        .AP_AXIMM_50_AWBURST(AP_AXIMM_50_AWBURST),
        .AP_AXIMM_50_AWLOCK(AP_AXIMM_50_AWLOCK),
        .AP_AXIMM_50_AWCACHE(AP_AXIMM_50_AWCACHE),
        .AP_AXIMM_50_AWPROT(AP_AXIMM_50_AWPROT),
        .AP_AXIMM_50_AWREGION(AP_AXIMM_50_AWREGION),
        .AP_AXIMM_50_AWQOS(AP_AXIMM_50_AWQOS),
        .AP_AXIMM_50_AWVALID(AP_AXIMM_50_AWVALID),
        .AP_AXIMM_50_AWREADY(AP_AXIMM_50_AWREADY),
        .AP_AXIMM_50_WDATA(AP_AXIMM_50_WDATA),
        .AP_AXIMM_50_WSTRB(AP_AXIMM_50_WSTRB),
        .AP_AXIMM_50_WLAST(AP_AXIMM_50_WLAST),
        .AP_AXIMM_50_WVALID(AP_AXIMM_50_WVALID),
        .AP_AXIMM_50_WREADY(AP_AXIMM_50_WREADY),
        .AP_AXIMM_50_BRESP(AP_AXIMM_50_BRESP),
        .AP_AXIMM_50_BVALID(AP_AXIMM_50_BVALID),
        .AP_AXIMM_50_BREADY(AP_AXIMM_50_BREADY),
        .AP_AXIMM_50_ARADDR(AP_AXIMM_50_ARADDR),
        .AP_AXIMM_50_ARLEN(AP_AXIMM_50_ARLEN),
        .AP_AXIMM_50_ARSIZE(AP_AXIMM_50_ARSIZE),
        .AP_AXIMM_50_ARBURST(AP_AXIMM_50_ARBURST),
        .AP_AXIMM_50_ARLOCK(AP_AXIMM_50_ARLOCK),
        .AP_AXIMM_50_ARCACHE(AP_AXIMM_50_ARCACHE),
        .AP_AXIMM_50_ARPROT(AP_AXIMM_50_ARPROT),
        .AP_AXIMM_50_ARREGION(AP_AXIMM_50_ARREGION),
        .AP_AXIMM_50_ARQOS(AP_AXIMM_50_ARQOS),
        .AP_AXIMM_50_ARVALID(AP_AXIMM_50_ARVALID),
        .AP_AXIMM_50_ARREADY(AP_AXIMM_50_ARREADY),
        .AP_AXIMM_50_RDATA(AP_AXIMM_50_RDATA),
        .AP_AXIMM_50_RRESP(AP_AXIMM_50_RRESP),
        .AP_AXIMM_50_RLAST(AP_AXIMM_50_RLAST),
        .AP_AXIMM_50_RVALID(AP_AXIMM_50_RVALID),
        .AP_AXIMM_50_RREADY(AP_AXIMM_50_RREADY),
        .M_AXIMM_50_AWADDR(M_AXIMM_50_AWADDR),
        .M_AXIMM_50_AWLEN(M_AXIMM_50_AWLEN),
        .M_AXIMM_50_AWSIZE(M_AXIMM_50_AWSIZE),
        .M_AXIMM_50_AWBURST(M_AXIMM_50_AWBURST),
        .M_AXIMM_50_AWLOCK(M_AXIMM_50_AWLOCK),
        .M_AXIMM_50_AWCACHE(M_AXIMM_50_AWCACHE),
        .M_AXIMM_50_AWPROT(M_AXIMM_50_AWPROT),
        .M_AXIMM_50_AWREGION(M_AXIMM_50_AWREGION),
        .M_AXIMM_50_AWQOS(M_AXIMM_50_AWQOS),
        .M_AXIMM_50_AWVALID(M_AXIMM_50_AWVALID),
        .M_AXIMM_50_AWREADY(M_AXIMM_50_AWREADY),
        .M_AXIMM_50_WDATA(M_AXIMM_50_WDATA),
        .M_AXIMM_50_WSTRB(M_AXIMM_50_WSTRB),
        .M_AXIMM_50_WLAST(M_AXIMM_50_WLAST),
        .M_AXIMM_50_WVALID(M_AXIMM_50_WVALID),
        .M_AXIMM_50_WREADY(M_AXIMM_50_WREADY),
        .M_AXIMM_50_BRESP(M_AXIMM_50_BRESP),
        .M_AXIMM_50_BVALID(M_AXIMM_50_BVALID),
        .M_AXIMM_50_BREADY(M_AXIMM_50_BREADY),
        .M_AXIMM_50_ARADDR(M_AXIMM_50_ARADDR),
        .M_AXIMM_50_ARLEN(M_AXIMM_50_ARLEN),
        .M_AXIMM_50_ARSIZE(M_AXIMM_50_ARSIZE),
        .M_AXIMM_50_ARBURST(M_AXIMM_50_ARBURST),
        .M_AXIMM_50_ARLOCK(M_AXIMM_50_ARLOCK),
        .M_AXIMM_50_ARCACHE(M_AXIMM_50_ARCACHE),
        .M_AXIMM_50_ARPROT(M_AXIMM_50_ARPROT),
        .M_AXIMM_50_ARREGION(M_AXIMM_50_ARREGION),
        .M_AXIMM_50_ARQOS(M_AXIMM_50_ARQOS),
        .M_AXIMM_50_ARVALID(M_AXIMM_50_ARVALID),
        .M_AXIMM_50_ARREADY(M_AXIMM_50_ARREADY),
        .M_AXIMM_50_RDATA(M_AXIMM_50_RDATA),
        .M_AXIMM_50_RRESP(M_AXIMM_50_RRESP),
        .M_AXIMM_50_RLAST(M_AXIMM_50_RLAST),
        .M_AXIMM_50_RVALID(M_AXIMM_50_RVALID),
        .M_AXIMM_50_RREADY(M_AXIMM_50_RREADY),
        .AP_AXIMM_51_AWADDR(AP_AXIMM_51_AWADDR),
        .AP_AXIMM_51_AWLEN(AP_AXIMM_51_AWLEN),
        .AP_AXIMM_51_AWSIZE(AP_AXIMM_51_AWSIZE),
        .AP_AXIMM_51_AWBURST(AP_AXIMM_51_AWBURST),
        .AP_AXIMM_51_AWLOCK(AP_AXIMM_51_AWLOCK),
        .AP_AXIMM_51_AWCACHE(AP_AXIMM_51_AWCACHE),
        .AP_AXIMM_51_AWPROT(AP_AXIMM_51_AWPROT),
        .AP_AXIMM_51_AWREGION(AP_AXIMM_51_AWREGION),
        .AP_AXIMM_51_AWQOS(AP_AXIMM_51_AWQOS),
        .AP_AXIMM_51_AWVALID(AP_AXIMM_51_AWVALID),
        .AP_AXIMM_51_AWREADY(AP_AXIMM_51_AWREADY),
        .AP_AXIMM_51_WDATA(AP_AXIMM_51_WDATA),
        .AP_AXIMM_51_WSTRB(AP_AXIMM_51_WSTRB),
        .AP_AXIMM_51_WLAST(AP_AXIMM_51_WLAST),
        .AP_AXIMM_51_WVALID(AP_AXIMM_51_WVALID),
        .AP_AXIMM_51_WREADY(AP_AXIMM_51_WREADY),
        .AP_AXIMM_51_BRESP(AP_AXIMM_51_BRESP),
        .AP_AXIMM_51_BVALID(AP_AXIMM_51_BVALID),
        .AP_AXIMM_51_BREADY(AP_AXIMM_51_BREADY),
        .AP_AXIMM_51_ARADDR(AP_AXIMM_51_ARADDR),
        .AP_AXIMM_51_ARLEN(AP_AXIMM_51_ARLEN),
        .AP_AXIMM_51_ARSIZE(AP_AXIMM_51_ARSIZE),
        .AP_AXIMM_51_ARBURST(AP_AXIMM_51_ARBURST),
        .AP_AXIMM_51_ARLOCK(AP_AXIMM_51_ARLOCK),
        .AP_AXIMM_51_ARCACHE(AP_AXIMM_51_ARCACHE),
        .AP_AXIMM_51_ARPROT(AP_AXIMM_51_ARPROT),
        .AP_AXIMM_51_ARREGION(AP_AXIMM_51_ARREGION),
        .AP_AXIMM_51_ARQOS(AP_AXIMM_51_ARQOS),
        .AP_AXIMM_51_ARVALID(AP_AXIMM_51_ARVALID),
        .AP_AXIMM_51_ARREADY(AP_AXIMM_51_ARREADY),
        .AP_AXIMM_51_RDATA(AP_AXIMM_51_RDATA),
        .AP_AXIMM_51_RRESP(AP_AXIMM_51_RRESP),
        .AP_AXIMM_51_RLAST(AP_AXIMM_51_RLAST),
        .AP_AXIMM_51_RVALID(AP_AXIMM_51_RVALID),
        .AP_AXIMM_51_RREADY(AP_AXIMM_51_RREADY),
        .M_AXIMM_51_AWADDR(M_AXIMM_51_AWADDR),
        .M_AXIMM_51_AWLEN(M_AXIMM_51_AWLEN),
        .M_AXIMM_51_AWSIZE(M_AXIMM_51_AWSIZE),
        .M_AXIMM_51_AWBURST(M_AXIMM_51_AWBURST),
        .M_AXIMM_51_AWLOCK(M_AXIMM_51_AWLOCK),
        .M_AXIMM_51_AWCACHE(M_AXIMM_51_AWCACHE),
        .M_AXIMM_51_AWPROT(M_AXIMM_51_AWPROT),
        .M_AXIMM_51_AWREGION(M_AXIMM_51_AWREGION),
        .M_AXIMM_51_AWQOS(M_AXIMM_51_AWQOS),
        .M_AXIMM_51_AWVALID(M_AXIMM_51_AWVALID),
        .M_AXIMM_51_AWREADY(M_AXIMM_51_AWREADY),
        .M_AXIMM_51_WDATA(M_AXIMM_51_WDATA),
        .M_AXIMM_51_WSTRB(M_AXIMM_51_WSTRB),
        .M_AXIMM_51_WLAST(M_AXIMM_51_WLAST),
        .M_AXIMM_51_WVALID(M_AXIMM_51_WVALID),
        .M_AXIMM_51_WREADY(M_AXIMM_51_WREADY),
        .M_AXIMM_51_BRESP(M_AXIMM_51_BRESP),
        .M_AXIMM_51_BVALID(M_AXIMM_51_BVALID),
        .M_AXIMM_51_BREADY(M_AXIMM_51_BREADY),
        .M_AXIMM_51_ARADDR(M_AXIMM_51_ARADDR),
        .M_AXIMM_51_ARLEN(M_AXIMM_51_ARLEN),
        .M_AXIMM_51_ARSIZE(M_AXIMM_51_ARSIZE),
        .M_AXIMM_51_ARBURST(M_AXIMM_51_ARBURST),
        .M_AXIMM_51_ARLOCK(M_AXIMM_51_ARLOCK),
        .M_AXIMM_51_ARCACHE(M_AXIMM_51_ARCACHE),
        .M_AXIMM_51_ARPROT(M_AXIMM_51_ARPROT),
        .M_AXIMM_51_ARREGION(M_AXIMM_51_ARREGION),
        .M_AXIMM_51_ARQOS(M_AXIMM_51_ARQOS),
        .M_AXIMM_51_ARVALID(M_AXIMM_51_ARVALID),
        .M_AXIMM_51_ARREADY(M_AXIMM_51_ARREADY),
        .M_AXIMM_51_RDATA(M_AXIMM_51_RDATA),
        .M_AXIMM_51_RRESP(M_AXIMM_51_RRESP),
        .M_AXIMM_51_RLAST(M_AXIMM_51_RLAST),
        .M_AXIMM_51_RVALID(M_AXIMM_51_RVALID),
        .M_AXIMM_51_RREADY(M_AXIMM_51_RREADY),
        .AP_AXIMM_52_AWADDR(AP_AXIMM_52_AWADDR),
        .AP_AXIMM_52_AWLEN(AP_AXIMM_52_AWLEN),
        .AP_AXIMM_52_AWSIZE(AP_AXIMM_52_AWSIZE),
        .AP_AXIMM_52_AWBURST(AP_AXIMM_52_AWBURST),
        .AP_AXIMM_52_AWLOCK(AP_AXIMM_52_AWLOCK),
        .AP_AXIMM_52_AWCACHE(AP_AXIMM_52_AWCACHE),
        .AP_AXIMM_52_AWPROT(AP_AXIMM_52_AWPROT),
        .AP_AXIMM_52_AWREGION(AP_AXIMM_52_AWREGION),
        .AP_AXIMM_52_AWQOS(AP_AXIMM_52_AWQOS),
        .AP_AXIMM_52_AWVALID(AP_AXIMM_52_AWVALID),
        .AP_AXIMM_52_AWREADY(AP_AXIMM_52_AWREADY),
        .AP_AXIMM_52_WDATA(AP_AXIMM_52_WDATA),
        .AP_AXIMM_52_WSTRB(AP_AXIMM_52_WSTRB),
        .AP_AXIMM_52_WLAST(AP_AXIMM_52_WLAST),
        .AP_AXIMM_52_WVALID(AP_AXIMM_52_WVALID),
        .AP_AXIMM_52_WREADY(AP_AXIMM_52_WREADY),
        .AP_AXIMM_52_BRESP(AP_AXIMM_52_BRESP),
        .AP_AXIMM_52_BVALID(AP_AXIMM_52_BVALID),
        .AP_AXIMM_52_BREADY(AP_AXIMM_52_BREADY),
        .AP_AXIMM_52_ARADDR(AP_AXIMM_52_ARADDR),
        .AP_AXIMM_52_ARLEN(AP_AXIMM_52_ARLEN),
        .AP_AXIMM_52_ARSIZE(AP_AXIMM_52_ARSIZE),
        .AP_AXIMM_52_ARBURST(AP_AXIMM_52_ARBURST),
        .AP_AXIMM_52_ARLOCK(AP_AXIMM_52_ARLOCK),
        .AP_AXIMM_52_ARCACHE(AP_AXIMM_52_ARCACHE),
        .AP_AXIMM_52_ARPROT(AP_AXIMM_52_ARPROT),
        .AP_AXIMM_52_ARREGION(AP_AXIMM_52_ARREGION),
        .AP_AXIMM_52_ARQOS(AP_AXIMM_52_ARQOS),
        .AP_AXIMM_52_ARVALID(AP_AXIMM_52_ARVALID),
        .AP_AXIMM_52_ARREADY(AP_AXIMM_52_ARREADY),
        .AP_AXIMM_52_RDATA(AP_AXIMM_52_RDATA),
        .AP_AXIMM_52_RRESP(AP_AXIMM_52_RRESP),
        .AP_AXIMM_52_RLAST(AP_AXIMM_52_RLAST),
        .AP_AXIMM_52_RVALID(AP_AXIMM_52_RVALID),
        .AP_AXIMM_52_RREADY(AP_AXIMM_52_RREADY),
        .M_AXIMM_52_AWADDR(M_AXIMM_52_AWADDR),
        .M_AXIMM_52_AWLEN(M_AXIMM_52_AWLEN),
        .M_AXIMM_52_AWSIZE(M_AXIMM_52_AWSIZE),
        .M_AXIMM_52_AWBURST(M_AXIMM_52_AWBURST),
        .M_AXIMM_52_AWLOCK(M_AXIMM_52_AWLOCK),
        .M_AXIMM_52_AWCACHE(M_AXIMM_52_AWCACHE),
        .M_AXIMM_52_AWPROT(M_AXIMM_52_AWPROT),
        .M_AXIMM_52_AWREGION(M_AXIMM_52_AWREGION),
        .M_AXIMM_52_AWQOS(M_AXIMM_52_AWQOS),
        .M_AXIMM_52_AWVALID(M_AXIMM_52_AWVALID),
        .M_AXIMM_52_AWREADY(M_AXIMM_52_AWREADY),
        .M_AXIMM_52_WDATA(M_AXIMM_52_WDATA),
        .M_AXIMM_52_WSTRB(M_AXIMM_52_WSTRB),
        .M_AXIMM_52_WLAST(M_AXIMM_52_WLAST),
        .M_AXIMM_52_WVALID(M_AXIMM_52_WVALID),
        .M_AXIMM_52_WREADY(M_AXIMM_52_WREADY),
        .M_AXIMM_52_BRESP(M_AXIMM_52_BRESP),
        .M_AXIMM_52_BVALID(M_AXIMM_52_BVALID),
        .M_AXIMM_52_BREADY(M_AXIMM_52_BREADY),
        .M_AXIMM_52_ARADDR(M_AXIMM_52_ARADDR),
        .M_AXIMM_52_ARLEN(M_AXIMM_52_ARLEN),
        .M_AXIMM_52_ARSIZE(M_AXIMM_52_ARSIZE),
        .M_AXIMM_52_ARBURST(M_AXIMM_52_ARBURST),
        .M_AXIMM_52_ARLOCK(M_AXIMM_52_ARLOCK),
        .M_AXIMM_52_ARCACHE(M_AXIMM_52_ARCACHE),
        .M_AXIMM_52_ARPROT(M_AXIMM_52_ARPROT),
        .M_AXIMM_52_ARREGION(M_AXIMM_52_ARREGION),
        .M_AXIMM_52_ARQOS(M_AXIMM_52_ARQOS),
        .M_AXIMM_52_ARVALID(M_AXIMM_52_ARVALID),
        .M_AXIMM_52_ARREADY(M_AXIMM_52_ARREADY),
        .M_AXIMM_52_RDATA(M_AXIMM_52_RDATA),
        .M_AXIMM_52_RRESP(M_AXIMM_52_RRESP),
        .M_AXIMM_52_RLAST(M_AXIMM_52_RLAST),
        .M_AXIMM_52_RVALID(M_AXIMM_52_RVALID),
        .M_AXIMM_52_RREADY(M_AXIMM_52_RREADY),
        .AP_AXIMM_53_AWADDR(AP_AXIMM_53_AWADDR),
        .AP_AXIMM_53_AWLEN(AP_AXIMM_53_AWLEN),
        .AP_AXIMM_53_AWSIZE(AP_AXIMM_53_AWSIZE),
        .AP_AXIMM_53_AWBURST(AP_AXIMM_53_AWBURST),
        .AP_AXIMM_53_AWLOCK(AP_AXIMM_53_AWLOCK),
        .AP_AXIMM_53_AWCACHE(AP_AXIMM_53_AWCACHE),
        .AP_AXIMM_53_AWPROT(AP_AXIMM_53_AWPROT),
        .AP_AXIMM_53_AWREGION(AP_AXIMM_53_AWREGION),
        .AP_AXIMM_53_AWQOS(AP_AXIMM_53_AWQOS),
        .AP_AXIMM_53_AWVALID(AP_AXIMM_53_AWVALID),
        .AP_AXIMM_53_AWREADY(AP_AXIMM_53_AWREADY),
        .AP_AXIMM_53_WDATA(AP_AXIMM_53_WDATA),
        .AP_AXIMM_53_WSTRB(AP_AXIMM_53_WSTRB),
        .AP_AXIMM_53_WLAST(AP_AXIMM_53_WLAST),
        .AP_AXIMM_53_WVALID(AP_AXIMM_53_WVALID),
        .AP_AXIMM_53_WREADY(AP_AXIMM_53_WREADY),
        .AP_AXIMM_53_BRESP(AP_AXIMM_53_BRESP),
        .AP_AXIMM_53_BVALID(AP_AXIMM_53_BVALID),
        .AP_AXIMM_53_BREADY(AP_AXIMM_53_BREADY),
        .AP_AXIMM_53_ARADDR(AP_AXIMM_53_ARADDR),
        .AP_AXIMM_53_ARLEN(AP_AXIMM_53_ARLEN),
        .AP_AXIMM_53_ARSIZE(AP_AXIMM_53_ARSIZE),
        .AP_AXIMM_53_ARBURST(AP_AXIMM_53_ARBURST),
        .AP_AXIMM_53_ARLOCK(AP_AXIMM_53_ARLOCK),
        .AP_AXIMM_53_ARCACHE(AP_AXIMM_53_ARCACHE),
        .AP_AXIMM_53_ARPROT(AP_AXIMM_53_ARPROT),
        .AP_AXIMM_53_ARREGION(AP_AXIMM_53_ARREGION),
        .AP_AXIMM_53_ARQOS(AP_AXIMM_53_ARQOS),
        .AP_AXIMM_53_ARVALID(AP_AXIMM_53_ARVALID),
        .AP_AXIMM_53_ARREADY(AP_AXIMM_53_ARREADY),
        .AP_AXIMM_53_RDATA(AP_AXIMM_53_RDATA),
        .AP_AXIMM_53_RRESP(AP_AXIMM_53_RRESP),
        .AP_AXIMM_53_RLAST(AP_AXIMM_53_RLAST),
        .AP_AXIMM_53_RVALID(AP_AXIMM_53_RVALID),
        .AP_AXIMM_53_RREADY(AP_AXIMM_53_RREADY),
        .M_AXIMM_53_AWADDR(M_AXIMM_53_AWADDR),
        .M_AXIMM_53_AWLEN(M_AXIMM_53_AWLEN),
        .M_AXIMM_53_AWSIZE(M_AXIMM_53_AWSIZE),
        .M_AXIMM_53_AWBURST(M_AXIMM_53_AWBURST),
        .M_AXIMM_53_AWLOCK(M_AXIMM_53_AWLOCK),
        .M_AXIMM_53_AWCACHE(M_AXIMM_53_AWCACHE),
        .M_AXIMM_53_AWPROT(M_AXIMM_53_AWPROT),
        .M_AXIMM_53_AWREGION(M_AXIMM_53_AWREGION),
        .M_AXIMM_53_AWQOS(M_AXIMM_53_AWQOS),
        .M_AXIMM_53_AWVALID(M_AXIMM_53_AWVALID),
        .M_AXIMM_53_AWREADY(M_AXIMM_53_AWREADY),
        .M_AXIMM_53_WDATA(M_AXIMM_53_WDATA),
        .M_AXIMM_53_WSTRB(M_AXIMM_53_WSTRB),
        .M_AXIMM_53_WLAST(M_AXIMM_53_WLAST),
        .M_AXIMM_53_WVALID(M_AXIMM_53_WVALID),
        .M_AXIMM_53_WREADY(M_AXIMM_53_WREADY),
        .M_AXIMM_53_BRESP(M_AXIMM_53_BRESP),
        .M_AXIMM_53_BVALID(M_AXIMM_53_BVALID),
        .M_AXIMM_53_BREADY(M_AXIMM_53_BREADY),
        .M_AXIMM_53_ARADDR(M_AXIMM_53_ARADDR),
        .M_AXIMM_53_ARLEN(M_AXIMM_53_ARLEN),
        .M_AXIMM_53_ARSIZE(M_AXIMM_53_ARSIZE),
        .M_AXIMM_53_ARBURST(M_AXIMM_53_ARBURST),
        .M_AXIMM_53_ARLOCK(M_AXIMM_53_ARLOCK),
        .M_AXIMM_53_ARCACHE(M_AXIMM_53_ARCACHE),
        .M_AXIMM_53_ARPROT(M_AXIMM_53_ARPROT),
        .M_AXIMM_53_ARREGION(M_AXIMM_53_ARREGION),
        .M_AXIMM_53_ARQOS(M_AXIMM_53_ARQOS),
        .M_AXIMM_53_ARVALID(M_AXIMM_53_ARVALID),
        .M_AXIMM_53_ARREADY(M_AXIMM_53_ARREADY),
        .M_AXIMM_53_RDATA(M_AXIMM_53_RDATA),
        .M_AXIMM_53_RRESP(M_AXIMM_53_RRESP),
        .M_AXIMM_53_RLAST(M_AXIMM_53_RLAST),
        .M_AXIMM_53_RVALID(M_AXIMM_53_RVALID),
        .M_AXIMM_53_RREADY(M_AXIMM_53_RREADY),
        .AP_AXIMM_54_AWADDR(AP_AXIMM_54_AWADDR),
        .AP_AXIMM_54_AWLEN(AP_AXIMM_54_AWLEN),
        .AP_AXIMM_54_AWSIZE(AP_AXIMM_54_AWSIZE),
        .AP_AXIMM_54_AWBURST(AP_AXIMM_54_AWBURST),
        .AP_AXIMM_54_AWLOCK(AP_AXIMM_54_AWLOCK),
        .AP_AXIMM_54_AWCACHE(AP_AXIMM_54_AWCACHE),
        .AP_AXIMM_54_AWPROT(AP_AXIMM_54_AWPROT),
        .AP_AXIMM_54_AWREGION(AP_AXIMM_54_AWREGION),
        .AP_AXIMM_54_AWQOS(AP_AXIMM_54_AWQOS),
        .AP_AXIMM_54_AWVALID(AP_AXIMM_54_AWVALID),
        .AP_AXIMM_54_AWREADY(AP_AXIMM_54_AWREADY),
        .AP_AXIMM_54_WDATA(AP_AXIMM_54_WDATA),
        .AP_AXIMM_54_WSTRB(AP_AXIMM_54_WSTRB),
        .AP_AXIMM_54_WLAST(AP_AXIMM_54_WLAST),
        .AP_AXIMM_54_WVALID(AP_AXIMM_54_WVALID),
        .AP_AXIMM_54_WREADY(AP_AXIMM_54_WREADY),
        .AP_AXIMM_54_BRESP(AP_AXIMM_54_BRESP),
        .AP_AXIMM_54_BVALID(AP_AXIMM_54_BVALID),
        .AP_AXIMM_54_BREADY(AP_AXIMM_54_BREADY),
        .AP_AXIMM_54_ARADDR(AP_AXIMM_54_ARADDR),
        .AP_AXIMM_54_ARLEN(AP_AXIMM_54_ARLEN),
        .AP_AXIMM_54_ARSIZE(AP_AXIMM_54_ARSIZE),
        .AP_AXIMM_54_ARBURST(AP_AXIMM_54_ARBURST),
        .AP_AXIMM_54_ARLOCK(AP_AXIMM_54_ARLOCK),
        .AP_AXIMM_54_ARCACHE(AP_AXIMM_54_ARCACHE),
        .AP_AXIMM_54_ARPROT(AP_AXIMM_54_ARPROT),
        .AP_AXIMM_54_ARREGION(AP_AXIMM_54_ARREGION),
        .AP_AXIMM_54_ARQOS(AP_AXIMM_54_ARQOS),
        .AP_AXIMM_54_ARVALID(AP_AXIMM_54_ARVALID),
        .AP_AXIMM_54_ARREADY(AP_AXIMM_54_ARREADY),
        .AP_AXIMM_54_RDATA(AP_AXIMM_54_RDATA),
        .AP_AXIMM_54_RRESP(AP_AXIMM_54_RRESP),
        .AP_AXIMM_54_RLAST(AP_AXIMM_54_RLAST),
        .AP_AXIMM_54_RVALID(AP_AXIMM_54_RVALID),
        .AP_AXIMM_54_RREADY(AP_AXIMM_54_RREADY),
        .M_AXIMM_54_AWADDR(M_AXIMM_54_AWADDR),
        .M_AXIMM_54_AWLEN(M_AXIMM_54_AWLEN),
        .M_AXIMM_54_AWSIZE(M_AXIMM_54_AWSIZE),
        .M_AXIMM_54_AWBURST(M_AXIMM_54_AWBURST),
        .M_AXIMM_54_AWLOCK(M_AXIMM_54_AWLOCK),
        .M_AXIMM_54_AWCACHE(M_AXIMM_54_AWCACHE),
        .M_AXIMM_54_AWPROT(M_AXIMM_54_AWPROT),
        .M_AXIMM_54_AWREGION(M_AXIMM_54_AWREGION),
        .M_AXIMM_54_AWQOS(M_AXIMM_54_AWQOS),
        .M_AXIMM_54_AWVALID(M_AXIMM_54_AWVALID),
        .M_AXIMM_54_AWREADY(M_AXIMM_54_AWREADY),
        .M_AXIMM_54_WDATA(M_AXIMM_54_WDATA),
        .M_AXIMM_54_WSTRB(M_AXIMM_54_WSTRB),
        .M_AXIMM_54_WLAST(M_AXIMM_54_WLAST),
        .M_AXIMM_54_WVALID(M_AXIMM_54_WVALID),
        .M_AXIMM_54_WREADY(M_AXIMM_54_WREADY),
        .M_AXIMM_54_BRESP(M_AXIMM_54_BRESP),
        .M_AXIMM_54_BVALID(M_AXIMM_54_BVALID),
        .M_AXIMM_54_BREADY(M_AXIMM_54_BREADY),
        .M_AXIMM_54_ARADDR(M_AXIMM_54_ARADDR),
        .M_AXIMM_54_ARLEN(M_AXIMM_54_ARLEN),
        .M_AXIMM_54_ARSIZE(M_AXIMM_54_ARSIZE),
        .M_AXIMM_54_ARBURST(M_AXIMM_54_ARBURST),
        .M_AXIMM_54_ARLOCK(M_AXIMM_54_ARLOCK),
        .M_AXIMM_54_ARCACHE(M_AXIMM_54_ARCACHE),
        .M_AXIMM_54_ARPROT(M_AXIMM_54_ARPROT),
        .M_AXIMM_54_ARREGION(M_AXIMM_54_ARREGION),
        .M_AXIMM_54_ARQOS(M_AXIMM_54_ARQOS),
        .M_AXIMM_54_ARVALID(M_AXIMM_54_ARVALID),
        .M_AXIMM_54_ARREADY(M_AXIMM_54_ARREADY),
        .M_AXIMM_54_RDATA(M_AXIMM_54_RDATA),
        .M_AXIMM_54_RRESP(M_AXIMM_54_RRESP),
        .M_AXIMM_54_RLAST(M_AXIMM_54_RLAST),
        .M_AXIMM_54_RVALID(M_AXIMM_54_RVALID),
        .M_AXIMM_54_RREADY(M_AXIMM_54_RREADY),
        .AP_AXIMM_55_AWADDR(AP_AXIMM_55_AWADDR),
        .AP_AXIMM_55_AWLEN(AP_AXIMM_55_AWLEN),
        .AP_AXIMM_55_AWSIZE(AP_AXIMM_55_AWSIZE),
        .AP_AXIMM_55_AWBURST(AP_AXIMM_55_AWBURST),
        .AP_AXIMM_55_AWLOCK(AP_AXIMM_55_AWLOCK),
        .AP_AXIMM_55_AWCACHE(AP_AXIMM_55_AWCACHE),
        .AP_AXIMM_55_AWPROT(AP_AXIMM_55_AWPROT),
        .AP_AXIMM_55_AWREGION(AP_AXIMM_55_AWREGION),
        .AP_AXIMM_55_AWQOS(AP_AXIMM_55_AWQOS),
        .AP_AXIMM_55_AWVALID(AP_AXIMM_55_AWVALID),
        .AP_AXIMM_55_AWREADY(AP_AXIMM_55_AWREADY),
        .AP_AXIMM_55_WDATA(AP_AXIMM_55_WDATA),
        .AP_AXIMM_55_WSTRB(AP_AXIMM_55_WSTRB),
        .AP_AXIMM_55_WLAST(AP_AXIMM_55_WLAST),
        .AP_AXIMM_55_WVALID(AP_AXIMM_55_WVALID),
        .AP_AXIMM_55_WREADY(AP_AXIMM_55_WREADY),
        .AP_AXIMM_55_BRESP(AP_AXIMM_55_BRESP),
        .AP_AXIMM_55_BVALID(AP_AXIMM_55_BVALID),
        .AP_AXIMM_55_BREADY(AP_AXIMM_55_BREADY),
        .AP_AXIMM_55_ARADDR(AP_AXIMM_55_ARADDR),
        .AP_AXIMM_55_ARLEN(AP_AXIMM_55_ARLEN),
        .AP_AXIMM_55_ARSIZE(AP_AXIMM_55_ARSIZE),
        .AP_AXIMM_55_ARBURST(AP_AXIMM_55_ARBURST),
        .AP_AXIMM_55_ARLOCK(AP_AXIMM_55_ARLOCK),
        .AP_AXIMM_55_ARCACHE(AP_AXIMM_55_ARCACHE),
        .AP_AXIMM_55_ARPROT(AP_AXIMM_55_ARPROT),
        .AP_AXIMM_55_ARREGION(AP_AXIMM_55_ARREGION),
        .AP_AXIMM_55_ARQOS(AP_AXIMM_55_ARQOS),
        .AP_AXIMM_55_ARVALID(AP_AXIMM_55_ARVALID),
        .AP_AXIMM_55_ARREADY(AP_AXIMM_55_ARREADY),
        .AP_AXIMM_55_RDATA(AP_AXIMM_55_RDATA),
        .AP_AXIMM_55_RRESP(AP_AXIMM_55_RRESP),
        .AP_AXIMM_55_RLAST(AP_AXIMM_55_RLAST),
        .AP_AXIMM_55_RVALID(AP_AXIMM_55_RVALID),
        .AP_AXIMM_55_RREADY(AP_AXIMM_55_RREADY),
        .M_AXIMM_55_AWADDR(M_AXIMM_55_AWADDR),
        .M_AXIMM_55_AWLEN(M_AXIMM_55_AWLEN),
        .M_AXIMM_55_AWSIZE(M_AXIMM_55_AWSIZE),
        .M_AXIMM_55_AWBURST(M_AXIMM_55_AWBURST),
        .M_AXIMM_55_AWLOCK(M_AXIMM_55_AWLOCK),
        .M_AXIMM_55_AWCACHE(M_AXIMM_55_AWCACHE),
        .M_AXIMM_55_AWPROT(M_AXIMM_55_AWPROT),
        .M_AXIMM_55_AWREGION(M_AXIMM_55_AWREGION),
        .M_AXIMM_55_AWQOS(M_AXIMM_55_AWQOS),
        .M_AXIMM_55_AWVALID(M_AXIMM_55_AWVALID),
        .M_AXIMM_55_AWREADY(M_AXIMM_55_AWREADY),
        .M_AXIMM_55_WDATA(M_AXIMM_55_WDATA),
        .M_AXIMM_55_WSTRB(M_AXIMM_55_WSTRB),
        .M_AXIMM_55_WLAST(M_AXIMM_55_WLAST),
        .M_AXIMM_55_WVALID(M_AXIMM_55_WVALID),
        .M_AXIMM_55_WREADY(M_AXIMM_55_WREADY),
        .M_AXIMM_55_BRESP(M_AXIMM_55_BRESP),
        .M_AXIMM_55_BVALID(M_AXIMM_55_BVALID),
        .M_AXIMM_55_BREADY(M_AXIMM_55_BREADY),
        .M_AXIMM_55_ARADDR(M_AXIMM_55_ARADDR),
        .M_AXIMM_55_ARLEN(M_AXIMM_55_ARLEN),
        .M_AXIMM_55_ARSIZE(M_AXIMM_55_ARSIZE),
        .M_AXIMM_55_ARBURST(M_AXIMM_55_ARBURST),
        .M_AXIMM_55_ARLOCK(M_AXIMM_55_ARLOCK),
        .M_AXIMM_55_ARCACHE(M_AXIMM_55_ARCACHE),
        .M_AXIMM_55_ARPROT(M_AXIMM_55_ARPROT),
        .M_AXIMM_55_ARREGION(M_AXIMM_55_ARREGION),
        .M_AXIMM_55_ARQOS(M_AXIMM_55_ARQOS),
        .M_AXIMM_55_ARVALID(M_AXIMM_55_ARVALID),
        .M_AXIMM_55_ARREADY(M_AXIMM_55_ARREADY),
        .M_AXIMM_55_RDATA(M_AXIMM_55_RDATA),
        .M_AXIMM_55_RRESP(M_AXIMM_55_RRESP),
        .M_AXIMM_55_RLAST(M_AXIMM_55_RLAST),
        .M_AXIMM_55_RVALID(M_AXIMM_55_RVALID),
        .M_AXIMM_55_RREADY(M_AXIMM_55_RREADY),
        .AP_AXIMM_56_AWADDR(AP_AXIMM_56_AWADDR),
        .AP_AXIMM_56_AWLEN(AP_AXIMM_56_AWLEN),
        .AP_AXIMM_56_AWSIZE(AP_AXIMM_56_AWSIZE),
        .AP_AXIMM_56_AWBURST(AP_AXIMM_56_AWBURST),
        .AP_AXIMM_56_AWLOCK(AP_AXIMM_56_AWLOCK),
        .AP_AXIMM_56_AWCACHE(AP_AXIMM_56_AWCACHE),
        .AP_AXIMM_56_AWPROT(AP_AXIMM_56_AWPROT),
        .AP_AXIMM_56_AWREGION(AP_AXIMM_56_AWREGION),
        .AP_AXIMM_56_AWQOS(AP_AXIMM_56_AWQOS),
        .AP_AXIMM_56_AWVALID(AP_AXIMM_56_AWVALID),
        .AP_AXIMM_56_AWREADY(AP_AXIMM_56_AWREADY),
        .AP_AXIMM_56_WDATA(AP_AXIMM_56_WDATA),
        .AP_AXIMM_56_WSTRB(AP_AXIMM_56_WSTRB),
        .AP_AXIMM_56_WLAST(AP_AXIMM_56_WLAST),
        .AP_AXIMM_56_WVALID(AP_AXIMM_56_WVALID),
        .AP_AXIMM_56_WREADY(AP_AXIMM_56_WREADY),
        .AP_AXIMM_56_BRESP(AP_AXIMM_56_BRESP),
        .AP_AXIMM_56_BVALID(AP_AXIMM_56_BVALID),
        .AP_AXIMM_56_BREADY(AP_AXIMM_56_BREADY),
        .AP_AXIMM_56_ARADDR(AP_AXIMM_56_ARADDR),
        .AP_AXIMM_56_ARLEN(AP_AXIMM_56_ARLEN),
        .AP_AXIMM_56_ARSIZE(AP_AXIMM_56_ARSIZE),
        .AP_AXIMM_56_ARBURST(AP_AXIMM_56_ARBURST),
        .AP_AXIMM_56_ARLOCK(AP_AXIMM_56_ARLOCK),
        .AP_AXIMM_56_ARCACHE(AP_AXIMM_56_ARCACHE),
        .AP_AXIMM_56_ARPROT(AP_AXIMM_56_ARPROT),
        .AP_AXIMM_56_ARREGION(AP_AXIMM_56_ARREGION),
        .AP_AXIMM_56_ARQOS(AP_AXIMM_56_ARQOS),
        .AP_AXIMM_56_ARVALID(AP_AXIMM_56_ARVALID),
        .AP_AXIMM_56_ARREADY(AP_AXIMM_56_ARREADY),
        .AP_AXIMM_56_RDATA(AP_AXIMM_56_RDATA),
        .AP_AXIMM_56_RRESP(AP_AXIMM_56_RRESP),
        .AP_AXIMM_56_RLAST(AP_AXIMM_56_RLAST),
        .AP_AXIMM_56_RVALID(AP_AXIMM_56_RVALID),
        .AP_AXIMM_56_RREADY(AP_AXIMM_56_RREADY),
        .M_AXIMM_56_AWADDR(M_AXIMM_56_AWADDR),
        .M_AXIMM_56_AWLEN(M_AXIMM_56_AWLEN),
        .M_AXIMM_56_AWSIZE(M_AXIMM_56_AWSIZE),
        .M_AXIMM_56_AWBURST(M_AXIMM_56_AWBURST),
        .M_AXIMM_56_AWLOCK(M_AXIMM_56_AWLOCK),
        .M_AXIMM_56_AWCACHE(M_AXIMM_56_AWCACHE),
        .M_AXIMM_56_AWPROT(M_AXIMM_56_AWPROT),
        .M_AXIMM_56_AWREGION(M_AXIMM_56_AWREGION),
        .M_AXIMM_56_AWQOS(M_AXIMM_56_AWQOS),
        .M_AXIMM_56_AWVALID(M_AXIMM_56_AWVALID),
        .M_AXIMM_56_AWREADY(M_AXIMM_56_AWREADY),
        .M_AXIMM_56_WDATA(M_AXIMM_56_WDATA),
        .M_AXIMM_56_WSTRB(M_AXIMM_56_WSTRB),
        .M_AXIMM_56_WLAST(M_AXIMM_56_WLAST),
        .M_AXIMM_56_WVALID(M_AXIMM_56_WVALID),
        .M_AXIMM_56_WREADY(M_AXIMM_56_WREADY),
        .M_AXIMM_56_BRESP(M_AXIMM_56_BRESP),
        .M_AXIMM_56_BVALID(M_AXIMM_56_BVALID),
        .M_AXIMM_56_BREADY(M_AXIMM_56_BREADY),
        .M_AXIMM_56_ARADDR(M_AXIMM_56_ARADDR),
        .M_AXIMM_56_ARLEN(M_AXIMM_56_ARLEN),
        .M_AXIMM_56_ARSIZE(M_AXIMM_56_ARSIZE),
        .M_AXIMM_56_ARBURST(M_AXIMM_56_ARBURST),
        .M_AXIMM_56_ARLOCK(M_AXIMM_56_ARLOCK),
        .M_AXIMM_56_ARCACHE(M_AXIMM_56_ARCACHE),
        .M_AXIMM_56_ARPROT(M_AXIMM_56_ARPROT),
        .M_AXIMM_56_ARREGION(M_AXIMM_56_ARREGION),
        .M_AXIMM_56_ARQOS(M_AXIMM_56_ARQOS),
        .M_AXIMM_56_ARVALID(M_AXIMM_56_ARVALID),
        .M_AXIMM_56_ARREADY(M_AXIMM_56_ARREADY),
        .M_AXIMM_56_RDATA(M_AXIMM_56_RDATA),
        .M_AXIMM_56_RRESP(M_AXIMM_56_RRESP),
        .M_AXIMM_56_RLAST(M_AXIMM_56_RLAST),
        .M_AXIMM_56_RVALID(M_AXIMM_56_RVALID),
        .M_AXIMM_56_RREADY(M_AXIMM_56_RREADY),
        .AP_AXIMM_57_AWADDR(AP_AXIMM_57_AWADDR),
        .AP_AXIMM_57_AWLEN(AP_AXIMM_57_AWLEN),
        .AP_AXIMM_57_AWSIZE(AP_AXIMM_57_AWSIZE),
        .AP_AXIMM_57_AWBURST(AP_AXIMM_57_AWBURST),
        .AP_AXIMM_57_AWLOCK(AP_AXIMM_57_AWLOCK),
        .AP_AXIMM_57_AWCACHE(AP_AXIMM_57_AWCACHE),
        .AP_AXIMM_57_AWPROT(AP_AXIMM_57_AWPROT),
        .AP_AXIMM_57_AWREGION(AP_AXIMM_57_AWREGION),
        .AP_AXIMM_57_AWQOS(AP_AXIMM_57_AWQOS),
        .AP_AXIMM_57_AWVALID(AP_AXIMM_57_AWVALID),
        .AP_AXIMM_57_AWREADY(AP_AXIMM_57_AWREADY),
        .AP_AXIMM_57_WDATA(AP_AXIMM_57_WDATA),
        .AP_AXIMM_57_WSTRB(AP_AXIMM_57_WSTRB),
        .AP_AXIMM_57_WLAST(AP_AXIMM_57_WLAST),
        .AP_AXIMM_57_WVALID(AP_AXIMM_57_WVALID),
        .AP_AXIMM_57_WREADY(AP_AXIMM_57_WREADY),
        .AP_AXIMM_57_BRESP(AP_AXIMM_57_BRESP),
        .AP_AXIMM_57_BVALID(AP_AXIMM_57_BVALID),
        .AP_AXIMM_57_BREADY(AP_AXIMM_57_BREADY),
        .AP_AXIMM_57_ARADDR(AP_AXIMM_57_ARADDR),
        .AP_AXIMM_57_ARLEN(AP_AXIMM_57_ARLEN),
        .AP_AXIMM_57_ARSIZE(AP_AXIMM_57_ARSIZE),
        .AP_AXIMM_57_ARBURST(AP_AXIMM_57_ARBURST),
        .AP_AXIMM_57_ARLOCK(AP_AXIMM_57_ARLOCK),
        .AP_AXIMM_57_ARCACHE(AP_AXIMM_57_ARCACHE),
        .AP_AXIMM_57_ARPROT(AP_AXIMM_57_ARPROT),
        .AP_AXIMM_57_ARREGION(AP_AXIMM_57_ARREGION),
        .AP_AXIMM_57_ARQOS(AP_AXIMM_57_ARQOS),
        .AP_AXIMM_57_ARVALID(AP_AXIMM_57_ARVALID),
        .AP_AXIMM_57_ARREADY(AP_AXIMM_57_ARREADY),
        .AP_AXIMM_57_RDATA(AP_AXIMM_57_RDATA),
        .AP_AXIMM_57_RRESP(AP_AXIMM_57_RRESP),
        .AP_AXIMM_57_RLAST(AP_AXIMM_57_RLAST),
        .AP_AXIMM_57_RVALID(AP_AXIMM_57_RVALID),
        .AP_AXIMM_57_RREADY(AP_AXIMM_57_RREADY),
        .M_AXIMM_57_AWADDR(M_AXIMM_57_AWADDR),
        .M_AXIMM_57_AWLEN(M_AXIMM_57_AWLEN),
        .M_AXIMM_57_AWSIZE(M_AXIMM_57_AWSIZE),
        .M_AXIMM_57_AWBURST(M_AXIMM_57_AWBURST),
        .M_AXIMM_57_AWLOCK(M_AXIMM_57_AWLOCK),
        .M_AXIMM_57_AWCACHE(M_AXIMM_57_AWCACHE),
        .M_AXIMM_57_AWPROT(M_AXIMM_57_AWPROT),
        .M_AXIMM_57_AWREGION(M_AXIMM_57_AWREGION),
        .M_AXIMM_57_AWQOS(M_AXIMM_57_AWQOS),
        .M_AXIMM_57_AWVALID(M_AXIMM_57_AWVALID),
        .M_AXIMM_57_AWREADY(M_AXIMM_57_AWREADY),
        .M_AXIMM_57_WDATA(M_AXIMM_57_WDATA),
        .M_AXIMM_57_WSTRB(M_AXIMM_57_WSTRB),
        .M_AXIMM_57_WLAST(M_AXIMM_57_WLAST),
        .M_AXIMM_57_WVALID(M_AXIMM_57_WVALID),
        .M_AXIMM_57_WREADY(M_AXIMM_57_WREADY),
        .M_AXIMM_57_BRESP(M_AXIMM_57_BRESP),
        .M_AXIMM_57_BVALID(M_AXIMM_57_BVALID),
        .M_AXIMM_57_BREADY(M_AXIMM_57_BREADY),
        .M_AXIMM_57_ARADDR(M_AXIMM_57_ARADDR),
        .M_AXIMM_57_ARLEN(M_AXIMM_57_ARLEN),
        .M_AXIMM_57_ARSIZE(M_AXIMM_57_ARSIZE),
        .M_AXIMM_57_ARBURST(M_AXIMM_57_ARBURST),
        .M_AXIMM_57_ARLOCK(M_AXIMM_57_ARLOCK),
        .M_AXIMM_57_ARCACHE(M_AXIMM_57_ARCACHE),
        .M_AXIMM_57_ARPROT(M_AXIMM_57_ARPROT),
        .M_AXIMM_57_ARREGION(M_AXIMM_57_ARREGION),
        .M_AXIMM_57_ARQOS(M_AXIMM_57_ARQOS),
        .M_AXIMM_57_ARVALID(M_AXIMM_57_ARVALID),
        .M_AXIMM_57_ARREADY(M_AXIMM_57_ARREADY),
        .M_AXIMM_57_RDATA(M_AXIMM_57_RDATA),
        .M_AXIMM_57_RRESP(M_AXIMM_57_RRESP),
        .M_AXIMM_57_RLAST(M_AXIMM_57_RLAST),
        .M_AXIMM_57_RVALID(M_AXIMM_57_RVALID),
        .M_AXIMM_57_RREADY(M_AXIMM_57_RREADY),
        .AP_AXIMM_58_AWADDR(AP_AXIMM_58_AWADDR),
        .AP_AXIMM_58_AWLEN(AP_AXIMM_58_AWLEN),
        .AP_AXIMM_58_AWSIZE(AP_AXIMM_58_AWSIZE),
        .AP_AXIMM_58_AWBURST(AP_AXIMM_58_AWBURST),
        .AP_AXIMM_58_AWLOCK(AP_AXIMM_58_AWLOCK),
        .AP_AXIMM_58_AWCACHE(AP_AXIMM_58_AWCACHE),
        .AP_AXIMM_58_AWPROT(AP_AXIMM_58_AWPROT),
        .AP_AXIMM_58_AWREGION(AP_AXIMM_58_AWREGION),
        .AP_AXIMM_58_AWQOS(AP_AXIMM_58_AWQOS),
        .AP_AXIMM_58_AWVALID(AP_AXIMM_58_AWVALID),
        .AP_AXIMM_58_AWREADY(AP_AXIMM_58_AWREADY),
        .AP_AXIMM_58_WDATA(AP_AXIMM_58_WDATA),
        .AP_AXIMM_58_WSTRB(AP_AXIMM_58_WSTRB),
        .AP_AXIMM_58_WLAST(AP_AXIMM_58_WLAST),
        .AP_AXIMM_58_WVALID(AP_AXIMM_58_WVALID),
        .AP_AXIMM_58_WREADY(AP_AXIMM_58_WREADY),
        .AP_AXIMM_58_BRESP(AP_AXIMM_58_BRESP),
        .AP_AXIMM_58_BVALID(AP_AXIMM_58_BVALID),
        .AP_AXIMM_58_BREADY(AP_AXIMM_58_BREADY),
        .AP_AXIMM_58_ARADDR(AP_AXIMM_58_ARADDR),
        .AP_AXIMM_58_ARLEN(AP_AXIMM_58_ARLEN),
        .AP_AXIMM_58_ARSIZE(AP_AXIMM_58_ARSIZE),
        .AP_AXIMM_58_ARBURST(AP_AXIMM_58_ARBURST),
        .AP_AXIMM_58_ARLOCK(AP_AXIMM_58_ARLOCK),
        .AP_AXIMM_58_ARCACHE(AP_AXIMM_58_ARCACHE),
        .AP_AXIMM_58_ARPROT(AP_AXIMM_58_ARPROT),
        .AP_AXIMM_58_ARREGION(AP_AXIMM_58_ARREGION),
        .AP_AXIMM_58_ARQOS(AP_AXIMM_58_ARQOS),
        .AP_AXIMM_58_ARVALID(AP_AXIMM_58_ARVALID),
        .AP_AXIMM_58_ARREADY(AP_AXIMM_58_ARREADY),
        .AP_AXIMM_58_RDATA(AP_AXIMM_58_RDATA),
        .AP_AXIMM_58_RRESP(AP_AXIMM_58_RRESP),
        .AP_AXIMM_58_RLAST(AP_AXIMM_58_RLAST),
        .AP_AXIMM_58_RVALID(AP_AXIMM_58_RVALID),
        .AP_AXIMM_58_RREADY(AP_AXIMM_58_RREADY),
        .M_AXIMM_58_AWADDR(M_AXIMM_58_AWADDR),
        .M_AXIMM_58_AWLEN(M_AXIMM_58_AWLEN),
        .M_AXIMM_58_AWSIZE(M_AXIMM_58_AWSIZE),
        .M_AXIMM_58_AWBURST(M_AXIMM_58_AWBURST),
        .M_AXIMM_58_AWLOCK(M_AXIMM_58_AWLOCK),
        .M_AXIMM_58_AWCACHE(M_AXIMM_58_AWCACHE),
        .M_AXIMM_58_AWPROT(M_AXIMM_58_AWPROT),
        .M_AXIMM_58_AWREGION(M_AXIMM_58_AWREGION),
        .M_AXIMM_58_AWQOS(M_AXIMM_58_AWQOS),
        .M_AXIMM_58_AWVALID(M_AXIMM_58_AWVALID),
        .M_AXIMM_58_AWREADY(M_AXIMM_58_AWREADY),
        .M_AXIMM_58_WDATA(M_AXIMM_58_WDATA),
        .M_AXIMM_58_WSTRB(M_AXIMM_58_WSTRB),
        .M_AXIMM_58_WLAST(M_AXIMM_58_WLAST),
        .M_AXIMM_58_WVALID(M_AXIMM_58_WVALID),
        .M_AXIMM_58_WREADY(M_AXIMM_58_WREADY),
        .M_AXIMM_58_BRESP(M_AXIMM_58_BRESP),
        .M_AXIMM_58_BVALID(M_AXIMM_58_BVALID),
        .M_AXIMM_58_BREADY(M_AXIMM_58_BREADY),
        .M_AXIMM_58_ARADDR(M_AXIMM_58_ARADDR),
        .M_AXIMM_58_ARLEN(M_AXIMM_58_ARLEN),
        .M_AXIMM_58_ARSIZE(M_AXIMM_58_ARSIZE),
        .M_AXIMM_58_ARBURST(M_AXIMM_58_ARBURST),
        .M_AXIMM_58_ARLOCK(M_AXIMM_58_ARLOCK),
        .M_AXIMM_58_ARCACHE(M_AXIMM_58_ARCACHE),
        .M_AXIMM_58_ARPROT(M_AXIMM_58_ARPROT),
        .M_AXIMM_58_ARREGION(M_AXIMM_58_ARREGION),
        .M_AXIMM_58_ARQOS(M_AXIMM_58_ARQOS),
        .M_AXIMM_58_ARVALID(M_AXIMM_58_ARVALID),
        .M_AXIMM_58_ARREADY(M_AXIMM_58_ARREADY),
        .M_AXIMM_58_RDATA(M_AXIMM_58_RDATA),
        .M_AXIMM_58_RRESP(M_AXIMM_58_RRESP),
        .M_AXIMM_58_RLAST(M_AXIMM_58_RLAST),
        .M_AXIMM_58_RVALID(M_AXIMM_58_RVALID),
        .M_AXIMM_58_RREADY(M_AXIMM_58_RREADY),
        .AP_AXIMM_59_AWADDR(AP_AXIMM_59_AWADDR),
        .AP_AXIMM_59_AWLEN(AP_AXIMM_59_AWLEN),
        .AP_AXIMM_59_AWSIZE(AP_AXIMM_59_AWSIZE),
        .AP_AXIMM_59_AWBURST(AP_AXIMM_59_AWBURST),
        .AP_AXIMM_59_AWLOCK(AP_AXIMM_59_AWLOCK),
        .AP_AXIMM_59_AWCACHE(AP_AXIMM_59_AWCACHE),
        .AP_AXIMM_59_AWPROT(AP_AXIMM_59_AWPROT),
        .AP_AXIMM_59_AWREGION(AP_AXIMM_59_AWREGION),
        .AP_AXIMM_59_AWQOS(AP_AXIMM_59_AWQOS),
        .AP_AXIMM_59_AWVALID(AP_AXIMM_59_AWVALID),
        .AP_AXIMM_59_AWREADY(AP_AXIMM_59_AWREADY),
        .AP_AXIMM_59_WDATA(AP_AXIMM_59_WDATA),
        .AP_AXIMM_59_WSTRB(AP_AXIMM_59_WSTRB),
        .AP_AXIMM_59_WLAST(AP_AXIMM_59_WLAST),
        .AP_AXIMM_59_WVALID(AP_AXIMM_59_WVALID),
        .AP_AXIMM_59_WREADY(AP_AXIMM_59_WREADY),
        .AP_AXIMM_59_BRESP(AP_AXIMM_59_BRESP),
        .AP_AXIMM_59_BVALID(AP_AXIMM_59_BVALID),
        .AP_AXIMM_59_BREADY(AP_AXIMM_59_BREADY),
        .AP_AXIMM_59_ARADDR(AP_AXIMM_59_ARADDR),
        .AP_AXIMM_59_ARLEN(AP_AXIMM_59_ARLEN),
        .AP_AXIMM_59_ARSIZE(AP_AXIMM_59_ARSIZE),
        .AP_AXIMM_59_ARBURST(AP_AXIMM_59_ARBURST),
        .AP_AXIMM_59_ARLOCK(AP_AXIMM_59_ARLOCK),
        .AP_AXIMM_59_ARCACHE(AP_AXIMM_59_ARCACHE),
        .AP_AXIMM_59_ARPROT(AP_AXIMM_59_ARPROT),
        .AP_AXIMM_59_ARREGION(AP_AXIMM_59_ARREGION),
        .AP_AXIMM_59_ARQOS(AP_AXIMM_59_ARQOS),
        .AP_AXIMM_59_ARVALID(AP_AXIMM_59_ARVALID),
        .AP_AXIMM_59_ARREADY(AP_AXIMM_59_ARREADY),
        .AP_AXIMM_59_RDATA(AP_AXIMM_59_RDATA),
        .AP_AXIMM_59_RRESP(AP_AXIMM_59_RRESP),
        .AP_AXIMM_59_RLAST(AP_AXIMM_59_RLAST),
        .AP_AXIMM_59_RVALID(AP_AXIMM_59_RVALID),
        .AP_AXIMM_59_RREADY(AP_AXIMM_59_RREADY),
        .M_AXIMM_59_AWADDR(M_AXIMM_59_AWADDR),
        .M_AXIMM_59_AWLEN(M_AXIMM_59_AWLEN),
        .M_AXIMM_59_AWSIZE(M_AXIMM_59_AWSIZE),
        .M_AXIMM_59_AWBURST(M_AXIMM_59_AWBURST),
        .M_AXIMM_59_AWLOCK(M_AXIMM_59_AWLOCK),
        .M_AXIMM_59_AWCACHE(M_AXIMM_59_AWCACHE),
        .M_AXIMM_59_AWPROT(M_AXIMM_59_AWPROT),
        .M_AXIMM_59_AWREGION(M_AXIMM_59_AWREGION),
        .M_AXIMM_59_AWQOS(M_AXIMM_59_AWQOS),
        .M_AXIMM_59_AWVALID(M_AXIMM_59_AWVALID),
        .M_AXIMM_59_AWREADY(M_AXIMM_59_AWREADY),
        .M_AXIMM_59_WDATA(M_AXIMM_59_WDATA),
        .M_AXIMM_59_WSTRB(M_AXIMM_59_WSTRB),
        .M_AXIMM_59_WLAST(M_AXIMM_59_WLAST),
        .M_AXIMM_59_WVALID(M_AXIMM_59_WVALID),
        .M_AXIMM_59_WREADY(M_AXIMM_59_WREADY),
        .M_AXIMM_59_BRESP(M_AXIMM_59_BRESP),
        .M_AXIMM_59_BVALID(M_AXIMM_59_BVALID),
        .M_AXIMM_59_BREADY(M_AXIMM_59_BREADY),
        .M_AXIMM_59_ARADDR(M_AXIMM_59_ARADDR),
        .M_AXIMM_59_ARLEN(M_AXIMM_59_ARLEN),
        .M_AXIMM_59_ARSIZE(M_AXIMM_59_ARSIZE),
        .M_AXIMM_59_ARBURST(M_AXIMM_59_ARBURST),
        .M_AXIMM_59_ARLOCK(M_AXIMM_59_ARLOCK),
        .M_AXIMM_59_ARCACHE(M_AXIMM_59_ARCACHE),
        .M_AXIMM_59_ARPROT(M_AXIMM_59_ARPROT),
        .M_AXIMM_59_ARREGION(M_AXIMM_59_ARREGION),
        .M_AXIMM_59_ARQOS(M_AXIMM_59_ARQOS),
        .M_AXIMM_59_ARVALID(M_AXIMM_59_ARVALID),
        .M_AXIMM_59_ARREADY(M_AXIMM_59_ARREADY),
        .M_AXIMM_59_RDATA(M_AXIMM_59_RDATA),
        .M_AXIMM_59_RRESP(M_AXIMM_59_RRESP),
        .M_AXIMM_59_RLAST(M_AXIMM_59_RLAST),
        .M_AXIMM_59_RVALID(M_AXIMM_59_RVALID),
        .M_AXIMM_59_RREADY(M_AXIMM_59_RREADY),
        .AP_AXIMM_60_AWADDR(AP_AXIMM_60_AWADDR),
        .AP_AXIMM_60_AWLEN(AP_AXIMM_60_AWLEN),
        .AP_AXIMM_60_AWSIZE(AP_AXIMM_60_AWSIZE),
        .AP_AXIMM_60_AWBURST(AP_AXIMM_60_AWBURST),
        .AP_AXIMM_60_AWLOCK(AP_AXIMM_60_AWLOCK),
        .AP_AXIMM_60_AWCACHE(AP_AXIMM_60_AWCACHE),
        .AP_AXIMM_60_AWPROT(AP_AXIMM_60_AWPROT),
        .AP_AXIMM_60_AWREGION(AP_AXIMM_60_AWREGION),
        .AP_AXIMM_60_AWQOS(AP_AXIMM_60_AWQOS),
        .AP_AXIMM_60_AWVALID(AP_AXIMM_60_AWVALID),
        .AP_AXIMM_60_AWREADY(AP_AXIMM_60_AWREADY),
        .AP_AXIMM_60_WDATA(AP_AXIMM_60_WDATA),
        .AP_AXIMM_60_WSTRB(AP_AXIMM_60_WSTRB),
        .AP_AXIMM_60_WLAST(AP_AXIMM_60_WLAST),
        .AP_AXIMM_60_WVALID(AP_AXIMM_60_WVALID),
        .AP_AXIMM_60_WREADY(AP_AXIMM_60_WREADY),
        .AP_AXIMM_60_BRESP(AP_AXIMM_60_BRESP),
        .AP_AXIMM_60_BVALID(AP_AXIMM_60_BVALID),
        .AP_AXIMM_60_BREADY(AP_AXIMM_60_BREADY),
        .AP_AXIMM_60_ARADDR(AP_AXIMM_60_ARADDR),
        .AP_AXIMM_60_ARLEN(AP_AXIMM_60_ARLEN),
        .AP_AXIMM_60_ARSIZE(AP_AXIMM_60_ARSIZE),
        .AP_AXIMM_60_ARBURST(AP_AXIMM_60_ARBURST),
        .AP_AXIMM_60_ARLOCK(AP_AXIMM_60_ARLOCK),
        .AP_AXIMM_60_ARCACHE(AP_AXIMM_60_ARCACHE),
        .AP_AXIMM_60_ARPROT(AP_AXIMM_60_ARPROT),
        .AP_AXIMM_60_ARREGION(AP_AXIMM_60_ARREGION),
        .AP_AXIMM_60_ARQOS(AP_AXIMM_60_ARQOS),
        .AP_AXIMM_60_ARVALID(AP_AXIMM_60_ARVALID),
        .AP_AXIMM_60_ARREADY(AP_AXIMM_60_ARREADY),
        .AP_AXIMM_60_RDATA(AP_AXIMM_60_RDATA),
        .AP_AXIMM_60_RRESP(AP_AXIMM_60_RRESP),
        .AP_AXIMM_60_RLAST(AP_AXIMM_60_RLAST),
        .AP_AXIMM_60_RVALID(AP_AXIMM_60_RVALID),
        .AP_AXIMM_60_RREADY(AP_AXIMM_60_RREADY),
        .M_AXIMM_60_AWADDR(M_AXIMM_60_AWADDR),
        .M_AXIMM_60_AWLEN(M_AXIMM_60_AWLEN),
        .M_AXIMM_60_AWSIZE(M_AXIMM_60_AWSIZE),
        .M_AXIMM_60_AWBURST(M_AXIMM_60_AWBURST),
        .M_AXIMM_60_AWLOCK(M_AXIMM_60_AWLOCK),
        .M_AXIMM_60_AWCACHE(M_AXIMM_60_AWCACHE),
        .M_AXIMM_60_AWPROT(M_AXIMM_60_AWPROT),
        .M_AXIMM_60_AWREGION(M_AXIMM_60_AWREGION),
        .M_AXIMM_60_AWQOS(M_AXIMM_60_AWQOS),
        .M_AXIMM_60_AWVALID(M_AXIMM_60_AWVALID),
        .M_AXIMM_60_AWREADY(M_AXIMM_60_AWREADY),
        .M_AXIMM_60_WDATA(M_AXIMM_60_WDATA),
        .M_AXIMM_60_WSTRB(M_AXIMM_60_WSTRB),
        .M_AXIMM_60_WLAST(M_AXIMM_60_WLAST),
        .M_AXIMM_60_WVALID(M_AXIMM_60_WVALID),
        .M_AXIMM_60_WREADY(M_AXIMM_60_WREADY),
        .M_AXIMM_60_BRESP(M_AXIMM_60_BRESP),
        .M_AXIMM_60_BVALID(M_AXIMM_60_BVALID),
        .M_AXIMM_60_BREADY(M_AXIMM_60_BREADY),
        .M_AXIMM_60_ARADDR(M_AXIMM_60_ARADDR),
        .M_AXIMM_60_ARLEN(M_AXIMM_60_ARLEN),
        .M_AXIMM_60_ARSIZE(M_AXIMM_60_ARSIZE),
        .M_AXIMM_60_ARBURST(M_AXIMM_60_ARBURST),
        .M_AXIMM_60_ARLOCK(M_AXIMM_60_ARLOCK),
        .M_AXIMM_60_ARCACHE(M_AXIMM_60_ARCACHE),
        .M_AXIMM_60_ARPROT(M_AXIMM_60_ARPROT),
        .M_AXIMM_60_ARREGION(M_AXIMM_60_ARREGION),
        .M_AXIMM_60_ARQOS(M_AXIMM_60_ARQOS),
        .M_AXIMM_60_ARVALID(M_AXIMM_60_ARVALID),
        .M_AXIMM_60_ARREADY(M_AXIMM_60_ARREADY),
        .M_AXIMM_60_RDATA(M_AXIMM_60_RDATA),
        .M_AXIMM_60_RRESP(M_AXIMM_60_RRESP),
        .M_AXIMM_60_RLAST(M_AXIMM_60_RLAST),
        .M_AXIMM_60_RVALID(M_AXIMM_60_RVALID),
        .M_AXIMM_60_RREADY(M_AXIMM_60_RREADY),
        .AP_AXIMM_61_AWADDR(AP_AXIMM_61_AWADDR),
        .AP_AXIMM_61_AWLEN(AP_AXIMM_61_AWLEN),
        .AP_AXIMM_61_AWSIZE(AP_AXIMM_61_AWSIZE),
        .AP_AXIMM_61_AWBURST(AP_AXIMM_61_AWBURST),
        .AP_AXIMM_61_AWLOCK(AP_AXIMM_61_AWLOCK),
        .AP_AXIMM_61_AWCACHE(AP_AXIMM_61_AWCACHE),
        .AP_AXIMM_61_AWPROT(AP_AXIMM_61_AWPROT),
        .AP_AXIMM_61_AWREGION(AP_AXIMM_61_AWREGION),
        .AP_AXIMM_61_AWQOS(AP_AXIMM_61_AWQOS),
        .AP_AXIMM_61_AWVALID(AP_AXIMM_61_AWVALID),
        .AP_AXIMM_61_AWREADY(AP_AXIMM_61_AWREADY),
        .AP_AXIMM_61_WDATA(AP_AXIMM_61_WDATA),
        .AP_AXIMM_61_WSTRB(AP_AXIMM_61_WSTRB),
        .AP_AXIMM_61_WLAST(AP_AXIMM_61_WLAST),
        .AP_AXIMM_61_WVALID(AP_AXIMM_61_WVALID),
        .AP_AXIMM_61_WREADY(AP_AXIMM_61_WREADY),
        .AP_AXIMM_61_BRESP(AP_AXIMM_61_BRESP),
        .AP_AXIMM_61_BVALID(AP_AXIMM_61_BVALID),
        .AP_AXIMM_61_BREADY(AP_AXIMM_61_BREADY),
        .AP_AXIMM_61_ARADDR(AP_AXIMM_61_ARADDR),
        .AP_AXIMM_61_ARLEN(AP_AXIMM_61_ARLEN),
        .AP_AXIMM_61_ARSIZE(AP_AXIMM_61_ARSIZE),
        .AP_AXIMM_61_ARBURST(AP_AXIMM_61_ARBURST),
        .AP_AXIMM_61_ARLOCK(AP_AXIMM_61_ARLOCK),
        .AP_AXIMM_61_ARCACHE(AP_AXIMM_61_ARCACHE),
        .AP_AXIMM_61_ARPROT(AP_AXIMM_61_ARPROT),
        .AP_AXIMM_61_ARREGION(AP_AXIMM_61_ARREGION),
        .AP_AXIMM_61_ARQOS(AP_AXIMM_61_ARQOS),
        .AP_AXIMM_61_ARVALID(AP_AXIMM_61_ARVALID),
        .AP_AXIMM_61_ARREADY(AP_AXIMM_61_ARREADY),
        .AP_AXIMM_61_RDATA(AP_AXIMM_61_RDATA),
        .AP_AXIMM_61_RRESP(AP_AXIMM_61_RRESP),
        .AP_AXIMM_61_RLAST(AP_AXIMM_61_RLAST),
        .AP_AXIMM_61_RVALID(AP_AXIMM_61_RVALID),
        .AP_AXIMM_61_RREADY(AP_AXIMM_61_RREADY),
        .M_AXIMM_61_AWADDR(M_AXIMM_61_AWADDR),
        .M_AXIMM_61_AWLEN(M_AXIMM_61_AWLEN),
        .M_AXIMM_61_AWSIZE(M_AXIMM_61_AWSIZE),
        .M_AXIMM_61_AWBURST(M_AXIMM_61_AWBURST),
        .M_AXIMM_61_AWLOCK(M_AXIMM_61_AWLOCK),
        .M_AXIMM_61_AWCACHE(M_AXIMM_61_AWCACHE),
        .M_AXIMM_61_AWPROT(M_AXIMM_61_AWPROT),
        .M_AXIMM_61_AWREGION(M_AXIMM_61_AWREGION),
        .M_AXIMM_61_AWQOS(M_AXIMM_61_AWQOS),
        .M_AXIMM_61_AWVALID(M_AXIMM_61_AWVALID),
        .M_AXIMM_61_AWREADY(M_AXIMM_61_AWREADY),
        .M_AXIMM_61_WDATA(M_AXIMM_61_WDATA),
        .M_AXIMM_61_WSTRB(M_AXIMM_61_WSTRB),
        .M_AXIMM_61_WLAST(M_AXIMM_61_WLAST),
        .M_AXIMM_61_WVALID(M_AXIMM_61_WVALID),
        .M_AXIMM_61_WREADY(M_AXIMM_61_WREADY),
        .M_AXIMM_61_BRESP(M_AXIMM_61_BRESP),
        .M_AXIMM_61_BVALID(M_AXIMM_61_BVALID),
        .M_AXIMM_61_BREADY(M_AXIMM_61_BREADY),
        .M_AXIMM_61_ARADDR(M_AXIMM_61_ARADDR),
        .M_AXIMM_61_ARLEN(M_AXIMM_61_ARLEN),
        .M_AXIMM_61_ARSIZE(M_AXIMM_61_ARSIZE),
        .M_AXIMM_61_ARBURST(M_AXIMM_61_ARBURST),
        .M_AXIMM_61_ARLOCK(M_AXIMM_61_ARLOCK),
        .M_AXIMM_61_ARCACHE(M_AXIMM_61_ARCACHE),
        .M_AXIMM_61_ARPROT(M_AXIMM_61_ARPROT),
        .M_AXIMM_61_ARREGION(M_AXIMM_61_ARREGION),
        .M_AXIMM_61_ARQOS(M_AXIMM_61_ARQOS),
        .M_AXIMM_61_ARVALID(M_AXIMM_61_ARVALID),
        .M_AXIMM_61_ARREADY(M_AXIMM_61_ARREADY),
        .M_AXIMM_61_RDATA(M_AXIMM_61_RDATA),
        .M_AXIMM_61_RRESP(M_AXIMM_61_RRESP),
        .M_AXIMM_61_RLAST(M_AXIMM_61_RLAST),
        .M_AXIMM_61_RVALID(M_AXIMM_61_RVALID),
        .M_AXIMM_61_RREADY(M_AXIMM_61_RREADY),
        .AP_AXIMM_62_AWADDR(AP_AXIMM_62_AWADDR),
        .AP_AXIMM_62_AWLEN(AP_AXIMM_62_AWLEN),
        .AP_AXIMM_62_AWSIZE(AP_AXIMM_62_AWSIZE),
        .AP_AXIMM_62_AWBURST(AP_AXIMM_62_AWBURST),
        .AP_AXIMM_62_AWLOCK(AP_AXIMM_62_AWLOCK),
        .AP_AXIMM_62_AWCACHE(AP_AXIMM_62_AWCACHE),
        .AP_AXIMM_62_AWPROT(AP_AXIMM_62_AWPROT),
        .AP_AXIMM_62_AWREGION(AP_AXIMM_62_AWREGION),
        .AP_AXIMM_62_AWQOS(AP_AXIMM_62_AWQOS),
        .AP_AXIMM_62_AWVALID(AP_AXIMM_62_AWVALID),
        .AP_AXIMM_62_AWREADY(AP_AXIMM_62_AWREADY),
        .AP_AXIMM_62_WDATA(AP_AXIMM_62_WDATA),
        .AP_AXIMM_62_WSTRB(AP_AXIMM_62_WSTRB),
        .AP_AXIMM_62_WLAST(AP_AXIMM_62_WLAST),
        .AP_AXIMM_62_WVALID(AP_AXIMM_62_WVALID),
        .AP_AXIMM_62_WREADY(AP_AXIMM_62_WREADY),
        .AP_AXIMM_62_BRESP(AP_AXIMM_62_BRESP),
        .AP_AXIMM_62_BVALID(AP_AXIMM_62_BVALID),
        .AP_AXIMM_62_BREADY(AP_AXIMM_62_BREADY),
        .AP_AXIMM_62_ARADDR(AP_AXIMM_62_ARADDR),
        .AP_AXIMM_62_ARLEN(AP_AXIMM_62_ARLEN),
        .AP_AXIMM_62_ARSIZE(AP_AXIMM_62_ARSIZE),
        .AP_AXIMM_62_ARBURST(AP_AXIMM_62_ARBURST),
        .AP_AXIMM_62_ARLOCK(AP_AXIMM_62_ARLOCK),
        .AP_AXIMM_62_ARCACHE(AP_AXIMM_62_ARCACHE),
        .AP_AXIMM_62_ARPROT(AP_AXIMM_62_ARPROT),
        .AP_AXIMM_62_ARREGION(AP_AXIMM_62_ARREGION),
        .AP_AXIMM_62_ARQOS(AP_AXIMM_62_ARQOS),
        .AP_AXIMM_62_ARVALID(AP_AXIMM_62_ARVALID),
        .AP_AXIMM_62_ARREADY(AP_AXIMM_62_ARREADY),
        .AP_AXIMM_62_RDATA(AP_AXIMM_62_RDATA),
        .AP_AXIMM_62_RRESP(AP_AXIMM_62_RRESP),
        .AP_AXIMM_62_RLAST(AP_AXIMM_62_RLAST),
        .AP_AXIMM_62_RVALID(AP_AXIMM_62_RVALID),
        .AP_AXIMM_62_RREADY(AP_AXIMM_62_RREADY),
        .M_AXIMM_62_AWADDR(M_AXIMM_62_AWADDR),
        .M_AXIMM_62_AWLEN(M_AXIMM_62_AWLEN),
        .M_AXIMM_62_AWSIZE(M_AXIMM_62_AWSIZE),
        .M_AXIMM_62_AWBURST(M_AXIMM_62_AWBURST),
        .M_AXIMM_62_AWLOCK(M_AXIMM_62_AWLOCK),
        .M_AXIMM_62_AWCACHE(M_AXIMM_62_AWCACHE),
        .M_AXIMM_62_AWPROT(M_AXIMM_62_AWPROT),
        .M_AXIMM_62_AWREGION(M_AXIMM_62_AWREGION),
        .M_AXIMM_62_AWQOS(M_AXIMM_62_AWQOS),
        .M_AXIMM_62_AWVALID(M_AXIMM_62_AWVALID),
        .M_AXIMM_62_AWREADY(M_AXIMM_62_AWREADY),
        .M_AXIMM_62_WDATA(M_AXIMM_62_WDATA),
        .M_AXIMM_62_WSTRB(M_AXIMM_62_WSTRB),
        .M_AXIMM_62_WLAST(M_AXIMM_62_WLAST),
        .M_AXIMM_62_WVALID(M_AXIMM_62_WVALID),
        .M_AXIMM_62_WREADY(M_AXIMM_62_WREADY),
        .M_AXIMM_62_BRESP(M_AXIMM_62_BRESP),
        .M_AXIMM_62_BVALID(M_AXIMM_62_BVALID),
        .M_AXIMM_62_BREADY(M_AXIMM_62_BREADY),
        .M_AXIMM_62_ARADDR(M_AXIMM_62_ARADDR),
        .M_AXIMM_62_ARLEN(M_AXIMM_62_ARLEN),
        .M_AXIMM_62_ARSIZE(M_AXIMM_62_ARSIZE),
        .M_AXIMM_62_ARBURST(M_AXIMM_62_ARBURST),
        .M_AXIMM_62_ARLOCK(M_AXIMM_62_ARLOCK),
        .M_AXIMM_62_ARCACHE(M_AXIMM_62_ARCACHE),
        .M_AXIMM_62_ARPROT(M_AXIMM_62_ARPROT),
        .M_AXIMM_62_ARREGION(M_AXIMM_62_ARREGION),
        .M_AXIMM_62_ARQOS(M_AXIMM_62_ARQOS),
        .M_AXIMM_62_ARVALID(M_AXIMM_62_ARVALID),
        .M_AXIMM_62_ARREADY(M_AXIMM_62_ARREADY),
        .M_AXIMM_62_RDATA(M_AXIMM_62_RDATA),
        .M_AXIMM_62_RRESP(M_AXIMM_62_RRESP),
        .M_AXIMM_62_RLAST(M_AXIMM_62_RLAST),
        .M_AXIMM_62_RVALID(M_AXIMM_62_RVALID),
        .M_AXIMM_62_RREADY(M_AXIMM_62_RREADY),
        .AP_AXIMM_63_AWADDR(AP_AXIMM_63_AWADDR),
        .AP_AXIMM_63_AWLEN(AP_AXIMM_63_AWLEN),
        .AP_AXIMM_63_AWSIZE(AP_AXIMM_63_AWSIZE),
        .AP_AXIMM_63_AWBURST(AP_AXIMM_63_AWBURST),
        .AP_AXIMM_63_AWLOCK(AP_AXIMM_63_AWLOCK),
        .AP_AXIMM_63_AWCACHE(AP_AXIMM_63_AWCACHE),
        .AP_AXIMM_63_AWPROT(AP_AXIMM_63_AWPROT),
        .AP_AXIMM_63_AWREGION(AP_AXIMM_63_AWREGION),
        .AP_AXIMM_63_AWQOS(AP_AXIMM_63_AWQOS),
        .AP_AXIMM_63_AWVALID(AP_AXIMM_63_AWVALID),
        .AP_AXIMM_63_AWREADY(AP_AXIMM_63_AWREADY),
        .AP_AXIMM_63_WDATA(AP_AXIMM_63_WDATA),
        .AP_AXIMM_63_WSTRB(AP_AXIMM_63_WSTRB),
        .AP_AXIMM_63_WLAST(AP_AXIMM_63_WLAST),
        .AP_AXIMM_63_WVALID(AP_AXIMM_63_WVALID),
        .AP_AXIMM_63_WREADY(AP_AXIMM_63_WREADY),
        .AP_AXIMM_63_BRESP(AP_AXIMM_63_BRESP),
        .AP_AXIMM_63_BVALID(AP_AXIMM_63_BVALID),
        .AP_AXIMM_63_BREADY(AP_AXIMM_63_BREADY),
        .AP_AXIMM_63_ARADDR(AP_AXIMM_63_ARADDR),
        .AP_AXIMM_63_ARLEN(AP_AXIMM_63_ARLEN),
        .AP_AXIMM_63_ARSIZE(AP_AXIMM_63_ARSIZE),
        .AP_AXIMM_63_ARBURST(AP_AXIMM_63_ARBURST),
        .AP_AXIMM_63_ARLOCK(AP_AXIMM_63_ARLOCK),
        .AP_AXIMM_63_ARCACHE(AP_AXIMM_63_ARCACHE),
        .AP_AXIMM_63_ARPROT(AP_AXIMM_63_ARPROT),
        .AP_AXIMM_63_ARREGION(AP_AXIMM_63_ARREGION),
        .AP_AXIMM_63_ARQOS(AP_AXIMM_63_ARQOS),
        .AP_AXIMM_63_ARVALID(AP_AXIMM_63_ARVALID),
        .AP_AXIMM_63_ARREADY(AP_AXIMM_63_ARREADY),
        .AP_AXIMM_63_RDATA(AP_AXIMM_63_RDATA),
        .AP_AXIMM_63_RRESP(AP_AXIMM_63_RRESP),
        .AP_AXIMM_63_RLAST(AP_AXIMM_63_RLAST),
        .AP_AXIMM_63_RVALID(AP_AXIMM_63_RVALID),
        .AP_AXIMM_63_RREADY(AP_AXIMM_63_RREADY),
        .M_AXIMM_63_AWADDR(M_AXIMM_63_AWADDR),
        .M_AXIMM_63_AWLEN(M_AXIMM_63_AWLEN),
        .M_AXIMM_63_AWSIZE(M_AXIMM_63_AWSIZE),
        .M_AXIMM_63_AWBURST(M_AXIMM_63_AWBURST),
        .M_AXIMM_63_AWLOCK(M_AXIMM_63_AWLOCK),
        .M_AXIMM_63_AWCACHE(M_AXIMM_63_AWCACHE),
        .M_AXIMM_63_AWPROT(M_AXIMM_63_AWPROT),
        .M_AXIMM_63_AWREGION(M_AXIMM_63_AWREGION),
        .M_AXIMM_63_AWQOS(M_AXIMM_63_AWQOS),
        .M_AXIMM_63_AWVALID(M_AXIMM_63_AWVALID),
        .M_AXIMM_63_AWREADY(M_AXIMM_63_AWREADY),
        .M_AXIMM_63_WDATA(M_AXIMM_63_WDATA),
        .M_AXIMM_63_WSTRB(M_AXIMM_63_WSTRB),
        .M_AXIMM_63_WLAST(M_AXIMM_63_WLAST),
        .M_AXIMM_63_WVALID(M_AXIMM_63_WVALID),
        .M_AXIMM_63_WREADY(M_AXIMM_63_WREADY),
        .M_AXIMM_63_BRESP(M_AXIMM_63_BRESP),
        .M_AXIMM_63_BVALID(M_AXIMM_63_BVALID),
        .M_AXIMM_63_BREADY(M_AXIMM_63_BREADY),
        .M_AXIMM_63_ARADDR(M_AXIMM_63_ARADDR),
        .M_AXIMM_63_ARLEN(M_AXIMM_63_ARLEN),
        .M_AXIMM_63_ARSIZE(M_AXIMM_63_ARSIZE),
        .M_AXIMM_63_ARBURST(M_AXIMM_63_ARBURST),
        .M_AXIMM_63_ARLOCK(M_AXIMM_63_ARLOCK),
        .M_AXIMM_63_ARCACHE(M_AXIMM_63_ARCACHE),
        .M_AXIMM_63_ARPROT(M_AXIMM_63_ARPROT),
        .M_AXIMM_63_ARREGION(M_AXIMM_63_ARREGION),
        .M_AXIMM_63_ARQOS(M_AXIMM_63_ARQOS),
        .M_AXIMM_63_ARVALID(M_AXIMM_63_ARVALID),
        .M_AXIMM_63_ARREADY(M_AXIMM_63_ARREADY),
        .M_AXIMM_63_RDATA(M_AXIMM_63_RDATA),
        .M_AXIMM_63_RRESP(M_AXIMM_63_RRESP),
        .M_AXIMM_63_RLAST(M_AXIMM_63_RLAST),
        .M_AXIMM_63_RVALID(M_AXIMM_63_RVALID),
        .M_AXIMM_63_RREADY(M_AXIMM_63_RREADY),
        .AP_AXIMM_64_AWADDR(AP_AXIMM_64_AWADDR),
        .AP_AXIMM_64_AWLEN(AP_AXIMM_64_AWLEN),
        .AP_AXIMM_64_AWSIZE(AP_AXIMM_64_AWSIZE),
        .AP_AXIMM_64_AWBURST(AP_AXIMM_64_AWBURST),
        .AP_AXIMM_64_AWLOCK(AP_AXIMM_64_AWLOCK),
        .AP_AXIMM_64_AWCACHE(AP_AXIMM_64_AWCACHE),
        .AP_AXIMM_64_AWPROT(AP_AXIMM_64_AWPROT),
        .AP_AXIMM_64_AWREGION(AP_AXIMM_64_AWREGION),
        .AP_AXIMM_64_AWQOS(AP_AXIMM_64_AWQOS),
        .AP_AXIMM_64_AWVALID(AP_AXIMM_64_AWVALID),
        .AP_AXIMM_64_AWREADY(AP_AXIMM_64_AWREADY),
        .AP_AXIMM_64_WDATA(AP_AXIMM_64_WDATA),
        .AP_AXIMM_64_WSTRB(AP_AXIMM_64_WSTRB),
        .AP_AXIMM_64_WLAST(AP_AXIMM_64_WLAST),
        .AP_AXIMM_64_WVALID(AP_AXIMM_64_WVALID),
        .AP_AXIMM_64_WREADY(AP_AXIMM_64_WREADY),
        .AP_AXIMM_64_BRESP(AP_AXIMM_64_BRESP),
        .AP_AXIMM_64_BVALID(AP_AXIMM_64_BVALID),
        .AP_AXIMM_64_BREADY(AP_AXIMM_64_BREADY),
        .AP_AXIMM_64_ARADDR(AP_AXIMM_64_ARADDR),
        .AP_AXIMM_64_ARLEN(AP_AXIMM_64_ARLEN),
        .AP_AXIMM_64_ARSIZE(AP_AXIMM_64_ARSIZE),
        .AP_AXIMM_64_ARBURST(AP_AXIMM_64_ARBURST),
        .AP_AXIMM_64_ARLOCK(AP_AXIMM_64_ARLOCK),
        .AP_AXIMM_64_ARCACHE(AP_AXIMM_64_ARCACHE),
        .AP_AXIMM_64_ARPROT(AP_AXIMM_64_ARPROT),
        .AP_AXIMM_64_ARREGION(AP_AXIMM_64_ARREGION),
        .AP_AXIMM_64_ARQOS(AP_AXIMM_64_ARQOS),
        .AP_AXIMM_64_ARVALID(AP_AXIMM_64_ARVALID),
        .AP_AXIMM_64_ARREADY(AP_AXIMM_64_ARREADY),
        .AP_AXIMM_64_RDATA(AP_AXIMM_64_RDATA),
        .AP_AXIMM_64_RRESP(AP_AXIMM_64_RRESP),
        .AP_AXIMM_64_RLAST(AP_AXIMM_64_RLAST),
        .AP_AXIMM_64_RVALID(AP_AXIMM_64_RVALID),
        .AP_AXIMM_64_RREADY(AP_AXIMM_64_RREADY),
        .M_AXIMM_64_AWADDR(M_AXIMM_64_AWADDR),
        .M_AXIMM_64_AWLEN(M_AXIMM_64_AWLEN),
        .M_AXIMM_64_AWSIZE(M_AXIMM_64_AWSIZE),
        .M_AXIMM_64_AWBURST(M_AXIMM_64_AWBURST),
        .M_AXIMM_64_AWLOCK(M_AXIMM_64_AWLOCK),
        .M_AXIMM_64_AWCACHE(M_AXIMM_64_AWCACHE),
        .M_AXIMM_64_AWPROT(M_AXIMM_64_AWPROT),
        .M_AXIMM_64_AWREGION(M_AXIMM_64_AWREGION),
        .M_AXIMM_64_AWQOS(M_AXIMM_64_AWQOS),
        .M_AXIMM_64_AWVALID(M_AXIMM_64_AWVALID),
        .M_AXIMM_64_AWREADY(M_AXIMM_64_AWREADY),
        .M_AXIMM_64_WDATA(M_AXIMM_64_WDATA),
        .M_AXIMM_64_WSTRB(M_AXIMM_64_WSTRB),
        .M_AXIMM_64_WLAST(M_AXIMM_64_WLAST),
        .M_AXIMM_64_WVALID(M_AXIMM_64_WVALID),
        .M_AXIMM_64_WREADY(M_AXIMM_64_WREADY),
        .M_AXIMM_64_BRESP(M_AXIMM_64_BRESP),
        .M_AXIMM_64_BVALID(M_AXIMM_64_BVALID),
        .M_AXIMM_64_BREADY(M_AXIMM_64_BREADY),
        .M_AXIMM_64_ARADDR(M_AXIMM_64_ARADDR),
        .M_AXIMM_64_ARLEN(M_AXIMM_64_ARLEN),
        .M_AXIMM_64_ARSIZE(M_AXIMM_64_ARSIZE),
        .M_AXIMM_64_ARBURST(M_AXIMM_64_ARBURST),
        .M_AXIMM_64_ARLOCK(M_AXIMM_64_ARLOCK),
        .M_AXIMM_64_ARCACHE(M_AXIMM_64_ARCACHE),
        .M_AXIMM_64_ARPROT(M_AXIMM_64_ARPROT),
        .M_AXIMM_64_ARREGION(M_AXIMM_64_ARREGION),
        .M_AXIMM_64_ARQOS(M_AXIMM_64_ARQOS),
        .M_AXIMM_64_ARVALID(M_AXIMM_64_ARVALID),
        .M_AXIMM_64_ARREADY(M_AXIMM_64_ARREADY),
        .M_AXIMM_64_RDATA(M_AXIMM_64_RDATA),
        .M_AXIMM_64_RRESP(M_AXIMM_64_RRESP),
        .M_AXIMM_64_RLAST(M_AXIMM_64_RLAST),
        .M_AXIMM_64_RVALID(M_AXIMM_64_RVALID),
        .M_AXIMM_64_RREADY(M_AXIMM_64_RREADY),
        .AP_AXIMM_65_AWADDR(AP_AXIMM_65_AWADDR),
        .AP_AXIMM_65_AWLEN(AP_AXIMM_65_AWLEN),
        .AP_AXIMM_65_AWSIZE(AP_AXIMM_65_AWSIZE),
        .AP_AXIMM_65_AWBURST(AP_AXIMM_65_AWBURST),
        .AP_AXIMM_65_AWLOCK(AP_AXIMM_65_AWLOCK),
        .AP_AXIMM_65_AWCACHE(AP_AXIMM_65_AWCACHE),
        .AP_AXIMM_65_AWPROT(AP_AXIMM_65_AWPROT),
        .AP_AXIMM_65_AWREGION(AP_AXIMM_65_AWREGION),
        .AP_AXIMM_65_AWQOS(AP_AXIMM_65_AWQOS),
        .AP_AXIMM_65_AWVALID(AP_AXIMM_65_AWVALID),
        .AP_AXIMM_65_AWREADY(AP_AXIMM_65_AWREADY),
        .AP_AXIMM_65_WDATA(AP_AXIMM_65_WDATA),
        .AP_AXIMM_65_WSTRB(AP_AXIMM_65_WSTRB),
        .AP_AXIMM_65_WLAST(AP_AXIMM_65_WLAST),
        .AP_AXIMM_65_WVALID(AP_AXIMM_65_WVALID),
        .AP_AXIMM_65_WREADY(AP_AXIMM_65_WREADY),
        .AP_AXIMM_65_BRESP(AP_AXIMM_65_BRESP),
        .AP_AXIMM_65_BVALID(AP_AXIMM_65_BVALID),
        .AP_AXIMM_65_BREADY(AP_AXIMM_65_BREADY),
        .AP_AXIMM_65_ARADDR(AP_AXIMM_65_ARADDR),
        .AP_AXIMM_65_ARLEN(AP_AXIMM_65_ARLEN),
        .AP_AXIMM_65_ARSIZE(AP_AXIMM_65_ARSIZE),
        .AP_AXIMM_65_ARBURST(AP_AXIMM_65_ARBURST),
        .AP_AXIMM_65_ARLOCK(AP_AXIMM_65_ARLOCK),
        .AP_AXIMM_65_ARCACHE(AP_AXIMM_65_ARCACHE),
        .AP_AXIMM_65_ARPROT(AP_AXIMM_65_ARPROT),
        .AP_AXIMM_65_ARREGION(AP_AXIMM_65_ARREGION),
        .AP_AXIMM_65_ARQOS(AP_AXIMM_65_ARQOS),
        .AP_AXIMM_65_ARVALID(AP_AXIMM_65_ARVALID),
        .AP_AXIMM_65_ARREADY(AP_AXIMM_65_ARREADY),
        .AP_AXIMM_65_RDATA(AP_AXIMM_65_RDATA),
        .AP_AXIMM_65_RRESP(AP_AXIMM_65_RRESP),
        .AP_AXIMM_65_RLAST(AP_AXIMM_65_RLAST),
        .AP_AXIMM_65_RVALID(AP_AXIMM_65_RVALID),
        .AP_AXIMM_65_RREADY(AP_AXIMM_65_RREADY),
        .M_AXIMM_65_AWADDR(M_AXIMM_65_AWADDR),
        .M_AXIMM_65_AWLEN(M_AXIMM_65_AWLEN),
        .M_AXIMM_65_AWSIZE(M_AXIMM_65_AWSIZE),
        .M_AXIMM_65_AWBURST(M_AXIMM_65_AWBURST),
        .M_AXIMM_65_AWLOCK(M_AXIMM_65_AWLOCK),
        .M_AXIMM_65_AWCACHE(M_AXIMM_65_AWCACHE),
        .M_AXIMM_65_AWPROT(M_AXIMM_65_AWPROT),
        .M_AXIMM_65_AWREGION(M_AXIMM_65_AWREGION),
        .M_AXIMM_65_AWQOS(M_AXIMM_65_AWQOS),
        .M_AXIMM_65_AWVALID(M_AXIMM_65_AWVALID),
        .M_AXIMM_65_AWREADY(M_AXIMM_65_AWREADY),
        .M_AXIMM_65_WDATA(M_AXIMM_65_WDATA),
        .M_AXIMM_65_WSTRB(M_AXIMM_65_WSTRB),
        .M_AXIMM_65_WLAST(M_AXIMM_65_WLAST),
        .M_AXIMM_65_WVALID(M_AXIMM_65_WVALID),
        .M_AXIMM_65_WREADY(M_AXIMM_65_WREADY),
        .M_AXIMM_65_BRESP(M_AXIMM_65_BRESP),
        .M_AXIMM_65_BVALID(M_AXIMM_65_BVALID),
        .M_AXIMM_65_BREADY(M_AXIMM_65_BREADY),
        .M_AXIMM_65_ARADDR(M_AXIMM_65_ARADDR),
        .M_AXIMM_65_ARLEN(M_AXIMM_65_ARLEN),
        .M_AXIMM_65_ARSIZE(M_AXIMM_65_ARSIZE),
        .M_AXIMM_65_ARBURST(M_AXIMM_65_ARBURST),
        .M_AXIMM_65_ARLOCK(M_AXIMM_65_ARLOCK),
        .M_AXIMM_65_ARCACHE(M_AXIMM_65_ARCACHE),
        .M_AXIMM_65_ARPROT(M_AXIMM_65_ARPROT),
        .M_AXIMM_65_ARREGION(M_AXIMM_65_ARREGION),
        .M_AXIMM_65_ARQOS(M_AXIMM_65_ARQOS),
        .M_AXIMM_65_ARVALID(M_AXIMM_65_ARVALID),
        .M_AXIMM_65_ARREADY(M_AXIMM_65_ARREADY),
        .M_AXIMM_65_RDATA(M_AXIMM_65_RDATA),
        .M_AXIMM_65_RRESP(M_AXIMM_65_RRESP),
        .M_AXIMM_65_RLAST(M_AXIMM_65_RLAST),
        .M_AXIMM_65_RVALID(M_AXIMM_65_RVALID),
        .M_AXIMM_65_RREADY(M_AXIMM_65_RREADY),
        .AP_AXIMM_66_AWADDR(AP_AXIMM_66_AWADDR),
        .AP_AXIMM_66_AWLEN(AP_AXIMM_66_AWLEN),
        .AP_AXIMM_66_AWSIZE(AP_AXIMM_66_AWSIZE),
        .AP_AXIMM_66_AWBURST(AP_AXIMM_66_AWBURST),
        .AP_AXIMM_66_AWLOCK(AP_AXIMM_66_AWLOCK),
        .AP_AXIMM_66_AWCACHE(AP_AXIMM_66_AWCACHE),
        .AP_AXIMM_66_AWPROT(AP_AXIMM_66_AWPROT),
        .AP_AXIMM_66_AWREGION(AP_AXIMM_66_AWREGION),
        .AP_AXIMM_66_AWQOS(AP_AXIMM_66_AWQOS),
        .AP_AXIMM_66_AWVALID(AP_AXIMM_66_AWVALID),
        .AP_AXIMM_66_AWREADY(AP_AXIMM_66_AWREADY),
        .AP_AXIMM_66_WDATA(AP_AXIMM_66_WDATA),
        .AP_AXIMM_66_WSTRB(AP_AXIMM_66_WSTRB),
        .AP_AXIMM_66_WLAST(AP_AXIMM_66_WLAST),
        .AP_AXIMM_66_WVALID(AP_AXIMM_66_WVALID),
        .AP_AXIMM_66_WREADY(AP_AXIMM_66_WREADY),
        .AP_AXIMM_66_BRESP(AP_AXIMM_66_BRESP),
        .AP_AXIMM_66_BVALID(AP_AXIMM_66_BVALID),
        .AP_AXIMM_66_BREADY(AP_AXIMM_66_BREADY),
        .AP_AXIMM_66_ARADDR(AP_AXIMM_66_ARADDR),
        .AP_AXIMM_66_ARLEN(AP_AXIMM_66_ARLEN),
        .AP_AXIMM_66_ARSIZE(AP_AXIMM_66_ARSIZE),
        .AP_AXIMM_66_ARBURST(AP_AXIMM_66_ARBURST),
        .AP_AXIMM_66_ARLOCK(AP_AXIMM_66_ARLOCK),
        .AP_AXIMM_66_ARCACHE(AP_AXIMM_66_ARCACHE),
        .AP_AXIMM_66_ARPROT(AP_AXIMM_66_ARPROT),
        .AP_AXIMM_66_ARREGION(AP_AXIMM_66_ARREGION),
        .AP_AXIMM_66_ARQOS(AP_AXIMM_66_ARQOS),
        .AP_AXIMM_66_ARVALID(AP_AXIMM_66_ARVALID),
        .AP_AXIMM_66_ARREADY(AP_AXIMM_66_ARREADY),
        .AP_AXIMM_66_RDATA(AP_AXIMM_66_RDATA),
        .AP_AXIMM_66_RRESP(AP_AXIMM_66_RRESP),
        .AP_AXIMM_66_RLAST(AP_AXIMM_66_RLAST),
        .AP_AXIMM_66_RVALID(AP_AXIMM_66_RVALID),
        .AP_AXIMM_66_RREADY(AP_AXIMM_66_RREADY),
        .M_AXIMM_66_AWADDR(M_AXIMM_66_AWADDR),
        .M_AXIMM_66_AWLEN(M_AXIMM_66_AWLEN),
        .M_AXIMM_66_AWSIZE(M_AXIMM_66_AWSIZE),
        .M_AXIMM_66_AWBURST(M_AXIMM_66_AWBURST),
        .M_AXIMM_66_AWLOCK(M_AXIMM_66_AWLOCK),
        .M_AXIMM_66_AWCACHE(M_AXIMM_66_AWCACHE),
        .M_AXIMM_66_AWPROT(M_AXIMM_66_AWPROT),
        .M_AXIMM_66_AWREGION(M_AXIMM_66_AWREGION),
        .M_AXIMM_66_AWQOS(M_AXIMM_66_AWQOS),
        .M_AXIMM_66_AWVALID(M_AXIMM_66_AWVALID),
        .M_AXIMM_66_AWREADY(M_AXIMM_66_AWREADY),
        .M_AXIMM_66_WDATA(M_AXIMM_66_WDATA),
        .M_AXIMM_66_WSTRB(M_AXIMM_66_WSTRB),
        .M_AXIMM_66_WLAST(M_AXIMM_66_WLAST),
        .M_AXIMM_66_WVALID(M_AXIMM_66_WVALID),
        .M_AXIMM_66_WREADY(M_AXIMM_66_WREADY),
        .M_AXIMM_66_BRESP(M_AXIMM_66_BRESP),
        .M_AXIMM_66_BVALID(M_AXIMM_66_BVALID),
        .M_AXIMM_66_BREADY(M_AXIMM_66_BREADY),
        .M_AXIMM_66_ARADDR(M_AXIMM_66_ARADDR),
        .M_AXIMM_66_ARLEN(M_AXIMM_66_ARLEN),
        .M_AXIMM_66_ARSIZE(M_AXIMM_66_ARSIZE),
        .M_AXIMM_66_ARBURST(M_AXIMM_66_ARBURST),
        .M_AXIMM_66_ARLOCK(M_AXIMM_66_ARLOCK),
        .M_AXIMM_66_ARCACHE(M_AXIMM_66_ARCACHE),
        .M_AXIMM_66_ARPROT(M_AXIMM_66_ARPROT),
        .M_AXIMM_66_ARREGION(M_AXIMM_66_ARREGION),
        .M_AXIMM_66_ARQOS(M_AXIMM_66_ARQOS),
        .M_AXIMM_66_ARVALID(M_AXIMM_66_ARVALID),
        .M_AXIMM_66_ARREADY(M_AXIMM_66_ARREADY),
        .M_AXIMM_66_RDATA(M_AXIMM_66_RDATA),
        .M_AXIMM_66_RRESP(M_AXIMM_66_RRESP),
        .M_AXIMM_66_RLAST(M_AXIMM_66_RLAST),
        .M_AXIMM_66_RVALID(M_AXIMM_66_RVALID),
        .M_AXIMM_66_RREADY(M_AXIMM_66_RREADY),
        .AP_AXIMM_67_AWADDR(AP_AXIMM_67_AWADDR),
        .AP_AXIMM_67_AWLEN(AP_AXIMM_67_AWLEN),
        .AP_AXIMM_67_AWSIZE(AP_AXIMM_67_AWSIZE),
        .AP_AXIMM_67_AWBURST(AP_AXIMM_67_AWBURST),
        .AP_AXIMM_67_AWLOCK(AP_AXIMM_67_AWLOCK),
        .AP_AXIMM_67_AWCACHE(AP_AXIMM_67_AWCACHE),
        .AP_AXIMM_67_AWPROT(AP_AXIMM_67_AWPROT),
        .AP_AXIMM_67_AWREGION(AP_AXIMM_67_AWREGION),
        .AP_AXIMM_67_AWQOS(AP_AXIMM_67_AWQOS),
        .AP_AXIMM_67_AWVALID(AP_AXIMM_67_AWVALID),
        .AP_AXIMM_67_AWREADY(AP_AXIMM_67_AWREADY),
        .AP_AXIMM_67_WDATA(AP_AXIMM_67_WDATA),
        .AP_AXIMM_67_WSTRB(AP_AXIMM_67_WSTRB),
        .AP_AXIMM_67_WLAST(AP_AXIMM_67_WLAST),
        .AP_AXIMM_67_WVALID(AP_AXIMM_67_WVALID),
        .AP_AXIMM_67_WREADY(AP_AXIMM_67_WREADY),
        .AP_AXIMM_67_BRESP(AP_AXIMM_67_BRESP),
        .AP_AXIMM_67_BVALID(AP_AXIMM_67_BVALID),
        .AP_AXIMM_67_BREADY(AP_AXIMM_67_BREADY),
        .AP_AXIMM_67_ARADDR(AP_AXIMM_67_ARADDR),
        .AP_AXIMM_67_ARLEN(AP_AXIMM_67_ARLEN),
        .AP_AXIMM_67_ARSIZE(AP_AXIMM_67_ARSIZE),
        .AP_AXIMM_67_ARBURST(AP_AXIMM_67_ARBURST),
        .AP_AXIMM_67_ARLOCK(AP_AXIMM_67_ARLOCK),
        .AP_AXIMM_67_ARCACHE(AP_AXIMM_67_ARCACHE),
        .AP_AXIMM_67_ARPROT(AP_AXIMM_67_ARPROT),
        .AP_AXIMM_67_ARREGION(AP_AXIMM_67_ARREGION),
        .AP_AXIMM_67_ARQOS(AP_AXIMM_67_ARQOS),
        .AP_AXIMM_67_ARVALID(AP_AXIMM_67_ARVALID),
        .AP_AXIMM_67_ARREADY(AP_AXIMM_67_ARREADY),
        .AP_AXIMM_67_RDATA(AP_AXIMM_67_RDATA),
        .AP_AXIMM_67_RRESP(AP_AXIMM_67_RRESP),
        .AP_AXIMM_67_RLAST(AP_AXIMM_67_RLAST),
        .AP_AXIMM_67_RVALID(AP_AXIMM_67_RVALID),
        .AP_AXIMM_67_RREADY(AP_AXIMM_67_RREADY),
        .M_AXIMM_67_AWADDR(M_AXIMM_67_AWADDR),
        .M_AXIMM_67_AWLEN(M_AXIMM_67_AWLEN),
        .M_AXIMM_67_AWSIZE(M_AXIMM_67_AWSIZE),
        .M_AXIMM_67_AWBURST(M_AXIMM_67_AWBURST),
        .M_AXIMM_67_AWLOCK(M_AXIMM_67_AWLOCK),
        .M_AXIMM_67_AWCACHE(M_AXIMM_67_AWCACHE),
        .M_AXIMM_67_AWPROT(M_AXIMM_67_AWPROT),
        .M_AXIMM_67_AWREGION(M_AXIMM_67_AWREGION),
        .M_AXIMM_67_AWQOS(M_AXIMM_67_AWQOS),
        .M_AXIMM_67_AWVALID(M_AXIMM_67_AWVALID),
        .M_AXIMM_67_AWREADY(M_AXIMM_67_AWREADY),
        .M_AXIMM_67_WDATA(M_AXIMM_67_WDATA),
        .M_AXIMM_67_WSTRB(M_AXIMM_67_WSTRB),
        .M_AXIMM_67_WLAST(M_AXIMM_67_WLAST),
        .M_AXIMM_67_WVALID(M_AXIMM_67_WVALID),
        .M_AXIMM_67_WREADY(M_AXIMM_67_WREADY),
        .M_AXIMM_67_BRESP(M_AXIMM_67_BRESP),
        .M_AXIMM_67_BVALID(M_AXIMM_67_BVALID),
        .M_AXIMM_67_BREADY(M_AXIMM_67_BREADY),
        .M_AXIMM_67_ARADDR(M_AXIMM_67_ARADDR),
        .M_AXIMM_67_ARLEN(M_AXIMM_67_ARLEN),
        .M_AXIMM_67_ARSIZE(M_AXIMM_67_ARSIZE),
        .M_AXIMM_67_ARBURST(M_AXIMM_67_ARBURST),
        .M_AXIMM_67_ARLOCK(M_AXIMM_67_ARLOCK),
        .M_AXIMM_67_ARCACHE(M_AXIMM_67_ARCACHE),
        .M_AXIMM_67_ARPROT(M_AXIMM_67_ARPROT),
        .M_AXIMM_67_ARREGION(M_AXIMM_67_ARREGION),
        .M_AXIMM_67_ARQOS(M_AXIMM_67_ARQOS),
        .M_AXIMM_67_ARVALID(M_AXIMM_67_ARVALID),
        .M_AXIMM_67_ARREADY(M_AXIMM_67_ARREADY),
        .M_AXIMM_67_RDATA(M_AXIMM_67_RDATA),
        .M_AXIMM_67_RRESP(M_AXIMM_67_RRESP),
        .M_AXIMM_67_RLAST(M_AXIMM_67_RLAST),
        .M_AXIMM_67_RVALID(M_AXIMM_67_RVALID),
        .M_AXIMM_67_RREADY(M_AXIMM_67_RREADY),
        .AP_AXIMM_68_AWADDR(AP_AXIMM_68_AWADDR),
        .AP_AXIMM_68_AWLEN(AP_AXIMM_68_AWLEN),
        .AP_AXIMM_68_AWSIZE(AP_AXIMM_68_AWSIZE),
        .AP_AXIMM_68_AWBURST(AP_AXIMM_68_AWBURST),
        .AP_AXIMM_68_AWLOCK(AP_AXIMM_68_AWLOCK),
        .AP_AXIMM_68_AWCACHE(AP_AXIMM_68_AWCACHE),
        .AP_AXIMM_68_AWPROT(AP_AXIMM_68_AWPROT),
        .AP_AXIMM_68_AWREGION(AP_AXIMM_68_AWREGION),
        .AP_AXIMM_68_AWQOS(AP_AXIMM_68_AWQOS),
        .AP_AXIMM_68_AWVALID(AP_AXIMM_68_AWVALID),
        .AP_AXIMM_68_AWREADY(AP_AXIMM_68_AWREADY),
        .AP_AXIMM_68_WDATA(AP_AXIMM_68_WDATA),
        .AP_AXIMM_68_WSTRB(AP_AXIMM_68_WSTRB),
        .AP_AXIMM_68_WLAST(AP_AXIMM_68_WLAST),
        .AP_AXIMM_68_WVALID(AP_AXIMM_68_WVALID),
        .AP_AXIMM_68_WREADY(AP_AXIMM_68_WREADY),
        .AP_AXIMM_68_BRESP(AP_AXIMM_68_BRESP),
        .AP_AXIMM_68_BVALID(AP_AXIMM_68_BVALID),
        .AP_AXIMM_68_BREADY(AP_AXIMM_68_BREADY),
        .AP_AXIMM_68_ARADDR(AP_AXIMM_68_ARADDR),
        .AP_AXIMM_68_ARLEN(AP_AXIMM_68_ARLEN),
        .AP_AXIMM_68_ARSIZE(AP_AXIMM_68_ARSIZE),
        .AP_AXIMM_68_ARBURST(AP_AXIMM_68_ARBURST),
        .AP_AXIMM_68_ARLOCK(AP_AXIMM_68_ARLOCK),
        .AP_AXIMM_68_ARCACHE(AP_AXIMM_68_ARCACHE),
        .AP_AXIMM_68_ARPROT(AP_AXIMM_68_ARPROT),
        .AP_AXIMM_68_ARREGION(AP_AXIMM_68_ARREGION),
        .AP_AXIMM_68_ARQOS(AP_AXIMM_68_ARQOS),
        .AP_AXIMM_68_ARVALID(AP_AXIMM_68_ARVALID),
        .AP_AXIMM_68_ARREADY(AP_AXIMM_68_ARREADY),
        .AP_AXIMM_68_RDATA(AP_AXIMM_68_RDATA),
        .AP_AXIMM_68_RRESP(AP_AXIMM_68_RRESP),
        .AP_AXIMM_68_RLAST(AP_AXIMM_68_RLAST),
        .AP_AXIMM_68_RVALID(AP_AXIMM_68_RVALID),
        .AP_AXIMM_68_RREADY(AP_AXIMM_68_RREADY),
        .M_AXIMM_68_AWADDR(M_AXIMM_68_AWADDR),
        .M_AXIMM_68_AWLEN(M_AXIMM_68_AWLEN),
        .M_AXIMM_68_AWSIZE(M_AXIMM_68_AWSIZE),
        .M_AXIMM_68_AWBURST(M_AXIMM_68_AWBURST),
        .M_AXIMM_68_AWLOCK(M_AXIMM_68_AWLOCK),
        .M_AXIMM_68_AWCACHE(M_AXIMM_68_AWCACHE),
        .M_AXIMM_68_AWPROT(M_AXIMM_68_AWPROT),
        .M_AXIMM_68_AWREGION(M_AXIMM_68_AWREGION),
        .M_AXIMM_68_AWQOS(M_AXIMM_68_AWQOS),
        .M_AXIMM_68_AWVALID(M_AXIMM_68_AWVALID),
        .M_AXIMM_68_AWREADY(M_AXIMM_68_AWREADY),
        .M_AXIMM_68_WDATA(M_AXIMM_68_WDATA),
        .M_AXIMM_68_WSTRB(M_AXIMM_68_WSTRB),
        .M_AXIMM_68_WLAST(M_AXIMM_68_WLAST),
        .M_AXIMM_68_WVALID(M_AXIMM_68_WVALID),
        .M_AXIMM_68_WREADY(M_AXIMM_68_WREADY),
        .M_AXIMM_68_BRESP(M_AXIMM_68_BRESP),
        .M_AXIMM_68_BVALID(M_AXIMM_68_BVALID),
        .M_AXIMM_68_BREADY(M_AXIMM_68_BREADY),
        .M_AXIMM_68_ARADDR(M_AXIMM_68_ARADDR),
        .M_AXIMM_68_ARLEN(M_AXIMM_68_ARLEN),
        .M_AXIMM_68_ARSIZE(M_AXIMM_68_ARSIZE),
        .M_AXIMM_68_ARBURST(M_AXIMM_68_ARBURST),
        .M_AXIMM_68_ARLOCK(M_AXIMM_68_ARLOCK),
        .M_AXIMM_68_ARCACHE(M_AXIMM_68_ARCACHE),
        .M_AXIMM_68_ARPROT(M_AXIMM_68_ARPROT),
        .M_AXIMM_68_ARREGION(M_AXIMM_68_ARREGION),
        .M_AXIMM_68_ARQOS(M_AXIMM_68_ARQOS),
        .M_AXIMM_68_ARVALID(M_AXIMM_68_ARVALID),
        .M_AXIMM_68_ARREADY(M_AXIMM_68_ARREADY),
        .M_AXIMM_68_RDATA(M_AXIMM_68_RDATA),
        .M_AXIMM_68_RRESP(M_AXIMM_68_RRESP),
        .M_AXIMM_68_RLAST(M_AXIMM_68_RLAST),
        .M_AXIMM_68_RVALID(M_AXIMM_68_RVALID),
        .M_AXIMM_68_RREADY(M_AXIMM_68_RREADY),
        .AP_AXIMM_69_AWADDR(AP_AXIMM_69_AWADDR),
        .AP_AXIMM_69_AWLEN(AP_AXIMM_69_AWLEN),
        .AP_AXIMM_69_AWSIZE(AP_AXIMM_69_AWSIZE),
        .AP_AXIMM_69_AWBURST(AP_AXIMM_69_AWBURST),
        .AP_AXIMM_69_AWLOCK(AP_AXIMM_69_AWLOCK),
        .AP_AXIMM_69_AWCACHE(AP_AXIMM_69_AWCACHE),
        .AP_AXIMM_69_AWPROT(AP_AXIMM_69_AWPROT),
        .AP_AXIMM_69_AWREGION(AP_AXIMM_69_AWREGION),
        .AP_AXIMM_69_AWQOS(AP_AXIMM_69_AWQOS),
        .AP_AXIMM_69_AWVALID(AP_AXIMM_69_AWVALID),
        .AP_AXIMM_69_AWREADY(AP_AXIMM_69_AWREADY),
        .AP_AXIMM_69_WDATA(AP_AXIMM_69_WDATA),
        .AP_AXIMM_69_WSTRB(AP_AXIMM_69_WSTRB),
        .AP_AXIMM_69_WLAST(AP_AXIMM_69_WLAST),
        .AP_AXIMM_69_WVALID(AP_AXIMM_69_WVALID),
        .AP_AXIMM_69_WREADY(AP_AXIMM_69_WREADY),
        .AP_AXIMM_69_BRESP(AP_AXIMM_69_BRESP),
        .AP_AXIMM_69_BVALID(AP_AXIMM_69_BVALID),
        .AP_AXIMM_69_BREADY(AP_AXIMM_69_BREADY),
        .AP_AXIMM_69_ARADDR(AP_AXIMM_69_ARADDR),
        .AP_AXIMM_69_ARLEN(AP_AXIMM_69_ARLEN),
        .AP_AXIMM_69_ARSIZE(AP_AXIMM_69_ARSIZE),
        .AP_AXIMM_69_ARBURST(AP_AXIMM_69_ARBURST),
        .AP_AXIMM_69_ARLOCK(AP_AXIMM_69_ARLOCK),
        .AP_AXIMM_69_ARCACHE(AP_AXIMM_69_ARCACHE),
        .AP_AXIMM_69_ARPROT(AP_AXIMM_69_ARPROT),
        .AP_AXIMM_69_ARREGION(AP_AXIMM_69_ARREGION),
        .AP_AXIMM_69_ARQOS(AP_AXIMM_69_ARQOS),
        .AP_AXIMM_69_ARVALID(AP_AXIMM_69_ARVALID),
        .AP_AXIMM_69_ARREADY(AP_AXIMM_69_ARREADY),
        .AP_AXIMM_69_RDATA(AP_AXIMM_69_RDATA),
        .AP_AXIMM_69_RRESP(AP_AXIMM_69_RRESP),
        .AP_AXIMM_69_RLAST(AP_AXIMM_69_RLAST),
        .AP_AXIMM_69_RVALID(AP_AXIMM_69_RVALID),
        .AP_AXIMM_69_RREADY(AP_AXIMM_69_RREADY),
        .M_AXIMM_69_AWADDR(M_AXIMM_69_AWADDR),
        .M_AXIMM_69_AWLEN(M_AXIMM_69_AWLEN),
        .M_AXIMM_69_AWSIZE(M_AXIMM_69_AWSIZE),
        .M_AXIMM_69_AWBURST(M_AXIMM_69_AWBURST),
        .M_AXIMM_69_AWLOCK(M_AXIMM_69_AWLOCK),
        .M_AXIMM_69_AWCACHE(M_AXIMM_69_AWCACHE),
        .M_AXIMM_69_AWPROT(M_AXIMM_69_AWPROT),
        .M_AXIMM_69_AWREGION(M_AXIMM_69_AWREGION),
        .M_AXIMM_69_AWQOS(M_AXIMM_69_AWQOS),
        .M_AXIMM_69_AWVALID(M_AXIMM_69_AWVALID),
        .M_AXIMM_69_AWREADY(M_AXIMM_69_AWREADY),
        .M_AXIMM_69_WDATA(M_AXIMM_69_WDATA),
        .M_AXIMM_69_WSTRB(M_AXIMM_69_WSTRB),
        .M_AXIMM_69_WLAST(M_AXIMM_69_WLAST),
        .M_AXIMM_69_WVALID(M_AXIMM_69_WVALID),
        .M_AXIMM_69_WREADY(M_AXIMM_69_WREADY),
        .M_AXIMM_69_BRESP(M_AXIMM_69_BRESP),
        .M_AXIMM_69_BVALID(M_AXIMM_69_BVALID),
        .M_AXIMM_69_BREADY(M_AXIMM_69_BREADY),
        .M_AXIMM_69_ARADDR(M_AXIMM_69_ARADDR),
        .M_AXIMM_69_ARLEN(M_AXIMM_69_ARLEN),
        .M_AXIMM_69_ARSIZE(M_AXIMM_69_ARSIZE),
        .M_AXIMM_69_ARBURST(M_AXIMM_69_ARBURST),
        .M_AXIMM_69_ARLOCK(M_AXIMM_69_ARLOCK),
        .M_AXIMM_69_ARCACHE(M_AXIMM_69_ARCACHE),
        .M_AXIMM_69_ARPROT(M_AXIMM_69_ARPROT),
        .M_AXIMM_69_ARREGION(M_AXIMM_69_ARREGION),
        .M_AXIMM_69_ARQOS(M_AXIMM_69_ARQOS),
        .M_AXIMM_69_ARVALID(M_AXIMM_69_ARVALID),
        .M_AXIMM_69_ARREADY(M_AXIMM_69_ARREADY),
        .M_AXIMM_69_RDATA(M_AXIMM_69_RDATA),
        .M_AXIMM_69_RRESP(M_AXIMM_69_RRESP),
        .M_AXIMM_69_RLAST(M_AXIMM_69_RLAST),
        .M_AXIMM_69_RVALID(M_AXIMM_69_RVALID),
        .M_AXIMM_69_RREADY(M_AXIMM_69_RREADY),
        .AP_AXIMM_70_AWADDR(AP_AXIMM_70_AWADDR),
        .AP_AXIMM_70_AWLEN(AP_AXIMM_70_AWLEN),
        .AP_AXIMM_70_AWSIZE(AP_AXIMM_70_AWSIZE),
        .AP_AXIMM_70_AWBURST(AP_AXIMM_70_AWBURST),
        .AP_AXIMM_70_AWLOCK(AP_AXIMM_70_AWLOCK),
        .AP_AXIMM_70_AWCACHE(AP_AXIMM_70_AWCACHE),
        .AP_AXIMM_70_AWPROT(AP_AXIMM_70_AWPROT),
        .AP_AXIMM_70_AWREGION(AP_AXIMM_70_AWREGION),
        .AP_AXIMM_70_AWQOS(AP_AXIMM_70_AWQOS),
        .AP_AXIMM_70_AWVALID(AP_AXIMM_70_AWVALID),
        .AP_AXIMM_70_AWREADY(AP_AXIMM_70_AWREADY),
        .AP_AXIMM_70_WDATA(AP_AXIMM_70_WDATA),
        .AP_AXIMM_70_WSTRB(AP_AXIMM_70_WSTRB),
        .AP_AXIMM_70_WLAST(AP_AXIMM_70_WLAST),
        .AP_AXIMM_70_WVALID(AP_AXIMM_70_WVALID),
        .AP_AXIMM_70_WREADY(AP_AXIMM_70_WREADY),
        .AP_AXIMM_70_BRESP(AP_AXIMM_70_BRESP),
        .AP_AXIMM_70_BVALID(AP_AXIMM_70_BVALID),
        .AP_AXIMM_70_BREADY(AP_AXIMM_70_BREADY),
        .AP_AXIMM_70_ARADDR(AP_AXIMM_70_ARADDR),
        .AP_AXIMM_70_ARLEN(AP_AXIMM_70_ARLEN),
        .AP_AXIMM_70_ARSIZE(AP_AXIMM_70_ARSIZE),
        .AP_AXIMM_70_ARBURST(AP_AXIMM_70_ARBURST),
        .AP_AXIMM_70_ARLOCK(AP_AXIMM_70_ARLOCK),
        .AP_AXIMM_70_ARCACHE(AP_AXIMM_70_ARCACHE),
        .AP_AXIMM_70_ARPROT(AP_AXIMM_70_ARPROT),
        .AP_AXIMM_70_ARREGION(AP_AXIMM_70_ARREGION),
        .AP_AXIMM_70_ARQOS(AP_AXIMM_70_ARQOS),
        .AP_AXIMM_70_ARVALID(AP_AXIMM_70_ARVALID),
        .AP_AXIMM_70_ARREADY(AP_AXIMM_70_ARREADY),
        .AP_AXIMM_70_RDATA(AP_AXIMM_70_RDATA),
        .AP_AXIMM_70_RRESP(AP_AXIMM_70_RRESP),
        .AP_AXIMM_70_RLAST(AP_AXIMM_70_RLAST),
        .AP_AXIMM_70_RVALID(AP_AXIMM_70_RVALID),
        .AP_AXIMM_70_RREADY(AP_AXIMM_70_RREADY),
        .M_AXIMM_70_AWADDR(M_AXIMM_70_AWADDR),
        .M_AXIMM_70_AWLEN(M_AXIMM_70_AWLEN),
        .M_AXIMM_70_AWSIZE(M_AXIMM_70_AWSIZE),
        .M_AXIMM_70_AWBURST(M_AXIMM_70_AWBURST),
        .M_AXIMM_70_AWLOCK(M_AXIMM_70_AWLOCK),
        .M_AXIMM_70_AWCACHE(M_AXIMM_70_AWCACHE),
        .M_AXIMM_70_AWPROT(M_AXIMM_70_AWPROT),
        .M_AXIMM_70_AWREGION(M_AXIMM_70_AWREGION),
        .M_AXIMM_70_AWQOS(M_AXIMM_70_AWQOS),
        .M_AXIMM_70_AWVALID(M_AXIMM_70_AWVALID),
        .M_AXIMM_70_AWREADY(M_AXIMM_70_AWREADY),
        .M_AXIMM_70_WDATA(M_AXIMM_70_WDATA),
        .M_AXIMM_70_WSTRB(M_AXIMM_70_WSTRB),
        .M_AXIMM_70_WLAST(M_AXIMM_70_WLAST),
        .M_AXIMM_70_WVALID(M_AXIMM_70_WVALID),
        .M_AXIMM_70_WREADY(M_AXIMM_70_WREADY),
        .M_AXIMM_70_BRESP(M_AXIMM_70_BRESP),
        .M_AXIMM_70_BVALID(M_AXIMM_70_BVALID),
        .M_AXIMM_70_BREADY(M_AXIMM_70_BREADY),
        .M_AXIMM_70_ARADDR(M_AXIMM_70_ARADDR),
        .M_AXIMM_70_ARLEN(M_AXIMM_70_ARLEN),
        .M_AXIMM_70_ARSIZE(M_AXIMM_70_ARSIZE),
        .M_AXIMM_70_ARBURST(M_AXIMM_70_ARBURST),
        .M_AXIMM_70_ARLOCK(M_AXIMM_70_ARLOCK),
        .M_AXIMM_70_ARCACHE(M_AXIMM_70_ARCACHE),
        .M_AXIMM_70_ARPROT(M_AXIMM_70_ARPROT),
        .M_AXIMM_70_ARREGION(M_AXIMM_70_ARREGION),
        .M_AXIMM_70_ARQOS(M_AXIMM_70_ARQOS),
        .M_AXIMM_70_ARVALID(M_AXIMM_70_ARVALID),
        .M_AXIMM_70_ARREADY(M_AXIMM_70_ARREADY),
        .M_AXIMM_70_RDATA(M_AXIMM_70_RDATA),
        .M_AXIMM_70_RRESP(M_AXIMM_70_RRESP),
        .M_AXIMM_70_RLAST(M_AXIMM_70_RLAST),
        .M_AXIMM_70_RVALID(M_AXIMM_70_RVALID),
        .M_AXIMM_70_RREADY(M_AXIMM_70_RREADY),
        .AP_AXIMM_71_AWADDR(AP_AXIMM_71_AWADDR),
        .AP_AXIMM_71_AWLEN(AP_AXIMM_71_AWLEN),
        .AP_AXIMM_71_AWSIZE(AP_AXIMM_71_AWSIZE),
        .AP_AXIMM_71_AWBURST(AP_AXIMM_71_AWBURST),
        .AP_AXIMM_71_AWLOCK(AP_AXIMM_71_AWLOCK),
        .AP_AXIMM_71_AWCACHE(AP_AXIMM_71_AWCACHE),
        .AP_AXIMM_71_AWPROT(AP_AXIMM_71_AWPROT),
        .AP_AXIMM_71_AWREGION(AP_AXIMM_71_AWREGION),
        .AP_AXIMM_71_AWQOS(AP_AXIMM_71_AWQOS),
        .AP_AXIMM_71_AWVALID(AP_AXIMM_71_AWVALID),
        .AP_AXIMM_71_AWREADY(AP_AXIMM_71_AWREADY),
        .AP_AXIMM_71_WDATA(AP_AXIMM_71_WDATA),
        .AP_AXIMM_71_WSTRB(AP_AXIMM_71_WSTRB),
        .AP_AXIMM_71_WLAST(AP_AXIMM_71_WLAST),
        .AP_AXIMM_71_WVALID(AP_AXIMM_71_WVALID),
        .AP_AXIMM_71_WREADY(AP_AXIMM_71_WREADY),
        .AP_AXIMM_71_BRESP(AP_AXIMM_71_BRESP),
        .AP_AXIMM_71_BVALID(AP_AXIMM_71_BVALID),
        .AP_AXIMM_71_BREADY(AP_AXIMM_71_BREADY),
        .AP_AXIMM_71_ARADDR(AP_AXIMM_71_ARADDR),
        .AP_AXIMM_71_ARLEN(AP_AXIMM_71_ARLEN),
        .AP_AXIMM_71_ARSIZE(AP_AXIMM_71_ARSIZE),
        .AP_AXIMM_71_ARBURST(AP_AXIMM_71_ARBURST),
        .AP_AXIMM_71_ARLOCK(AP_AXIMM_71_ARLOCK),
        .AP_AXIMM_71_ARCACHE(AP_AXIMM_71_ARCACHE),
        .AP_AXIMM_71_ARPROT(AP_AXIMM_71_ARPROT),
        .AP_AXIMM_71_ARREGION(AP_AXIMM_71_ARREGION),
        .AP_AXIMM_71_ARQOS(AP_AXIMM_71_ARQOS),
        .AP_AXIMM_71_ARVALID(AP_AXIMM_71_ARVALID),
        .AP_AXIMM_71_ARREADY(AP_AXIMM_71_ARREADY),
        .AP_AXIMM_71_RDATA(AP_AXIMM_71_RDATA),
        .AP_AXIMM_71_RRESP(AP_AXIMM_71_RRESP),
        .AP_AXIMM_71_RLAST(AP_AXIMM_71_RLAST),
        .AP_AXIMM_71_RVALID(AP_AXIMM_71_RVALID),
        .AP_AXIMM_71_RREADY(AP_AXIMM_71_RREADY),
        .M_AXIMM_71_AWADDR(M_AXIMM_71_AWADDR),
        .M_AXIMM_71_AWLEN(M_AXIMM_71_AWLEN),
        .M_AXIMM_71_AWSIZE(M_AXIMM_71_AWSIZE),
        .M_AXIMM_71_AWBURST(M_AXIMM_71_AWBURST),
        .M_AXIMM_71_AWLOCK(M_AXIMM_71_AWLOCK),
        .M_AXIMM_71_AWCACHE(M_AXIMM_71_AWCACHE),
        .M_AXIMM_71_AWPROT(M_AXIMM_71_AWPROT),
        .M_AXIMM_71_AWREGION(M_AXIMM_71_AWREGION),
        .M_AXIMM_71_AWQOS(M_AXIMM_71_AWQOS),
        .M_AXIMM_71_AWVALID(M_AXIMM_71_AWVALID),
        .M_AXIMM_71_AWREADY(M_AXIMM_71_AWREADY),
        .M_AXIMM_71_WDATA(M_AXIMM_71_WDATA),
        .M_AXIMM_71_WSTRB(M_AXIMM_71_WSTRB),
        .M_AXIMM_71_WLAST(M_AXIMM_71_WLAST),
        .M_AXIMM_71_WVALID(M_AXIMM_71_WVALID),
        .M_AXIMM_71_WREADY(M_AXIMM_71_WREADY),
        .M_AXIMM_71_BRESP(M_AXIMM_71_BRESP),
        .M_AXIMM_71_BVALID(M_AXIMM_71_BVALID),
        .M_AXIMM_71_BREADY(M_AXIMM_71_BREADY),
        .M_AXIMM_71_ARADDR(M_AXIMM_71_ARADDR),
        .M_AXIMM_71_ARLEN(M_AXIMM_71_ARLEN),
        .M_AXIMM_71_ARSIZE(M_AXIMM_71_ARSIZE),
        .M_AXIMM_71_ARBURST(M_AXIMM_71_ARBURST),
        .M_AXIMM_71_ARLOCK(M_AXIMM_71_ARLOCK),
        .M_AXIMM_71_ARCACHE(M_AXIMM_71_ARCACHE),
        .M_AXIMM_71_ARPROT(M_AXIMM_71_ARPROT),
        .M_AXIMM_71_ARREGION(M_AXIMM_71_ARREGION),
        .M_AXIMM_71_ARQOS(M_AXIMM_71_ARQOS),
        .M_AXIMM_71_ARVALID(M_AXIMM_71_ARVALID),
        .M_AXIMM_71_ARREADY(M_AXIMM_71_ARREADY),
        .M_AXIMM_71_RDATA(M_AXIMM_71_RDATA),
        .M_AXIMM_71_RRESP(M_AXIMM_71_RRESP),
        .M_AXIMM_71_RLAST(M_AXIMM_71_RLAST),
        .M_AXIMM_71_RVALID(M_AXIMM_71_RVALID),
        .M_AXIMM_71_RREADY(M_AXIMM_71_RREADY),
        .AP_AXIMM_72_AWADDR(AP_AXIMM_72_AWADDR),
        .AP_AXIMM_72_AWLEN(AP_AXIMM_72_AWLEN),
        .AP_AXIMM_72_AWSIZE(AP_AXIMM_72_AWSIZE),
        .AP_AXIMM_72_AWBURST(AP_AXIMM_72_AWBURST),
        .AP_AXIMM_72_AWLOCK(AP_AXIMM_72_AWLOCK),
        .AP_AXIMM_72_AWCACHE(AP_AXIMM_72_AWCACHE),
        .AP_AXIMM_72_AWPROT(AP_AXIMM_72_AWPROT),
        .AP_AXIMM_72_AWREGION(AP_AXIMM_72_AWREGION),
        .AP_AXIMM_72_AWQOS(AP_AXIMM_72_AWQOS),
        .AP_AXIMM_72_AWVALID(AP_AXIMM_72_AWVALID),
        .AP_AXIMM_72_AWREADY(AP_AXIMM_72_AWREADY),
        .AP_AXIMM_72_WDATA(AP_AXIMM_72_WDATA),
        .AP_AXIMM_72_WSTRB(AP_AXIMM_72_WSTRB),
        .AP_AXIMM_72_WLAST(AP_AXIMM_72_WLAST),
        .AP_AXIMM_72_WVALID(AP_AXIMM_72_WVALID),
        .AP_AXIMM_72_WREADY(AP_AXIMM_72_WREADY),
        .AP_AXIMM_72_BRESP(AP_AXIMM_72_BRESP),
        .AP_AXIMM_72_BVALID(AP_AXIMM_72_BVALID),
        .AP_AXIMM_72_BREADY(AP_AXIMM_72_BREADY),
        .AP_AXIMM_72_ARADDR(AP_AXIMM_72_ARADDR),
        .AP_AXIMM_72_ARLEN(AP_AXIMM_72_ARLEN),
        .AP_AXIMM_72_ARSIZE(AP_AXIMM_72_ARSIZE),
        .AP_AXIMM_72_ARBURST(AP_AXIMM_72_ARBURST),
        .AP_AXIMM_72_ARLOCK(AP_AXIMM_72_ARLOCK),
        .AP_AXIMM_72_ARCACHE(AP_AXIMM_72_ARCACHE),
        .AP_AXIMM_72_ARPROT(AP_AXIMM_72_ARPROT),
        .AP_AXIMM_72_ARREGION(AP_AXIMM_72_ARREGION),
        .AP_AXIMM_72_ARQOS(AP_AXIMM_72_ARQOS),
        .AP_AXIMM_72_ARVALID(AP_AXIMM_72_ARVALID),
        .AP_AXIMM_72_ARREADY(AP_AXIMM_72_ARREADY),
        .AP_AXIMM_72_RDATA(AP_AXIMM_72_RDATA),
        .AP_AXIMM_72_RRESP(AP_AXIMM_72_RRESP),
        .AP_AXIMM_72_RLAST(AP_AXIMM_72_RLAST),
        .AP_AXIMM_72_RVALID(AP_AXIMM_72_RVALID),
        .AP_AXIMM_72_RREADY(AP_AXIMM_72_RREADY),
        .M_AXIMM_72_AWADDR(M_AXIMM_72_AWADDR),
        .M_AXIMM_72_AWLEN(M_AXIMM_72_AWLEN),
        .M_AXIMM_72_AWSIZE(M_AXIMM_72_AWSIZE),
        .M_AXIMM_72_AWBURST(M_AXIMM_72_AWBURST),
        .M_AXIMM_72_AWLOCK(M_AXIMM_72_AWLOCK),
        .M_AXIMM_72_AWCACHE(M_AXIMM_72_AWCACHE),
        .M_AXIMM_72_AWPROT(M_AXIMM_72_AWPROT),
        .M_AXIMM_72_AWREGION(M_AXIMM_72_AWREGION),
        .M_AXIMM_72_AWQOS(M_AXIMM_72_AWQOS),
        .M_AXIMM_72_AWVALID(M_AXIMM_72_AWVALID),
        .M_AXIMM_72_AWREADY(M_AXIMM_72_AWREADY),
        .M_AXIMM_72_WDATA(M_AXIMM_72_WDATA),
        .M_AXIMM_72_WSTRB(M_AXIMM_72_WSTRB),
        .M_AXIMM_72_WLAST(M_AXIMM_72_WLAST),
        .M_AXIMM_72_WVALID(M_AXIMM_72_WVALID),
        .M_AXIMM_72_WREADY(M_AXIMM_72_WREADY),
        .M_AXIMM_72_BRESP(M_AXIMM_72_BRESP),
        .M_AXIMM_72_BVALID(M_AXIMM_72_BVALID),
        .M_AXIMM_72_BREADY(M_AXIMM_72_BREADY),
        .M_AXIMM_72_ARADDR(M_AXIMM_72_ARADDR),
        .M_AXIMM_72_ARLEN(M_AXIMM_72_ARLEN),
        .M_AXIMM_72_ARSIZE(M_AXIMM_72_ARSIZE),
        .M_AXIMM_72_ARBURST(M_AXIMM_72_ARBURST),
        .M_AXIMM_72_ARLOCK(M_AXIMM_72_ARLOCK),
        .M_AXIMM_72_ARCACHE(M_AXIMM_72_ARCACHE),
        .M_AXIMM_72_ARPROT(M_AXIMM_72_ARPROT),
        .M_AXIMM_72_ARREGION(M_AXIMM_72_ARREGION),
        .M_AXIMM_72_ARQOS(M_AXIMM_72_ARQOS),
        .M_AXIMM_72_ARVALID(M_AXIMM_72_ARVALID),
        .M_AXIMM_72_ARREADY(M_AXIMM_72_ARREADY),
        .M_AXIMM_72_RDATA(M_AXIMM_72_RDATA),
        .M_AXIMM_72_RRESP(M_AXIMM_72_RRESP),
        .M_AXIMM_72_RLAST(M_AXIMM_72_RLAST),
        .M_AXIMM_72_RVALID(M_AXIMM_72_RVALID),
        .M_AXIMM_72_RREADY(M_AXIMM_72_RREADY),
        .AP_AXIMM_73_AWADDR(AP_AXIMM_73_AWADDR),
        .AP_AXIMM_73_AWLEN(AP_AXIMM_73_AWLEN),
        .AP_AXIMM_73_AWSIZE(AP_AXIMM_73_AWSIZE),
        .AP_AXIMM_73_AWBURST(AP_AXIMM_73_AWBURST),
        .AP_AXIMM_73_AWLOCK(AP_AXIMM_73_AWLOCK),
        .AP_AXIMM_73_AWCACHE(AP_AXIMM_73_AWCACHE),
        .AP_AXIMM_73_AWPROT(AP_AXIMM_73_AWPROT),
        .AP_AXIMM_73_AWREGION(AP_AXIMM_73_AWREGION),
        .AP_AXIMM_73_AWQOS(AP_AXIMM_73_AWQOS),
        .AP_AXIMM_73_AWVALID(AP_AXIMM_73_AWVALID),
        .AP_AXIMM_73_AWREADY(AP_AXIMM_73_AWREADY),
        .AP_AXIMM_73_WDATA(AP_AXIMM_73_WDATA),
        .AP_AXIMM_73_WSTRB(AP_AXIMM_73_WSTRB),
        .AP_AXIMM_73_WLAST(AP_AXIMM_73_WLAST),
        .AP_AXIMM_73_WVALID(AP_AXIMM_73_WVALID),
        .AP_AXIMM_73_WREADY(AP_AXIMM_73_WREADY),
        .AP_AXIMM_73_BRESP(AP_AXIMM_73_BRESP),
        .AP_AXIMM_73_BVALID(AP_AXIMM_73_BVALID),
        .AP_AXIMM_73_BREADY(AP_AXIMM_73_BREADY),
        .AP_AXIMM_73_ARADDR(AP_AXIMM_73_ARADDR),
        .AP_AXIMM_73_ARLEN(AP_AXIMM_73_ARLEN),
        .AP_AXIMM_73_ARSIZE(AP_AXIMM_73_ARSIZE),
        .AP_AXIMM_73_ARBURST(AP_AXIMM_73_ARBURST),
        .AP_AXIMM_73_ARLOCK(AP_AXIMM_73_ARLOCK),
        .AP_AXIMM_73_ARCACHE(AP_AXIMM_73_ARCACHE),
        .AP_AXIMM_73_ARPROT(AP_AXIMM_73_ARPROT),
        .AP_AXIMM_73_ARREGION(AP_AXIMM_73_ARREGION),
        .AP_AXIMM_73_ARQOS(AP_AXIMM_73_ARQOS),
        .AP_AXIMM_73_ARVALID(AP_AXIMM_73_ARVALID),
        .AP_AXIMM_73_ARREADY(AP_AXIMM_73_ARREADY),
        .AP_AXIMM_73_RDATA(AP_AXIMM_73_RDATA),
        .AP_AXIMM_73_RRESP(AP_AXIMM_73_RRESP),
        .AP_AXIMM_73_RLAST(AP_AXIMM_73_RLAST),
        .AP_AXIMM_73_RVALID(AP_AXIMM_73_RVALID),
        .AP_AXIMM_73_RREADY(AP_AXIMM_73_RREADY),
        .M_AXIMM_73_AWADDR(M_AXIMM_73_AWADDR),
        .M_AXIMM_73_AWLEN(M_AXIMM_73_AWLEN),
        .M_AXIMM_73_AWSIZE(M_AXIMM_73_AWSIZE),
        .M_AXIMM_73_AWBURST(M_AXIMM_73_AWBURST),
        .M_AXIMM_73_AWLOCK(M_AXIMM_73_AWLOCK),
        .M_AXIMM_73_AWCACHE(M_AXIMM_73_AWCACHE),
        .M_AXIMM_73_AWPROT(M_AXIMM_73_AWPROT),
        .M_AXIMM_73_AWREGION(M_AXIMM_73_AWREGION),
        .M_AXIMM_73_AWQOS(M_AXIMM_73_AWQOS),
        .M_AXIMM_73_AWVALID(M_AXIMM_73_AWVALID),
        .M_AXIMM_73_AWREADY(M_AXIMM_73_AWREADY),
        .M_AXIMM_73_WDATA(M_AXIMM_73_WDATA),
        .M_AXIMM_73_WSTRB(M_AXIMM_73_WSTRB),
        .M_AXIMM_73_WLAST(M_AXIMM_73_WLAST),
        .M_AXIMM_73_WVALID(M_AXIMM_73_WVALID),
        .M_AXIMM_73_WREADY(M_AXIMM_73_WREADY),
        .M_AXIMM_73_BRESP(M_AXIMM_73_BRESP),
        .M_AXIMM_73_BVALID(M_AXIMM_73_BVALID),
        .M_AXIMM_73_BREADY(M_AXIMM_73_BREADY),
        .M_AXIMM_73_ARADDR(M_AXIMM_73_ARADDR),
        .M_AXIMM_73_ARLEN(M_AXIMM_73_ARLEN),
        .M_AXIMM_73_ARSIZE(M_AXIMM_73_ARSIZE),
        .M_AXIMM_73_ARBURST(M_AXIMM_73_ARBURST),
        .M_AXIMM_73_ARLOCK(M_AXIMM_73_ARLOCK),
        .M_AXIMM_73_ARCACHE(M_AXIMM_73_ARCACHE),
        .M_AXIMM_73_ARPROT(M_AXIMM_73_ARPROT),
        .M_AXIMM_73_ARREGION(M_AXIMM_73_ARREGION),
        .M_AXIMM_73_ARQOS(M_AXIMM_73_ARQOS),
        .M_AXIMM_73_ARVALID(M_AXIMM_73_ARVALID),
        .M_AXIMM_73_ARREADY(M_AXIMM_73_ARREADY),
        .M_AXIMM_73_RDATA(M_AXIMM_73_RDATA),
        .M_AXIMM_73_RRESP(M_AXIMM_73_RRESP),
        .M_AXIMM_73_RLAST(M_AXIMM_73_RLAST),
        .M_AXIMM_73_RVALID(M_AXIMM_73_RVALID),
        .M_AXIMM_73_RREADY(M_AXIMM_73_RREADY),
        .AP_AXIMM_74_AWADDR(AP_AXIMM_74_AWADDR),
        .AP_AXIMM_74_AWLEN(AP_AXIMM_74_AWLEN),
        .AP_AXIMM_74_AWSIZE(AP_AXIMM_74_AWSIZE),
        .AP_AXIMM_74_AWBURST(AP_AXIMM_74_AWBURST),
        .AP_AXIMM_74_AWLOCK(AP_AXIMM_74_AWLOCK),
        .AP_AXIMM_74_AWCACHE(AP_AXIMM_74_AWCACHE),
        .AP_AXIMM_74_AWPROT(AP_AXIMM_74_AWPROT),
        .AP_AXIMM_74_AWREGION(AP_AXIMM_74_AWREGION),
        .AP_AXIMM_74_AWQOS(AP_AXIMM_74_AWQOS),
        .AP_AXIMM_74_AWVALID(AP_AXIMM_74_AWVALID),
        .AP_AXIMM_74_AWREADY(AP_AXIMM_74_AWREADY),
        .AP_AXIMM_74_WDATA(AP_AXIMM_74_WDATA),
        .AP_AXIMM_74_WSTRB(AP_AXIMM_74_WSTRB),
        .AP_AXIMM_74_WLAST(AP_AXIMM_74_WLAST),
        .AP_AXIMM_74_WVALID(AP_AXIMM_74_WVALID),
        .AP_AXIMM_74_WREADY(AP_AXIMM_74_WREADY),
        .AP_AXIMM_74_BRESP(AP_AXIMM_74_BRESP),
        .AP_AXIMM_74_BVALID(AP_AXIMM_74_BVALID),
        .AP_AXIMM_74_BREADY(AP_AXIMM_74_BREADY),
        .AP_AXIMM_74_ARADDR(AP_AXIMM_74_ARADDR),
        .AP_AXIMM_74_ARLEN(AP_AXIMM_74_ARLEN),
        .AP_AXIMM_74_ARSIZE(AP_AXIMM_74_ARSIZE),
        .AP_AXIMM_74_ARBURST(AP_AXIMM_74_ARBURST),
        .AP_AXIMM_74_ARLOCK(AP_AXIMM_74_ARLOCK),
        .AP_AXIMM_74_ARCACHE(AP_AXIMM_74_ARCACHE),
        .AP_AXIMM_74_ARPROT(AP_AXIMM_74_ARPROT),
        .AP_AXIMM_74_ARREGION(AP_AXIMM_74_ARREGION),
        .AP_AXIMM_74_ARQOS(AP_AXIMM_74_ARQOS),
        .AP_AXIMM_74_ARVALID(AP_AXIMM_74_ARVALID),
        .AP_AXIMM_74_ARREADY(AP_AXIMM_74_ARREADY),
        .AP_AXIMM_74_RDATA(AP_AXIMM_74_RDATA),
        .AP_AXIMM_74_RRESP(AP_AXIMM_74_RRESP),
        .AP_AXIMM_74_RLAST(AP_AXIMM_74_RLAST),
        .AP_AXIMM_74_RVALID(AP_AXIMM_74_RVALID),
        .AP_AXIMM_74_RREADY(AP_AXIMM_74_RREADY),
        .M_AXIMM_74_AWADDR(M_AXIMM_74_AWADDR),
        .M_AXIMM_74_AWLEN(M_AXIMM_74_AWLEN),
        .M_AXIMM_74_AWSIZE(M_AXIMM_74_AWSIZE),
        .M_AXIMM_74_AWBURST(M_AXIMM_74_AWBURST),
        .M_AXIMM_74_AWLOCK(M_AXIMM_74_AWLOCK),
        .M_AXIMM_74_AWCACHE(M_AXIMM_74_AWCACHE),
        .M_AXIMM_74_AWPROT(M_AXIMM_74_AWPROT),
        .M_AXIMM_74_AWREGION(M_AXIMM_74_AWREGION),
        .M_AXIMM_74_AWQOS(M_AXIMM_74_AWQOS),
        .M_AXIMM_74_AWVALID(M_AXIMM_74_AWVALID),
        .M_AXIMM_74_AWREADY(M_AXIMM_74_AWREADY),
        .M_AXIMM_74_WDATA(M_AXIMM_74_WDATA),
        .M_AXIMM_74_WSTRB(M_AXIMM_74_WSTRB),
        .M_AXIMM_74_WLAST(M_AXIMM_74_WLAST),
        .M_AXIMM_74_WVALID(M_AXIMM_74_WVALID),
        .M_AXIMM_74_WREADY(M_AXIMM_74_WREADY),
        .M_AXIMM_74_BRESP(M_AXIMM_74_BRESP),
        .M_AXIMM_74_BVALID(M_AXIMM_74_BVALID),
        .M_AXIMM_74_BREADY(M_AXIMM_74_BREADY),
        .M_AXIMM_74_ARADDR(M_AXIMM_74_ARADDR),
        .M_AXIMM_74_ARLEN(M_AXIMM_74_ARLEN),
        .M_AXIMM_74_ARSIZE(M_AXIMM_74_ARSIZE),
        .M_AXIMM_74_ARBURST(M_AXIMM_74_ARBURST),
        .M_AXIMM_74_ARLOCK(M_AXIMM_74_ARLOCK),
        .M_AXIMM_74_ARCACHE(M_AXIMM_74_ARCACHE),
        .M_AXIMM_74_ARPROT(M_AXIMM_74_ARPROT),
        .M_AXIMM_74_ARREGION(M_AXIMM_74_ARREGION),
        .M_AXIMM_74_ARQOS(M_AXIMM_74_ARQOS),
        .M_AXIMM_74_ARVALID(M_AXIMM_74_ARVALID),
        .M_AXIMM_74_ARREADY(M_AXIMM_74_ARREADY),
        .M_AXIMM_74_RDATA(M_AXIMM_74_RDATA),
        .M_AXIMM_74_RRESP(M_AXIMM_74_RRESP),
        .M_AXIMM_74_RLAST(M_AXIMM_74_RLAST),
        .M_AXIMM_74_RVALID(M_AXIMM_74_RVALID),
        .M_AXIMM_74_RREADY(M_AXIMM_74_RREADY),
        .AP_AXIMM_75_AWADDR(AP_AXIMM_75_AWADDR),
        .AP_AXIMM_75_AWLEN(AP_AXIMM_75_AWLEN),
        .AP_AXIMM_75_AWSIZE(AP_AXIMM_75_AWSIZE),
        .AP_AXIMM_75_AWBURST(AP_AXIMM_75_AWBURST),
        .AP_AXIMM_75_AWLOCK(AP_AXIMM_75_AWLOCK),
        .AP_AXIMM_75_AWCACHE(AP_AXIMM_75_AWCACHE),
        .AP_AXIMM_75_AWPROT(AP_AXIMM_75_AWPROT),
        .AP_AXIMM_75_AWREGION(AP_AXIMM_75_AWREGION),
        .AP_AXIMM_75_AWQOS(AP_AXIMM_75_AWQOS),
        .AP_AXIMM_75_AWVALID(AP_AXIMM_75_AWVALID),
        .AP_AXIMM_75_AWREADY(AP_AXIMM_75_AWREADY),
        .AP_AXIMM_75_WDATA(AP_AXIMM_75_WDATA),
        .AP_AXIMM_75_WSTRB(AP_AXIMM_75_WSTRB),
        .AP_AXIMM_75_WLAST(AP_AXIMM_75_WLAST),
        .AP_AXIMM_75_WVALID(AP_AXIMM_75_WVALID),
        .AP_AXIMM_75_WREADY(AP_AXIMM_75_WREADY),
        .AP_AXIMM_75_BRESP(AP_AXIMM_75_BRESP),
        .AP_AXIMM_75_BVALID(AP_AXIMM_75_BVALID),
        .AP_AXIMM_75_BREADY(AP_AXIMM_75_BREADY),
        .AP_AXIMM_75_ARADDR(AP_AXIMM_75_ARADDR),
        .AP_AXIMM_75_ARLEN(AP_AXIMM_75_ARLEN),
        .AP_AXIMM_75_ARSIZE(AP_AXIMM_75_ARSIZE),
        .AP_AXIMM_75_ARBURST(AP_AXIMM_75_ARBURST),
        .AP_AXIMM_75_ARLOCK(AP_AXIMM_75_ARLOCK),
        .AP_AXIMM_75_ARCACHE(AP_AXIMM_75_ARCACHE),
        .AP_AXIMM_75_ARPROT(AP_AXIMM_75_ARPROT),
        .AP_AXIMM_75_ARREGION(AP_AXIMM_75_ARREGION),
        .AP_AXIMM_75_ARQOS(AP_AXIMM_75_ARQOS),
        .AP_AXIMM_75_ARVALID(AP_AXIMM_75_ARVALID),
        .AP_AXIMM_75_ARREADY(AP_AXIMM_75_ARREADY),
        .AP_AXIMM_75_RDATA(AP_AXIMM_75_RDATA),
        .AP_AXIMM_75_RRESP(AP_AXIMM_75_RRESP),
        .AP_AXIMM_75_RLAST(AP_AXIMM_75_RLAST),
        .AP_AXIMM_75_RVALID(AP_AXIMM_75_RVALID),
        .AP_AXIMM_75_RREADY(AP_AXIMM_75_RREADY),
        .M_AXIMM_75_AWADDR(M_AXIMM_75_AWADDR),
        .M_AXIMM_75_AWLEN(M_AXIMM_75_AWLEN),
        .M_AXIMM_75_AWSIZE(M_AXIMM_75_AWSIZE),
        .M_AXIMM_75_AWBURST(M_AXIMM_75_AWBURST),
        .M_AXIMM_75_AWLOCK(M_AXIMM_75_AWLOCK),
        .M_AXIMM_75_AWCACHE(M_AXIMM_75_AWCACHE),
        .M_AXIMM_75_AWPROT(M_AXIMM_75_AWPROT),
        .M_AXIMM_75_AWREGION(M_AXIMM_75_AWREGION),
        .M_AXIMM_75_AWQOS(M_AXIMM_75_AWQOS),
        .M_AXIMM_75_AWVALID(M_AXIMM_75_AWVALID),
        .M_AXIMM_75_AWREADY(M_AXIMM_75_AWREADY),
        .M_AXIMM_75_WDATA(M_AXIMM_75_WDATA),
        .M_AXIMM_75_WSTRB(M_AXIMM_75_WSTRB),
        .M_AXIMM_75_WLAST(M_AXIMM_75_WLAST),
        .M_AXIMM_75_WVALID(M_AXIMM_75_WVALID),
        .M_AXIMM_75_WREADY(M_AXIMM_75_WREADY),
        .M_AXIMM_75_BRESP(M_AXIMM_75_BRESP),
        .M_AXIMM_75_BVALID(M_AXIMM_75_BVALID),
        .M_AXIMM_75_BREADY(M_AXIMM_75_BREADY),
        .M_AXIMM_75_ARADDR(M_AXIMM_75_ARADDR),
        .M_AXIMM_75_ARLEN(M_AXIMM_75_ARLEN),
        .M_AXIMM_75_ARSIZE(M_AXIMM_75_ARSIZE),
        .M_AXIMM_75_ARBURST(M_AXIMM_75_ARBURST),
        .M_AXIMM_75_ARLOCK(M_AXIMM_75_ARLOCK),
        .M_AXIMM_75_ARCACHE(M_AXIMM_75_ARCACHE),
        .M_AXIMM_75_ARPROT(M_AXIMM_75_ARPROT),
        .M_AXIMM_75_ARREGION(M_AXIMM_75_ARREGION),
        .M_AXIMM_75_ARQOS(M_AXIMM_75_ARQOS),
        .M_AXIMM_75_ARVALID(M_AXIMM_75_ARVALID),
        .M_AXIMM_75_ARREADY(M_AXIMM_75_ARREADY),
        .M_AXIMM_75_RDATA(M_AXIMM_75_RDATA),
        .M_AXIMM_75_RRESP(M_AXIMM_75_RRESP),
        .M_AXIMM_75_RLAST(M_AXIMM_75_RLAST),
        .M_AXIMM_75_RVALID(M_AXIMM_75_RVALID),
        .M_AXIMM_75_RREADY(M_AXIMM_75_RREADY),
        .AP_AXIMM_76_AWADDR(AP_AXIMM_76_AWADDR),
        .AP_AXIMM_76_AWLEN(AP_AXIMM_76_AWLEN),
        .AP_AXIMM_76_AWSIZE(AP_AXIMM_76_AWSIZE),
        .AP_AXIMM_76_AWBURST(AP_AXIMM_76_AWBURST),
        .AP_AXIMM_76_AWLOCK(AP_AXIMM_76_AWLOCK),
        .AP_AXIMM_76_AWCACHE(AP_AXIMM_76_AWCACHE),
        .AP_AXIMM_76_AWPROT(AP_AXIMM_76_AWPROT),
        .AP_AXIMM_76_AWREGION(AP_AXIMM_76_AWREGION),
        .AP_AXIMM_76_AWQOS(AP_AXIMM_76_AWQOS),
        .AP_AXIMM_76_AWVALID(AP_AXIMM_76_AWVALID),
        .AP_AXIMM_76_AWREADY(AP_AXIMM_76_AWREADY),
        .AP_AXIMM_76_WDATA(AP_AXIMM_76_WDATA),
        .AP_AXIMM_76_WSTRB(AP_AXIMM_76_WSTRB),
        .AP_AXIMM_76_WLAST(AP_AXIMM_76_WLAST),
        .AP_AXIMM_76_WVALID(AP_AXIMM_76_WVALID),
        .AP_AXIMM_76_WREADY(AP_AXIMM_76_WREADY),
        .AP_AXIMM_76_BRESP(AP_AXIMM_76_BRESP),
        .AP_AXIMM_76_BVALID(AP_AXIMM_76_BVALID),
        .AP_AXIMM_76_BREADY(AP_AXIMM_76_BREADY),
        .AP_AXIMM_76_ARADDR(AP_AXIMM_76_ARADDR),
        .AP_AXIMM_76_ARLEN(AP_AXIMM_76_ARLEN),
        .AP_AXIMM_76_ARSIZE(AP_AXIMM_76_ARSIZE),
        .AP_AXIMM_76_ARBURST(AP_AXIMM_76_ARBURST),
        .AP_AXIMM_76_ARLOCK(AP_AXIMM_76_ARLOCK),
        .AP_AXIMM_76_ARCACHE(AP_AXIMM_76_ARCACHE),
        .AP_AXIMM_76_ARPROT(AP_AXIMM_76_ARPROT),
        .AP_AXIMM_76_ARREGION(AP_AXIMM_76_ARREGION),
        .AP_AXIMM_76_ARQOS(AP_AXIMM_76_ARQOS),
        .AP_AXIMM_76_ARVALID(AP_AXIMM_76_ARVALID),
        .AP_AXIMM_76_ARREADY(AP_AXIMM_76_ARREADY),
        .AP_AXIMM_76_RDATA(AP_AXIMM_76_RDATA),
        .AP_AXIMM_76_RRESP(AP_AXIMM_76_RRESP),
        .AP_AXIMM_76_RLAST(AP_AXIMM_76_RLAST),
        .AP_AXIMM_76_RVALID(AP_AXIMM_76_RVALID),
        .AP_AXIMM_76_RREADY(AP_AXIMM_76_RREADY),
        .M_AXIMM_76_AWADDR(M_AXIMM_76_AWADDR),
        .M_AXIMM_76_AWLEN(M_AXIMM_76_AWLEN),
        .M_AXIMM_76_AWSIZE(M_AXIMM_76_AWSIZE),
        .M_AXIMM_76_AWBURST(M_AXIMM_76_AWBURST),
        .M_AXIMM_76_AWLOCK(M_AXIMM_76_AWLOCK),
        .M_AXIMM_76_AWCACHE(M_AXIMM_76_AWCACHE),
        .M_AXIMM_76_AWPROT(M_AXIMM_76_AWPROT),
        .M_AXIMM_76_AWREGION(M_AXIMM_76_AWREGION),
        .M_AXIMM_76_AWQOS(M_AXIMM_76_AWQOS),
        .M_AXIMM_76_AWVALID(M_AXIMM_76_AWVALID),
        .M_AXIMM_76_AWREADY(M_AXIMM_76_AWREADY),
        .M_AXIMM_76_WDATA(M_AXIMM_76_WDATA),
        .M_AXIMM_76_WSTRB(M_AXIMM_76_WSTRB),
        .M_AXIMM_76_WLAST(M_AXIMM_76_WLAST),
        .M_AXIMM_76_WVALID(M_AXIMM_76_WVALID),
        .M_AXIMM_76_WREADY(M_AXIMM_76_WREADY),
        .M_AXIMM_76_BRESP(M_AXIMM_76_BRESP),
        .M_AXIMM_76_BVALID(M_AXIMM_76_BVALID),
        .M_AXIMM_76_BREADY(M_AXIMM_76_BREADY),
        .M_AXIMM_76_ARADDR(M_AXIMM_76_ARADDR),
        .M_AXIMM_76_ARLEN(M_AXIMM_76_ARLEN),
        .M_AXIMM_76_ARSIZE(M_AXIMM_76_ARSIZE),
        .M_AXIMM_76_ARBURST(M_AXIMM_76_ARBURST),
        .M_AXIMM_76_ARLOCK(M_AXIMM_76_ARLOCK),
        .M_AXIMM_76_ARCACHE(M_AXIMM_76_ARCACHE),
        .M_AXIMM_76_ARPROT(M_AXIMM_76_ARPROT),
        .M_AXIMM_76_ARREGION(M_AXIMM_76_ARREGION),
        .M_AXIMM_76_ARQOS(M_AXIMM_76_ARQOS),
        .M_AXIMM_76_ARVALID(M_AXIMM_76_ARVALID),
        .M_AXIMM_76_ARREADY(M_AXIMM_76_ARREADY),
        .M_AXIMM_76_RDATA(M_AXIMM_76_RDATA),
        .M_AXIMM_76_RRESP(M_AXIMM_76_RRESP),
        .M_AXIMM_76_RLAST(M_AXIMM_76_RLAST),
        .M_AXIMM_76_RVALID(M_AXIMM_76_RVALID),
        .M_AXIMM_76_RREADY(M_AXIMM_76_RREADY),
        .AP_AXIMM_77_AWADDR(AP_AXIMM_77_AWADDR),
        .AP_AXIMM_77_AWLEN(AP_AXIMM_77_AWLEN),
        .AP_AXIMM_77_AWSIZE(AP_AXIMM_77_AWSIZE),
        .AP_AXIMM_77_AWBURST(AP_AXIMM_77_AWBURST),
        .AP_AXIMM_77_AWLOCK(AP_AXIMM_77_AWLOCK),
        .AP_AXIMM_77_AWCACHE(AP_AXIMM_77_AWCACHE),
        .AP_AXIMM_77_AWPROT(AP_AXIMM_77_AWPROT),
        .AP_AXIMM_77_AWREGION(AP_AXIMM_77_AWREGION),
        .AP_AXIMM_77_AWQOS(AP_AXIMM_77_AWQOS),
        .AP_AXIMM_77_AWVALID(AP_AXIMM_77_AWVALID),
        .AP_AXIMM_77_AWREADY(AP_AXIMM_77_AWREADY),
        .AP_AXIMM_77_WDATA(AP_AXIMM_77_WDATA),
        .AP_AXIMM_77_WSTRB(AP_AXIMM_77_WSTRB),
        .AP_AXIMM_77_WLAST(AP_AXIMM_77_WLAST),
        .AP_AXIMM_77_WVALID(AP_AXIMM_77_WVALID),
        .AP_AXIMM_77_WREADY(AP_AXIMM_77_WREADY),
        .AP_AXIMM_77_BRESP(AP_AXIMM_77_BRESP),
        .AP_AXIMM_77_BVALID(AP_AXIMM_77_BVALID),
        .AP_AXIMM_77_BREADY(AP_AXIMM_77_BREADY),
        .AP_AXIMM_77_ARADDR(AP_AXIMM_77_ARADDR),
        .AP_AXIMM_77_ARLEN(AP_AXIMM_77_ARLEN),
        .AP_AXIMM_77_ARSIZE(AP_AXIMM_77_ARSIZE),
        .AP_AXIMM_77_ARBURST(AP_AXIMM_77_ARBURST),
        .AP_AXIMM_77_ARLOCK(AP_AXIMM_77_ARLOCK),
        .AP_AXIMM_77_ARCACHE(AP_AXIMM_77_ARCACHE),
        .AP_AXIMM_77_ARPROT(AP_AXIMM_77_ARPROT),
        .AP_AXIMM_77_ARREGION(AP_AXIMM_77_ARREGION),
        .AP_AXIMM_77_ARQOS(AP_AXIMM_77_ARQOS),
        .AP_AXIMM_77_ARVALID(AP_AXIMM_77_ARVALID),
        .AP_AXIMM_77_ARREADY(AP_AXIMM_77_ARREADY),
        .AP_AXIMM_77_RDATA(AP_AXIMM_77_RDATA),
        .AP_AXIMM_77_RRESP(AP_AXIMM_77_RRESP),
        .AP_AXIMM_77_RLAST(AP_AXIMM_77_RLAST),
        .AP_AXIMM_77_RVALID(AP_AXIMM_77_RVALID),
        .AP_AXIMM_77_RREADY(AP_AXIMM_77_RREADY),
        .M_AXIMM_77_AWADDR(M_AXIMM_77_AWADDR),
        .M_AXIMM_77_AWLEN(M_AXIMM_77_AWLEN),
        .M_AXIMM_77_AWSIZE(M_AXIMM_77_AWSIZE),
        .M_AXIMM_77_AWBURST(M_AXIMM_77_AWBURST),
        .M_AXIMM_77_AWLOCK(M_AXIMM_77_AWLOCK),
        .M_AXIMM_77_AWCACHE(M_AXIMM_77_AWCACHE),
        .M_AXIMM_77_AWPROT(M_AXIMM_77_AWPROT),
        .M_AXIMM_77_AWREGION(M_AXIMM_77_AWREGION),
        .M_AXIMM_77_AWQOS(M_AXIMM_77_AWQOS),
        .M_AXIMM_77_AWVALID(M_AXIMM_77_AWVALID),
        .M_AXIMM_77_AWREADY(M_AXIMM_77_AWREADY),
        .M_AXIMM_77_WDATA(M_AXIMM_77_WDATA),
        .M_AXIMM_77_WSTRB(M_AXIMM_77_WSTRB),
        .M_AXIMM_77_WLAST(M_AXIMM_77_WLAST),
        .M_AXIMM_77_WVALID(M_AXIMM_77_WVALID),
        .M_AXIMM_77_WREADY(M_AXIMM_77_WREADY),
        .M_AXIMM_77_BRESP(M_AXIMM_77_BRESP),
        .M_AXIMM_77_BVALID(M_AXIMM_77_BVALID),
        .M_AXIMM_77_BREADY(M_AXIMM_77_BREADY),
        .M_AXIMM_77_ARADDR(M_AXIMM_77_ARADDR),
        .M_AXIMM_77_ARLEN(M_AXIMM_77_ARLEN),
        .M_AXIMM_77_ARSIZE(M_AXIMM_77_ARSIZE),
        .M_AXIMM_77_ARBURST(M_AXIMM_77_ARBURST),
        .M_AXIMM_77_ARLOCK(M_AXIMM_77_ARLOCK),
        .M_AXIMM_77_ARCACHE(M_AXIMM_77_ARCACHE),
        .M_AXIMM_77_ARPROT(M_AXIMM_77_ARPROT),
        .M_AXIMM_77_ARREGION(M_AXIMM_77_ARREGION),
        .M_AXIMM_77_ARQOS(M_AXIMM_77_ARQOS),
        .M_AXIMM_77_ARVALID(M_AXIMM_77_ARVALID),
        .M_AXIMM_77_ARREADY(M_AXIMM_77_ARREADY),
        .M_AXIMM_77_RDATA(M_AXIMM_77_RDATA),
        .M_AXIMM_77_RRESP(M_AXIMM_77_RRESP),
        .M_AXIMM_77_RLAST(M_AXIMM_77_RLAST),
        .M_AXIMM_77_RVALID(M_AXIMM_77_RVALID),
        .M_AXIMM_77_RREADY(M_AXIMM_77_RREADY),
        .AP_AXIMM_78_AWADDR(AP_AXIMM_78_AWADDR),
        .AP_AXIMM_78_AWLEN(AP_AXIMM_78_AWLEN),
        .AP_AXIMM_78_AWSIZE(AP_AXIMM_78_AWSIZE),
        .AP_AXIMM_78_AWBURST(AP_AXIMM_78_AWBURST),
        .AP_AXIMM_78_AWLOCK(AP_AXIMM_78_AWLOCK),
        .AP_AXIMM_78_AWCACHE(AP_AXIMM_78_AWCACHE),
        .AP_AXIMM_78_AWPROT(AP_AXIMM_78_AWPROT),
        .AP_AXIMM_78_AWREGION(AP_AXIMM_78_AWREGION),
        .AP_AXIMM_78_AWQOS(AP_AXIMM_78_AWQOS),
        .AP_AXIMM_78_AWVALID(AP_AXIMM_78_AWVALID),
        .AP_AXIMM_78_AWREADY(AP_AXIMM_78_AWREADY),
        .AP_AXIMM_78_WDATA(AP_AXIMM_78_WDATA),
        .AP_AXIMM_78_WSTRB(AP_AXIMM_78_WSTRB),
        .AP_AXIMM_78_WLAST(AP_AXIMM_78_WLAST),
        .AP_AXIMM_78_WVALID(AP_AXIMM_78_WVALID),
        .AP_AXIMM_78_WREADY(AP_AXIMM_78_WREADY),
        .AP_AXIMM_78_BRESP(AP_AXIMM_78_BRESP),
        .AP_AXIMM_78_BVALID(AP_AXIMM_78_BVALID),
        .AP_AXIMM_78_BREADY(AP_AXIMM_78_BREADY),
        .AP_AXIMM_78_ARADDR(AP_AXIMM_78_ARADDR),
        .AP_AXIMM_78_ARLEN(AP_AXIMM_78_ARLEN),
        .AP_AXIMM_78_ARSIZE(AP_AXIMM_78_ARSIZE),
        .AP_AXIMM_78_ARBURST(AP_AXIMM_78_ARBURST),
        .AP_AXIMM_78_ARLOCK(AP_AXIMM_78_ARLOCK),
        .AP_AXIMM_78_ARCACHE(AP_AXIMM_78_ARCACHE),
        .AP_AXIMM_78_ARPROT(AP_AXIMM_78_ARPROT),
        .AP_AXIMM_78_ARREGION(AP_AXIMM_78_ARREGION),
        .AP_AXIMM_78_ARQOS(AP_AXIMM_78_ARQOS),
        .AP_AXIMM_78_ARVALID(AP_AXIMM_78_ARVALID),
        .AP_AXIMM_78_ARREADY(AP_AXIMM_78_ARREADY),
        .AP_AXIMM_78_RDATA(AP_AXIMM_78_RDATA),
        .AP_AXIMM_78_RRESP(AP_AXIMM_78_RRESP),
        .AP_AXIMM_78_RLAST(AP_AXIMM_78_RLAST),
        .AP_AXIMM_78_RVALID(AP_AXIMM_78_RVALID),
        .AP_AXIMM_78_RREADY(AP_AXIMM_78_RREADY),
        .M_AXIMM_78_AWADDR(M_AXIMM_78_AWADDR),
        .M_AXIMM_78_AWLEN(M_AXIMM_78_AWLEN),
        .M_AXIMM_78_AWSIZE(M_AXIMM_78_AWSIZE),
        .M_AXIMM_78_AWBURST(M_AXIMM_78_AWBURST),
        .M_AXIMM_78_AWLOCK(M_AXIMM_78_AWLOCK),
        .M_AXIMM_78_AWCACHE(M_AXIMM_78_AWCACHE),
        .M_AXIMM_78_AWPROT(M_AXIMM_78_AWPROT),
        .M_AXIMM_78_AWREGION(M_AXIMM_78_AWREGION),
        .M_AXIMM_78_AWQOS(M_AXIMM_78_AWQOS),
        .M_AXIMM_78_AWVALID(M_AXIMM_78_AWVALID),
        .M_AXIMM_78_AWREADY(M_AXIMM_78_AWREADY),
        .M_AXIMM_78_WDATA(M_AXIMM_78_WDATA),
        .M_AXIMM_78_WSTRB(M_AXIMM_78_WSTRB),
        .M_AXIMM_78_WLAST(M_AXIMM_78_WLAST),
        .M_AXIMM_78_WVALID(M_AXIMM_78_WVALID),
        .M_AXIMM_78_WREADY(M_AXIMM_78_WREADY),
        .M_AXIMM_78_BRESP(M_AXIMM_78_BRESP),
        .M_AXIMM_78_BVALID(M_AXIMM_78_BVALID),
        .M_AXIMM_78_BREADY(M_AXIMM_78_BREADY),
        .M_AXIMM_78_ARADDR(M_AXIMM_78_ARADDR),
        .M_AXIMM_78_ARLEN(M_AXIMM_78_ARLEN),
        .M_AXIMM_78_ARSIZE(M_AXIMM_78_ARSIZE),
        .M_AXIMM_78_ARBURST(M_AXIMM_78_ARBURST),
        .M_AXIMM_78_ARLOCK(M_AXIMM_78_ARLOCK),
        .M_AXIMM_78_ARCACHE(M_AXIMM_78_ARCACHE),
        .M_AXIMM_78_ARPROT(M_AXIMM_78_ARPROT),
        .M_AXIMM_78_ARREGION(M_AXIMM_78_ARREGION),
        .M_AXIMM_78_ARQOS(M_AXIMM_78_ARQOS),
        .M_AXIMM_78_ARVALID(M_AXIMM_78_ARVALID),
        .M_AXIMM_78_ARREADY(M_AXIMM_78_ARREADY),
        .M_AXIMM_78_RDATA(M_AXIMM_78_RDATA),
        .M_AXIMM_78_RRESP(M_AXIMM_78_RRESP),
        .M_AXIMM_78_RLAST(M_AXIMM_78_RLAST),
        .M_AXIMM_78_RVALID(M_AXIMM_78_RVALID),
        .M_AXIMM_78_RREADY(M_AXIMM_78_RREADY),
        .AP_AXIMM_79_AWADDR(AP_AXIMM_79_AWADDR),
        .AP_AXIMM_79_AWLEN(AP_AXIMM_79_AWLEN),
        .AP_AXIMM_79_AWSIZE(AP_AXIMM_79_AWSIZE),
        .AP_AXIMM_79_AWBURST(AP_AXIMM_79_AWBURST),
        .AP_AXIMM_79_AWLOCK(AP_AXIMM_79_AWLOCK),
        .AP_AXIMM_79_AWCACHE(AP_AXIMM_79_AWCACHE),
        .AP_AXIMM_79_AWPROT(AP_AXIMM_79_AWPROT),
        .AP_AXIMM_79_AWREGION(AP_AXIMM_79_AWREGION),
        .AP_AXIMM_79_AWQOS(AP_AXIMM_79_AWQOS),
        .AP_AXIMM_79_AWVALID(AP_AXIMM_79_AWVALID),
        .AP_AXIMM_79_AWREADY(AP_AXIMM_79_AWREADY),
        .AP_AXIMM_79_WDATA(AP_AXIMM_79_WDATA),
        .AP_AXIMM_79_WSTRB(AP_AXIMM_79_WSTRB),
        .AP_AXIMM_79_WLAST(AP_AXIMM_79_WLAST),
        .AP_AXIMM_79_WVALID(AP_AXIMM_79_WVALID),
        .AP_AXIMM_79_WREADY(AP_AXIMM_79_WREADY),
        .AP_AXIMM_79_BRESP(AP_AXIMM_79_BRESP),
        .AP_AXIMM_79_BVALID(AP_AXIMM_79_BVALID),
        .AP_AXIMM_79_BREADY(AP_AXIMM_79_BREADY),
        .AP_AXIMM_79_ARADDR(AP_AXIMM_79_ARADDR),
        .AP_AXIMM_79_ARLEN(AP_AXIMM_79_ARLEN),
        .AP_AXIMM_79_ARSIZE(AP_AXIMM_79_ARSIZE),
        .AP_AXIMM_79_ARBURST(AP_AXIMM_79_ARBURST),
        .AP_AXIMM_79_ARLOCK(AP_AXIMM_79_ARLOCK),
        .AP_AXIMM_79_ARCACHE(AP_AXIMM_79_ARCACHE),
        .AP_AXIMM_79_ARPROT(AP_AXIMM_79_ARPROT),
        .AP_AXIMM_79_ARREGION(AP_AXIMM_79_ARREGION),
        .AP_AXIMM_79_ARQOS(AP_AXIMM_79_ARQOS),
        .AP_AXIMM_79_ARVALID(AP_AXIMM_79_ARVALID),
        .AP_AXIMM_79_ARREADY(AP_AXIMM_79_ARREADY),
        .AP_AXIMM_79_RDATA(AP_AXIMM_79_RDATA),
        .AP_AXIMM_79_RRESP(AP_AXIMM_79_RRESP),
        .AP_AXIMM_79_RLAST(AP_AXIMM_79_RLAST),
        .AP_AXIMM_79_RVALID(AP_AXIMM_79_RVALID),
        .AP_AXIMM_79_RREADY(AP_AXIMM_79_RREADY),
        .M_AXIMM_79_AWADDR(M_AXIMM_79_AWADDR),
        .M_AXIMM_79_AWLEN(M_AXIMM_79_AWLEN),
        .M_AXIMM_79_AWSIZE(M_AXIMM_79_AWSIZE),
        .M_AXIMM_79_AWBURST(M_AXIMM_79_AWBURST),
        .M_AXIMM_79_AWLOCK(M_AXIMM_79_AWLOCK),
        .M_AXIMM_79_AWCACHE(M_AXIMM_79_AWCACHE),
        .M_AXIMM_79_AWPROT(M_AXIMM_79_AWPROT),
        .M_AXIMM_79_AWREGION(M_AXIMM_79_AWREGION),
        .M_AXIMM_79_AWQOS(M_AXIMM_79_AWQOS),
        .M_AXIMM_79_AWVALID(M_AXIMM_79_AWVALID),
        .M_AXIMM_79_AWREADY(M_AXIMM_79_AWREADY),
        .M_AXIMM_79_WDATA(M_AXIMM_79_WDATA),
        .M_AXIMM_79_WSTRB(M_AXIMM_79_WSTRB),
        .M_AXIMM_79_WLAST(M_AXIMM_79_WLAST),
        .M_AXIMM_79_WVALID(M_AXIMM_79_WVALID),
        .M_AXIMM_79_WREADY(M_AXIMM_79_WREADY),
        .M_AXIMM_79_BRESP(M_AXIMM_79_BRESP),
        .M_AXIMM_79_BVALID(M_AXIMM_79_BVALID),
        .M_AXIMM_79_BREADY(M_AXIMM_79_BREADY),
        .M_AXIMM_79_ARADDR(M_AXIMM_79_ARADDR),
        .M_AXIMM_79_ARLEN(M_AXIMM_79_ARLEN),
        .M_AXIMM_79_ARSIZE(M_AXIMM_79_ARSIZE),
        .M_AXIMM_79_ARBURST(M_AXIMM_79_ARBURST),
        .M_AXIMM_79_ARLOCK(M_AXIMM_79_ARLOCK),
        .M_AXIMM_79_ARCACHE(M_AXIMM_79_ARCACHE),
        .M_AXIMM_79_ARPROT(M_AXIMM_79_ARPROT),
        .M_AXIMM_79_ARREGION(M_AXIMM_79_ARREGION),
        .M_AXIMM_79_ARQOS(M_AXIMM_79_ARQOS),
        .M_AXIMM_79_ARVALID(M_AXIMM_79_ARVALID),
        .M_AXIMM_79_ARREADY(M_AXIMM_79_ARREADY),
        .M_AXIMM_79_RDATA(M_AXIMM_79_RDATA),
        .M_AXIMM_79_RRESP(M_AXIMM_79_RRESP),
        .M_AXIMM_79_RLAST(M_AXIMM_79_RLAST),
        .M_AXIMM_79_RVALID(M_AXIMM_79_RVALID),
        .M_AXIMM_79_RREADY(M_AXIMM_79_RREADY),
        .AP_AXIMM_80_AWADDR(AP_AXIMM_80_AWADDR),
        .AP_AXIMM_80_AWLEN(AP_AXIMM_80_AWLEN),
        .AP_AXIMM_80_AWSIZE(AP_AXIMM_80_AWSIZE),
        .AP_AXIMM_80_AWBURST(AP_AXIMM_80_AWBURST),
        .AP_AXIMM_80_AWLOCK(AP_AXIMM_80_AWLOCK),
        .AP_AXIMM_80_AWCACHE(AP_AXIMM_80_AWCACHE),
        .AP_AXIMM_80_AWPROT(AP_AXIMM_80_AWPROT),
        .AP_AXIMM_80_AWREGION(AP_AXIMM_80_AWREGION),
        .AP_AXIMM_80_AWQOS(AP_AXIMM_80_AWQOS),
        .AP_AXIMM_80_AWVALID(AP_AXIMM_80_AWVALID),
        .AP_AXIMM_80_AWREADY(AP_AXIMM_80_AWREADY),
        .AP_AXIMM_80_WDATA(AP_AXIMM_80_WDATA),
        .AP_AXIMM_80_WSTRB(AP_AXIMM_80_WSTRB),
        .AP_AXIMM_80_WLAST(AP_AXIMM_80_WLAST),
        .AP_AXIMM_80_WVALID(AP_AXIMM_80_WVALID),
        .AP_AXIMM_80_WREADY(AP_AXIMM_80_WREADY),
        .AP_AXIMM_80_BRESP(AP_AXIMM_80_BRESP),
        .AP_AXIMM_80_BVALID(AP_AXIMM_80_BVALID),
        .AP_AXIMM_80_BREADY(AP_AXIMM_80_BREADY),
        .AP_AXIMM_80_ARADDR(AP_AXIMM_80_ARADDR),
        .AP_AXIMM_80_ARLEN(AP_AXIMM_80_ARLEN),
        .AP_AXIMM_80_ARSIZE(AP_AXIMM_80_ARSIZE),
        .AP_AXIMM_80_ARBURST(AP_AXIMM_80_ARBURST),
        .AP_AXIMM_80_ARLOCK(AP_AXIMM_80_ARLOCK),
        .AP_AXIMM_80_ARCACHE(AP_AXIMM_80_ARCACHE),
        .AP_AXIMM_80_ARPROT(AP_AXIMM_80_ARPROT),
        .AP_AXIMM_80_ARREGION(AP_AXIMM_80_ARREGION),
        .AP_AXIMM_80_ARQOS(AP_AXIMM_80_ARQOS),
        .AP_AXIMM_80_ARVALID(AP_AXIMM_80_ARVALID),
        .AP_AXIMM_80_ARREADY(AP_AXIMM_80_ARREADY),
        .AP_AXIMM_80_RDATA(AP_AXIMM_80_RDATA),
        .AP_AXIMM_80_RRESP(AP_AXIMM_80_RRESP),
        .AP_AXIMM_80_RLAST(AP_AXIMM_80_RLAST),
        .AP_AXIMM_80_RVALID(AP_AXIMM_80_RVALID),
        .AP_AXIMM_80_RREADY(AP_AXIMM_80_RREADY),
        .M_AXIMM_80_AWADDR(M_AXIMM_80_AWADDR),
        .M_AXIMM_80_AWLEN(M_AXIMM_80_AWLEN),
        .M_AXIMM_80_AWSIZE(M_AXIMM_80_AWSIZE),
        .M_AXIMM_80_AWBURST(M_AXIMM_80_AWBURST),
        .M_AXIMM_80_AWLOCK(M_AXIMM_80_AWLOCK),
        .M_AXIMM_80_AWCACHE(M_AXIMM_80_AWCACHE),
        .M_AXIMM_80_AWPROT(M_AXIMM_80_AWPROT),
        .M_AXIMM_80_AWREGION(M_AXIMM_80_AWREGION),
        .M_AXIMM_80_AWQOS(M_AXIMM_80_AWQOS),
        .M_AXIMM_80_AWVALID(M_AXIMM_80_AWVALID),
        .M_AXIMM_80_AWREADY(M_AXIMM_80_AWREADY),
        .M_AXIMM_80_WDATA(M_AXIMM_80_WDATA),
        .M_AXIMM_80_WSTRB(M_AXIMM_80_WSTRB),
        .M_AXIMM_80_WLAST(M_AXIMM_80_WLAST),
        .M_AXIMM_80_WVALID(M_AXIMM_80_WVALID),
        .M_AXIMM_80_WREADY(M_AXIMM_80_WREADY),
        .M_AXIMM_80_BRESP(M_AXIMM_80_BRESP),
        .M_AXIMM_80_BVALID(M_AXIMM_80_BVALID),
        .M_AXIMM_80_BREADY(M_AXIMM_80_BREADY),
        .M_AXIMM_80_ARADDR(M_AXIMM_80_ARADDR),
        .M_AXIMM_80_ARLEN(M_AXIMM_80_ARLEN),
        .M_AXIMM_80_ARSIZE(M_AXIMM_80_ARSIZE),
        .M_AXIMM_80_ARBURST(M_AXIMM_80_ARBURST),
        .M_AXIMM_80_ARLOCK(M_AXIMM_80_ARLOCK),
        .M_AXIMM_80_ARCACHE(M_AXIMM_80_ARCACHE),
        .M_AXIMM_80_ARPROT(M_AXIMM_80_ARPROT),
        .M_AXIMM_80_ARREGION(M_AXIMM_80_ARREGION),
        .M_AXIMM_80_ARQOS(M_AXIMM_80_ARQOS),
        .M_AXIMM_80_ARVALID(M_AXIMM_80_ARVALID),
        .M_AXIMM_80_ARREADY(M_AXIMM_80_ARREADY),
        .M_AXIMM_80_RDATA(M_AXIMM_80_RDATA),
        .M_AXIMM_80_RRESP(M_AXIMM_80_RRESP),
        .M_AXIMM_80_RLAST(M_AXIMM_80_RLAST),
        .M_AXIMM_80_RVALID(M_AXIMM_80_RVALID),
        .M_AXIMM_80_RREADY(M_AXIMM_80_RREADY),
        .AP_AXIMM_81_AWADDR(AP_AXIMM_81_AWADDR),
        .AP_AXIMM_81_AWLEN(AP_AXIMM_81_AWLEN),
        .AP_AXIMM_81_AWSIZE(AP_AXIMM_81_AWSIZE),
        .AP_AXIMM_81_AWBURST(AP_AXIMM_81_AWBURST),
        .AP_AXIMM_81_AWLOCK(AP_AXIMM_81_AWLOCK),
        .AP_AXIMM_81_AWCACHE(AP_AXIMM_81_AWCACHE),
        .AP_AXIMM_81_AWPROT(AP_AXIMM_81_AWPROT),
        .AP_AXIMM_81_AWREGION(AP_AXIMM_81_AWREGION),
        .AP_AXIMM_81_AWQOS(AP_AXIMM_81_AWQOS),
        .AP_AXIMM_81_AWVALID(AP_AXIMM_81_AWVALID),
        .AP_AXIMM_81_AWREADY(AP_AXIMM_81_AWREADY),
        .AP_AXIMM_81_WDATA(AP_AXIMM_81_WDATA),
        .AP_AXIMM_81_WSTRB(AP_AXIMM_81_WSTRB),
        .AP_AXIMM_81_WLAST(AP_AXIMM_81_WLAST),
        .AP_AXIMM_81_WVALID(AP_AXIMM_81_WVALID),
        .AP_AXIMM_81_WREADY(AP_AXIMM_81_WREADY),
        .AP_AXIMM_81_BRESP(AP_AXIMM_81_BRESP),
        .AP_AXIMM_81_BVALID(AP_AXIMM_81_BVALID),
        .AP_AXIMM_81_BREADY(AP_AXIMM_81_BREADY),
        .AP_AXIMM_81_ARADDR(AP_AXIMM_81_ARADDR),
        .AP_AXIMM_81_ARLEN(AP_AXIMM_81_ARLEN),
        .AP_AXIMM_81_ARSIZE(AP_AXIMM_81_ARSIZE),
        .AP_AXIMM_81_ARBURST(AP_AXIMM_81_ARBURST),
        .AP_AXIMM_81_ARLOCK(AP_AXIMM_81_ARLOCK),
        .AP_AXIMM_81_ARCACHE(AP_AXIMM_81_ARCACHE),
        .AP_AXIMM_81_ARPROT(AP_AXIMM_81_ARPROT),
        .AP_AXIMM_81_ARREGION(AP_AXIMM_81_ARREGION),
        .AP_AXIMM_81_ARQOS(AP_AXIMM_81_ARQOS),
        .AP_AXIMM_81_ARVALID(AP_AXIMM_81_ARVALID),
        .AP_AXIMM_81_ARREADY(AP_AXIMM_81_ARREADY),
        .AP_AXIMM_81_RDATA(AP_AXIMM_81_RDATA),
        .AP_AXIMM_81_RRESP(AP_AXIMM_81_RRESP),
        .AP_AXIMM_81_RLAST(AP_AXIMM_81_RLAST),
        .AP_AXIMM_81_RVALID(AP_AXIMM_81_RVALID),
        .AP_AXIMM_81_RREADY(AP_AXIMM_81_RREADY),
        .M_AXIMM_81_AWADDR(M_AXIMM_81_AWADDR),
        .M_AXIMM_81_AWLEN(M_AXIMM_81_AWLEN),
        .M_AXIMM_81_AWSIZE(M_AXIMM_81_AWSIZE),
        .M_AXIMM_81_AWBURST(M_AXIMM_81_AWBURST),
        .M_AXIMM_81_AWLOCK(M_AXIMM_81_AWLOCK),
        .M_AXIMM_81_AWCACHE(M_AXIMM_81_AWCACHE),
        .M_AXIMM_81_AWPROT(M_AXIMM_81_AWPROT),
        .M_AXIMM_81_AWREGION(M_AXIMM_81_AWREGION),
        .M_AXIMM_81_AWQOS(M_AXIMM_81_AWQOS),
        .M_AXIMM_81_AWVALID(M_AXIMM_81_AWVALID),
        .M_AXIMM_81_AWREADY(M_AXIMM_81_AWREADY),
        .M_AXIMM_81_WDATA(M_AXIMM_81_WDATA),
        .M_AXIMM_81_WSTRB(M_AXIMM_81_WSTRB),
        .M_AXIMM_81_WLAST(M_AXIMM_81_WLAST),
        .M_AXIMM_81_WVALID(M_AXIMM_81_WVALID),
        .M_AXIMM_81_WREADY(M_AXIMM_81_WREADY),
        .M_AXIMM_81_BRESP(M_AXIMM_81_BRESP),
        .M_AXIMM_81_BVALID(M_AXIMM_81_BVALID),
        .M_AXIMM_81_BREADY(M_AXIMM_81_BREADY),
        .M_AXIMM_81_ARADDR(M_AXIMM_81_ARADDR),
        .M_AXIMM_81_ARLEN(M_AXIMM_81_ARLEN),
        .M_AXIMM_81_ARSIZE(M_AXIMM_81_ARSIZE),
        .M_AXIMM_81_ARBURST(M_AXIMM_81_ARBURST),
        .M_AXIMM_81_ARLOCK(M_AXIMM_81_ARLOCK),
        .M_AXIMM_81_ARCACHE(M_AXIMM_81_ARCACHE),
        .M_AXIMM_81_ARPROT(M_AXIMM_81_ARPROT),
        .M_AXIMM_81_ARREGION(M_AXIMM_81_ARREGION),
        .M_AXIMM_81_ARQOS(M_AXIMM_81_ARQOS),
        .M_AXIMM_81_ARVALID(M_AXIMM_81_ARVALID),
        .M_AXIMM_81_ARREADY(M_AXIMM_81_ARREADY),
        .M_AXIMM_81_RDATA(M_AXIMM_81_RDATA),
        .M_AXIMM_81_RRESP(M_AXIMM_81_RRESP),
        .M_AXIMM_81_RLAST(M_AXIMM_81_RLAST),
        .M_AXIMM_81_RVALID(M_AXIMM_81_RVALID),
        .M_AXIMM_81_RREADY(M_AXIMM_81_RREADY),
        .AP_AXIMM_82_AWADDR(AP_AXIMM_82_AWADDR),
        .AP_AXIMM_82_AWLEN(AP_AXIMM_82_AWLEN),
        .AP_AXIMM_82_AWSIZE(AP_AXIMM_82_AWSIZE),
        .AP_AXIMM_82_AWBURST(AP_AXIMM_82_AWBURST),
        .AP_AXIMM_82_AWLOCK(AP_AXIMM_82_AWLOCK),
        .AP_AXIMM_82_AWCACHE(AP_AXIMM_82_AWCACHE),
        .AP_AXIMM_82_AWPROT(AP_AXIMM_82_AWPROT),
        .AP_AXIMM_82_AWREGION(AP_AXIMM_82_AWREGION),
        .AP_AXIMM_82_AWQOS(AP_AXIMM_82_AWQOS),
        .AP_AXIMM_82_AWVALID(AP_AXIMM_82_AWVALID),
        .AP_AXIMM_82_AWREADY(AP_AXIMM_82_AWREADY),
        .AP_AXIMM_82_WDATA(AP_AXIMM_82_WDATA),
        .AP_AXIMM_82_WSTRB(AP_AXIMM_82_WSTRB),
        .AP_AXIMM_82_WLAST(AP_AXIMM_82_WLAST),
        .AP_AXIMM_82_WVALID(AP_AXIMM_82_WVALID),
        .AP_AXIMM_82_WREADY(AP_AXIMM_82_WREADY),
        .AP_AXIMM_82_BRESP(AP_AXIMM_82_BRESP),
        .AP_AXIMM_82_BVALID(AP_AXIMM_82_BVALID),
        .AP_AXIMM_82_BREADY(AP_AXIMM_82_BREADY),
        .AP_AXIMM_82_ARADDR(AP_AXIMM_82_ARADDR),
        .AP_AXIMM_82_ARLEN(AP_AXIMM_82_ARLEN),
        .AP_AXIMM_82_ARSIZE(AP_AXIMM_82_ARSIZE),
        .AP_AXIMM_82_ARBURST(AP_AXIMM_82_ARBURST),
        .AP_AXIMM_82_ARLOCK(AP_AXIMM_82_ARLOCK),
        .AP_AXIMM_82_ARCACHE(AP_AXIMM_82_ARCACHE),
        .AP_AXIMM_82_ARPROT(AP_AXIMM_82_ARPROT),
        .AP_AXIMM_82_ARREGION(AP_AXIMM_82_ARREGION),
        .AP_AXIMM_82_ARQOS(AP_AXIMM_82_ARQOS),
        .AP_AXIMM_82_ARVALID(AP_AXIMM_82_ARVALID),
        .AP_AXIMM_82_ARREADY(AP_AXIMM_82_ARREADY),
        .AP_AXIMM_82_RDATA(AP_AXIMM_82_RDATA),
        .AP_AXIMM_82_RRESP(AP_AXIMM_82_RRESP),
        .AP_AXIMM_82_RLAST(AP_AXIMM_82_RLAST),
        .AP_AXIMM_82_RVALID(AP_AXIMM_82_RVALID),
        .AP_AXIMM_82_RREADY(AP_AXIMM_82_RREADY),
        .M_AXIMM_82_AWADDR(M_AXIMM_82_AWADDR),
        .M_AXIMM_82_AWLEN(M_AXIMM_82_AWLEN),
        .M_AXIMM_82_AWSIZE(M_AXIMM_82_AWSIZE),
        .M_AXIMM_82_AWBURST(M_AXIMM_82_AWBURST),
        .M_AXIMM_82_AWLOCK(M_AXIMM_82_AWLOCK),
        .M_AXIMM_82_AWCACHE(M_AXIMM_82_AWCACHE),
        .M_AXIMM_82_AWPROT(M_AXIMM_82_AWPROT),
        .M_AXIMM_82_AWREGION(M_AXIMM_82_AWREGION),
        .M_AXIMM_82_AWQOS(M_AXIMM_82_AWQOS),
        .M_AXIMM_82_AWVALID(M_AXIMM_82_AWVALID),
        .M_AXIMM_82_AWREADY(M_AXIMM_82_AWREADY),
        .M_AXIMM_82_WDATA(M_AXIMM_82_WDATA),
        .M_AXIMM_82_WSTRB(M_AXIMM_82_WSTRB),
        .M_AXIMM_82_WLAST(M_AXIMM_82_WLAST),
        .M_AXIMM_82_WVALID(M_AXIMM_82_WVALID),
        .M_AXIMM_82_WREADY(M_AXIMM_82_WREADY),
        .M_AXIMM_82_BRESP(M_AXIMM_82_BRESP),
        .M_AXIMM_82_BVALID(M_AXIMM_82_BVALID),
        .M_AXIMM_82_BREADY(M_AXIMM_82_BREADY),
        .M_AXIMM_82_ARADDR(M_AXIMM_82_ARADDR),
        .M_AXIMM_82_ARLEN(M_AXIMM_82_ARLEN),
        .M_AXIMM_82_ARSIZE(M_AXIMM_82_ARSIZE),
        .M_AXIMM_82_ARBURST(M_AXIMM_82_ARBURST),
        .M_AXIMM_82_ARLOCK(M_AXIMM_82_ARLOCK),
        .M_AXIMM_82_ARCACHE(M_AXIMM_82_ARCACHE),
        .M_AXIMM_82_ARPROT(M_AXIMM_82_ARPROT),
        .M_AXIMM_82_ARREGION(M_AXIMM_82_ARREGION),
        .M_AXIMM_82_ARQOS(M_AXIMM_82_ARQOS),
        .M_AXIMM_82_ARVALID(M_AXIMM_82_ARVALID),
        .M_AXIMM_82_ARREADY(M_AXIMM_82_ARREADY),
        .M_AXIMM_82_RDATA(M_AXIMM_82_RDATA),
        .M_AXIMM_82_RRESP(M_AXIMM_82_RRESP),
        .M_AXIMM_82_RLAST(M_AXIMM_82_RLAST),
        .M_AXIMM_82_RVALID(M_AXIMM_82_RVALID),
        .M_AXIMM_82_RREADY(M_AXIMM_82_RREADY),
        .AP_AXIMM_83_AWADDR(AP_AXIMM_83_AWADDR),
        .AP_AXIMM_83_AWLEN(AP_AXIMM_83_AWLEN),
        .AP_AXIMM_83_AWSIZE(AP_AXIMM_83_AWSIZE),
        .AP_AXIMM_83_AWBURST(AP_AXIMM_83_AWBURST),
        .AP_AXIMM_83_AWLOCK(AP_AXIMM_83_AWLOCK),
        .AP_AXIMM_83_AWCACHE(AP_AXIMM_83_AWCACHE),
        .AP_AXIMM_83_AWPROT(AP_AXIMM_83_AWPROT),
        .AP_AXIMM_83_AWREGION(AP_AXIMM_83_AWREGION),
        .AP_AXIMM_83_AWQOS(AP_AXIMM_83_AWQOS),
        .AP_AXIMM_83_AWVALID(AP_AXIMM_83_AWVALID),
        .AP_AXIMM_83_AWREADY(AP_AXIMM_83_AWREADY),
        .AP_AXIMM_83_WDATA(AP_AXIMM_83_WDATA),
        .AP_AXIMM_83_WSTRB(AP_AXIMM_83_WSTRB),
        .AP_AXIMM_83_WLAST(AP_AXIMM_83_WLAST),
        .AP_AXIMM_83_WVALID(AP_AXIMM_83_WVALID),
        .AP_AXIMM_83_WREADY(AP_AXIMM_83_WREADY),
        .AP_AXIMM_83_BRESP(AP_AXIMM_83_BRESP),
        .AP_AXIMM_83_BVALID(AP_AXIMM_83_BVALID),
        .AP_AXIMM_83_BREADY(AP_AXIMM_83_BREADY),
        .AP_AXIMM_83_ARADDR(AP_AXIMM_83_ARADDR),
        .AP_AXIMM_83_ARLEN(AP_AXIMM_83_ARLEN),
        .AP_AXIMM_83_ARSIZE(AP_AXIMM_83_ARSIZE),
        .AP_AXIMM_83_ARBURST(AP_AXIMM_83_ARBURST),
        .AP_AXIMM_83_ARLOCK(AP_AXIMM_83_ARLOCK),
        .AP_AXIMM_83_ARCACHE(AP_AXIMM_83_ARCACHE),
        .AP_AXIMM_83_ARPROT(AP_AXIMM_83_ARPROT),
        .AP_AXIMM_83_ARREGION(AP_AXIMM_83_ARREGION),
        .AP_AXIMM_83_ARQOS(AP_AXIMM_83_ARQOS),
        .AP_AXIMM_83_ARVALID(AP_AXIMM_83_ARVALID),
        .AP_AXIMM_83_ARREADY(AP_AXIMM_83_ARREADY),
        .AP_AXIMM_83_RDATA(AP_AXIMM_83_RDATA),
        .AP_AXIMM_83_RRESP(AP_AXIMM_83_RRESP),
        .AP_AXIMM_83_RLAST(AP_AXIMM_83_RLAST),
        .AP_AXIMM_83_RVALID(AP_AXIMM_83_RVALID),
        .AP_AXIMM_83_RREADY(AP_AXIMM_83_RREADY),
        .M_AXIMM_83_AWADDR(M_AXIMM_83_AWADDR),
        .M_AXIMM_83_AWLEN(M_AXIMM_83_AWLEN),
        .M_AXIMM_83_AWSIZE(M_AXIMM_83_AWSIZE),
        .M_AXIMM_83_AWBURST(M_AXIMM_83_AWBURST),
        .M_AXIMM_83_AWLOCK(M_AXIMM_83_AWLOCK),
        .M_AXIMM_83_AWCACHE(M_AXIMM_83_AWCACHE),
        .M_AXIMM_83_AWPROT(M_AXIMM_83_AWPROT),
        .M_AXIMM_83_AWREGION(M_AXIMM_83_AWREGION),
        .M_AXIMM_83_AWQOS(M_AXIMM_83_AWQOS),
        .M_AXIMM_83_AWVALID(M_AXIMM_83_AWVALID),
        .M_AXIMM_83_AWREADY(M_AXIMM_83_AWREADY),
        .M_AXIMM_83_WDATA(M_AXIMM_83_WDATA),
        .M_AXIMM_83_WSTRB(M_AXIMM_83_WSTRB),
        .M_AXIMM_83_WLAST(M_AXIMM_83_WLAST),
        .M_AXIMM_83_WVALID(M_AXIMM_83_WVALID),
        .M_AXIMM_83_WREADY(M_AXIMM_83_WREADY),
        .M_AXIMM_83_BRESP(M_AXIMM_83_BRESP),
        .M_AXIMM_83_BVALID(M_AXIMM_83_BVALID),
        .M_AXIMM_83_BREADY(M_AXIMM_83_BREADY),
        .M_AXIMM_83_ARADDR(M_AXIMM_83_ARADDR),
        .M_AXIMM_83_ARLEN(M_AXIMM_83_ARLEN),
        .M_AXIMM_83_ARSIZE(M_AXIMM_83_ARSIZE),
        .M_AXIMM_83_ARBURST(M_AXIMM_83_ARBURST),
        .M_AXIMM_83_ARLOCK(M_AXIMM_83_ARLOCK),
        .M_AXIMM_83_ARCACHE(M_AXIMM_83_ARCACHE),
        .M_AXIMM_83_ARPROT(M_AXIMM_83_ARPROT),
        .M_AXIMM_83_ARREGION(M_AXIMM_83_ARREGION),
        .M_AXIMM_83_ARQOS(M_AXIMM_83_ARQOS),
        .M_AXIMM_83_ARVALID(M_AXIMM_83_ARVALID),
        .M_AXIMM_83_ARREADY(M_AXIMM_83_ARREADY),
        .M_AXIMM_83_RDATA(M_AXIMM_83_RDATA),
        .M_AXIMM_83_RRESP(M_AXIMM_83_RRESP),
        .M_AXIMM_83_RLAST(M_AXIMM_83_RLAST),
        .M_AXIMM_83_RVALID(M_AXIMM_83_RVALID),
        .M_AXIMM_83_RREADY(M_AXIMM_83_RREADY),
        .AP_AXIMM_84_AWADDR(AP_AXIMM_84_AWADDR),
        .AP_AXIMM_84_AWLEN(AP_AXIMM_84_AWLEN),
        .AP_AXIMM_84_AWSIZE(AP_AXIMM_84_AWSIZE),
        .AP_AXIMM_84_AWBURST(AP_AXIMM_84_AWBURST),
        .AP_AXIMM_84_AWLOCK(AP_AXIMM_84_AWLOCK),
        .AP_AXIMM_84_AWCACHE(AP_AXIMM_84_AWCACHE),
        .AP_AXIMM_84_AWPROT(AP_AXIMM_84_AWPROT),
        .AP_AXIMM_84_AWREGION(AP_AXIMM_84_AWREGION),
        .AP_AXIMM_84_AWQOS(AP_AXIMM_84_AWQOS),
        .AP_AXIMM_84_AWVALID(AP_AXIMM_84_AWVALID),
        .AP_AXIMM_84_AWREADY(AP_AXIMM_84_AWREADY),
        .AP_AXIMM_84_WDATA(AP_AXIMM_84_WDATA),
        .AP_AXIMM_84_WSTRB(AP_AXIMM_84_WSTRB),
        .AP_AXIMM_84_WLAST(AP_AXIMM_84_WLAST),
        .AP_AXIMM_84_WVALID(AP_AXIMM_84_WVALID),
        .AP_AXIMM_84_WREADY(AP_AXIMM_84_WREADY),
        .AP_AXIMM_84_BRESP(AP_AXIMM_84_BRESP),
        .AP_AXIMM_84_BVALID(AP_AXIMM_84_BVALID),
        .AP_AXIMM_84_BREADY(AP_AXIMM_84_BREADY),
        .AP_AXIMM_84_ARADDR(AP_AXIMM_84_ARADDR),
        .AP_AXIMM_84_ARLEN(AP_AXIMM_84_ARLEN),
        .AP_AXIMM_84_ARSIZE(AP_AXIMM_84_ARSIZE),
        .AP_AXIMM_84_ARBURST(AP_AXIMM_84_ARBURST),
        .AP_AXIMM_84_ARLOCK(AP_AXIMM_84_ARLOCK),
        .AP_AXIMM_84_ARCACHE(AP_AXIMM_84_ARCACHE),
        .AP_AXIMM_84_ARPROT(AP_AXIMM_84_ARPROT),
        .AP_AXIMM_84_ARREGION(AP_AXIMM_84_ARREGION),
        .AP_AXIMM_84_ARQOS(AP_AXIMM_84_ARQOS),
        .AP_AXIMM_84_ARVALID(AP_AXIMM_84_ARVALID),
        .AP_AXIMM_84_ARREADY(AP_AXIMM_84_ARREADY),
        .AP_AXIMM_84_RDATA(AP_AXIMM_84_RDATA),
        .AP_AXIMM_84_RRESP(AP_AXIMM_84_RRESP),
        .AP_AXIMM_84_RLAST(AP_AXIMM_84_RLAST),
        .AP_AXIMM_84_RVALID(AP_AXIMM_84_RVALID),
        .AP_AXIMM_84_RREADY(AP_AXIMM_84_RREADY),
        .M_AXIMM_84_AWADDR(M_AXIMM_84_AWADDR),
        .M_AXIMM_84_AWLEN(M_AXIMM_84_AWLEN),
        .M_AXIMM_84_AWSIZE(M_AXIMM_84_AWSIZE),
        .M_AXIMM_84_AWBURST(M_AXIMM_84_AWBURST),
        .M_AXIMM_84_AWLOCK(M_AXIMM_84_AWLOCK),
        .M_AXIMM_84_AWCACHE(M_AXIMM_84_AWCACHE),
        .M_AXIMM_84_AWPROT(M_AXIMM_84_AWPROT),
        .M_AXIMM_84_AWREGION(M_AXIMM_84_AWREGION),
        .M_AXIMM_84_AWQOS(M_AXIMM_84_AWQOS),
        .M_AXIMM_84_AWVALID(M_AXIMM_84_AWVALID),
        .M_AXIMM_84_AWREADY(M_AXIMM_84_AWREADY),
        .M_AXIMM_84_WDATA(M_AXIMM_84_WDATA),
        .M_AXIMM_84_WSTRB(M_AXIMM_84_WSTRB),
        .M_AXIMM_84_WLAST(M_AXIMM_84_WLAST),
        .M_AXIMM_84_WVALID(M_AXIMM_84_WVALID),
        .M_AXIMM_84_WREADY(M_AXIMM_84_WREADY),
        .M_AXIMM_84_BRESP(M_AXIMM_84_BRESP),
        .M_AXIMM_84_BVALID(M_AXIMM_84_BVALID),
        .M_AXIMM_84_BREADY(M_AXIMM_84_BREADY),
        .M_AXIMM_84_ARADDR(M_AXIMM_84_ARADDR),
        .M_AXIMM_84_ARLEN(M_AXIMM_84_ARLEN),
        .M_AXIMM_84_ARSIZE(M_AXIMM_84_ARSIZE),
        .M_AXIMM_84_ARBURST(M_AXIMM_84_ARBURST),
        .M_AXIMM_84_ARLOCK(M_AXIMM_84_ARLOCK),
        .M_AXIMM_84_ARCACHE(M_AXIMM_84_ARCACHE),
        .M_AXIMM_84_ARPROT(M_AXIMM_84_ARPROT),
        .M_AXIMM_84_ARREGION(M_AXIMM_84_ARREGION),
        .M_AXIMM_84_ARQOS(M_AXIMM_84_ARQOS),
        .M_AXIMM_84_ARVALID(M_AXIMM_84_ARVALID),
        .M_AXIMM_84_ARREADY(M_AXIMM_84_ARREADY),
        .M_AXIMM_84_RDATA(M_AXIMM_84_RDATA),
        .M_AXIMM_84_RRESP(M_AXIMM_84_RRESP),
        .M_AXIMM_84_RLAST(M_AXIMM_84_RLAST),
        .M_AXIMM_84_RVALID(M_AXIMM_84_RVALID),
        .M_AXIMM_84_RREADY(M_AXIMM_84_RREADY),
        .AP_AXIMM_85_AWADDR(AP_AXIMM_85_AWADDR),
        .AP_AXIMM_85_AWLEN(AP_AXIMM_85_AWLEN),
        .AP_AXIMM_85_AWSIZE(AP_AXIMM_85_AWSIZE),
        .AP_AXIMM_85_AWBURST(AP_AXIMM_85_AWBURST),
        .AP_AXIMM_85_AWLOCK(AP_AXIMM_85_AWLOCK),
        .AP_AXIMM_85_AWCACHE(AP_AXIMM_85_AWCACHE),
        .AP_AXIMM_85_AWPROT(AP_AXIMM_85_AWPROT),
        .AP_AXIMM_85_AWREGION(AP_AXIMM_85_AWREGION),
        .AP_AXIMM_85_AWQOS(AP_AXIMM_85_AWQOS),
        .AP_AXIMM_85_AWVALID(AP_AXIMM_85_AWVALID),
        .AP_AXIMM_85_AWREADY(AP_AXIMM_85_AWREADY),
        .AP_AXIMM_85_WDATA(AP_AXIMM_85_WDATA),
        .AP_AXIMM_85_WSTRB(AP_AXIMM_85_WSTRB),
        .AP_AXIMM_85_WLAST(AP_AXIMM_85_WLAST),
        .AP_AXIMM_85_WVALID(AP_AXIMM_85_WVALID),
        .AP_AXIMM_85_WREADY(AP_AXIMM_85_WREADY),
        .AP_AXIMM_85_BRESP(AP_AXIMM_85_BRESP),
        .AP_AXIMM_85_BVALID(AP_AXIMM_85_BVALID),
        .AP_AXIMM_85_BREADY(AP_AXIMM_85_BREADY),
        .AP_AXIMM_85_ARADDR(AP_AXIMM_85_ARADDR),
        .AP_AXIMM_85_ARLEN(AP_AXIMM_85_ARLEN),
        .AP_AXIMM_85_ARSIZE(AP_AXIMM_85_ARSIZE),
        .AP_AXIMM_85_ARBURST(AP_AXIMM_85_ARBURST),
        .AP_AXIMM_85_ARLOCK(AP_AXIMM_85_ARLOCK),
        .AP_AXIMM_85_ARCACHE(AP_AXIMM_85_ARCACHE),
        .AP_AXIMM_85_ARPROT(AP_AXIMM_85_ARPROT),
        .AP_AXIMM_85_ARREGION(AP_AXIMM_85_ARREGION),
        .AP_AXIMM_85_ARQOS(AP_AXIMM_85_ARQOS),
        .AP_AXIMM_85_ARVALID(AP_AXIMM_85_ARVALID),
        .AP_AXIMM_85_ARREADY(AP_AXIMM_85_ARREADY),
        .AP_AXIMM_85_RDATA(AP_AXIMM_85_RDATA),
        .AP_AXIMM_85_RRESP(AP_AXIMM_85_RRESP),
        .AP_AXIMM_85_RLAST(AP_AXIMM_85_RLAST),
        .AP_AXIMM_85_RVALID(AP_AXIMM_85_RVALID),
        .AP_AXIMM_85_RREADY(AP_AXIMM_85_RREADY),
        .M_AXIMM_85_AWADDR(M_AXIMM_85_AWADDR),
        .M_AXIMM_85_AWLEN(M_AXIMM_85_AWLEN),
        .M_AXIMM_85_AWSIZE(M_AXIMM_85_AWSIZE),
        .M_AXIMM_85_AWBURST(M_AXIMM_85_AWBURST),
        .M_AXIMM_85_AWLOCK(M_AXIMM_85_AWLOCK),
        .M_AXIMM_85_AWCACHE(M_AXIMM_85_AWCACHE),
        .M_AXIMM_85_AWPROT(M_AXIMM_85_AWPROT),
        .M_AXIMM_85_AWREGION(M_AXIMM_85_AWREGION),
        .M_AXIMM_85_AWQOS(M_AXIMM_85_AWQOS),
        .M_AXIMM_85_AWVALID(M_AXIMM_85_AWVALID),
        .M_AXIMM_85_AWREADY(M_AXIMM_85_AWREADY),
        .M_AXIMM_85_WDATA(M_AXIMM_85_WDATA),
        .M_AXIMM_85_WSTRB(M_AXIMM_85_WSTRB),
        .M_AXIMM_85_WLAST(M_AXIMM_85_WLAST),
        .M_AXIMM_85_WVALID(M_AXIMM_85_WVALID),
        .M_AXIMM_85_WREADY(M_AXIMM_85_WREADY),
        .M_AXIMM_85_BRESP(M_AXIMM_85_BRESP),
        .M_AXIMM_85_BVALID(M_AXIMM_85_BVALID),
        .M_AXIMM_85_BREADY(M_AXIMM_85_BREADY),
        .M_AXIMM_85_ARADDR(M_AXIMM_85_ARADDR),
        .M_AXIMM_85_ARLEN(M_AXIMM_85_ARLEN),
        .M_AXIMM_85_ARSIZE(M_AXIMM_85_ARSIZE),
        .M_AXIMM_85_ARBURST(M_AXIMM_85_ARBURST),
        .M_AXIMM_85_ARLOCK(M_AXIMM_85_ARLOCK),
        .M_AXIMM_85_ARCACHE(M_AXIMM_85_ARCACHE),
        .M_AXIMM_85_ARPROT(M_AXIMM_85_ARPROT),
        .M_AXIMM_85_ARREGION(M_AXIMM_85_ARREGION),
        .M_AXIMM_85_ARQOS(M_AXIMM_85_ARQOS),
        .M_AXIMM_85_ARVALID(M_AXIMM_85_ARVALID),
        .M_AXIMM_85_ARREADY(M_AXIMM_85_ARREADY),
        .M_AXIMM_85_RDATA(M_AXIMM_85_RDATA),
        .M_AXIMM_85_RRESP(M_AXIMM_85_RRESP),
        .M_AXIMM_85_RLAST(M_AXIMM_85_RLAST),
        .M_AXIMM_85_RVALID(M_AXIMM_85_RVALID),
        .M_AXIMM_85_RREADY(M_AXIMM_85_RREADY),
        .AP_AXIMM_86_AWADDR(AP_AXIMM_86_AWADDR),
        .AP_AXIMM_86_AWLEN(AP_AXIMM_86_AWLEN),
        .AP_AXIMM_86_AWSIZE(AP_AXIMM_86_AWSIZE),
        .AP_AXIMM_86_AWBURST(AP_AXIMM_86_AWBURST),
        .AP_AXIMM_86_AWLOCK(AP_AXIMM_86_AWLOCK),
        .AP_AXIMM_86_AWCACHE(AP_AXIMM_86_AWCACHE),
        .AP_AXIMM_86_AWPROT(AP_AXIMM_86_AWPROT),
        .AP_AXIMM_86_AWREGION(AP_AXIMM_86_AWREGION),
        .AP_AXIMM_86_AWQOS(AP_AXIMM_86_AWQOS),
        .AP_AXIMM_86_AWVALID(AP_AXIMM_86_AWVALID),
        .AP_AXIMM_86_AWREADY(AP_AXIMM_86_AWREADY),
        .AP_AXIMM_86_WDATA(AP_AXIMM_86_WDATA),
        .AP_AXIMM_86_WSTRB(AP_AXIMM_86_WSTRB),
        .AP_AXIMM_86_WLAST(AP_AXIMM_86_WLAST),
        .AP_AXIMM_86_WVALID(AP_AXIMM_86_WVALID),
        .AP_AXIMM_86_WREADY(AP_AXIMM_86_WREADY),
        .AP_AXIMM_86_BRESP(AP_AXIMM_86_BRESP),
        .AP_AXIMM_86_BVALID(AP_AXIMM_86_BVALID),
        .AP_AXIMM_86_BREADY(AP_AXIMM_86_BREADY),
        .AP_AXIMM_86_ARADDR(AP_AXIMM_86_ARADDR),
        .AP_AXIMM_86_ARLEN(AP_AXIMM_86_ARLEN),
        .AP_AXIMM_86_ARSIZE(AP_AXIMM_86_ARSIZE),
        .AP_AXIMM_86_ARBURST(AP_AXIMM_86_ARBURST),
        .AP_AXIMM_86_ARLOCK(AP_AXIMM_86_ARLOCK),
        .AP_AXIMM_86_ARCACHE(AP_AXIMM_86_ARCACHE),
        .AP_AXIMM_86_ARPROT(AP_AXIMM_86_ARPROT),
        .AP_AXIMM_86_ARREGION(AP_AXIMM_86_ARREGION),
        .AP_AXIMM_86_ARQOS(AP_AXIMM_86_ARQOS),
        .AP_AXIMM_86_ARVALID(AP_AXIMM_86_ARVALID),
        .AP_AXIMM_86_ARREADY(AP_AXIMM_86_ARREADY),
        .AP_AXIMM_86_RDATA(AP_AXIMM_86_RDATA),
        .AP_AXIMM_86_RRESP(AP_AXIMM_86_RRESP),
        .AP_AXIMM_86_RLAST(AP_AXIMM_86_RLAST),
        .AP_AXIMM_86_RVALID(AP_AXIMM_86_RVALID),
        .AP_AXIMM_86_RREADY(AP_AXIMM_86_RREADY),
        .M_AXIMM_86_AWADDR(M_AXIMM_86_AWADDR),
        .M_AXIMM_86_AWLEN(M_AXIMM_86_AWLEN),
        .M_AXIMM_86_AWSIZE(M_AXIMM_86_AWSIZE),
        .M_AXIMM_86_AWBURST(M_AXIMM_86_AWBURST),
        .M_AXIMM_86_AWLOCK(M_AXIMM_86_AWLOCK),
        .M_AXIMM_86_AWCACHE(M_AXIMM_86_AWCACHE),
        .M_AXIMM_86_AWPROT(M_AXIMM_86_AWPROT),
        .M_AXIMM_86_AWREGION(M_AXIMM_86_AWREGION),
        .M_AXIMM_86_AWQOS(M_AXIMM_86_AWQOS),
        .M_AXIMM_86_AWVALID(M_AXIMM_86_AWVALID),
        .M_AXIMM_86_AWREADY(M_AXIMM_86_AWREADY),
        .M_AXIMM_86_WDATA(M_AXIMM_86_WDATA),
        .M_AXIMM_86_WSTRB(M_AXIMM_86_WSTRB),
        .M_AXIMM_86_WLAST(M_AXIMM_86_WLAST),
        .M_AXIMM_86_WVALID(M_AXIMM_86_WVALID),
        .M_AXIMM_86_WREADY(M_AXIMM_86_WREADY),
        .M_AXIMM_86_BRESP(M_AXIMM_86_BRESP),
        .M_AXIMM_86_BVALID(M_AXIMM_86_BVALID),
        .M_AXIMM_86_BREADY(M_AXIMM_86_BREADY),
        .M_AXIMM_86_ARADDR(M_AXIMM_86_ARADDR),
        .M_AXIMM_86_ARLEN(M_AXIMM_86_ARLEN),
        .M_AXIMM_86_ARSIZE(M_AXIMM_86_ARSIZE),
        .M_AXIMM_86_ARBURST(M_AXIMM_86_ARBURST),
        .M_AXIMM_86_ARLOCK(M_AXIMM_86_ARLOCK),
        .M_AXIMM_86_ARCACHE(M_AXIMM_86_ARCACHE),
        .M_AXIMM_86_ARPROT(M_AXIMM_86_ARPROT),
        .M_AXIMM_86_ARREGION(M_AXIMM_86_ARREGION),
        .M_AXIMM_86_ARQOS(M_AXIMM_86_ARQOS),
        .M_AXIMM_86_ARVALID(M_AXIMM_86_ARVALID),
        .M_AXIMM_86_ARREADY(M_AXIMM_86_ARREADY),
        .M_AXIMM_86_RDATA(M_AXIMM_86_RDATA),
        .M_AXIMM_86_RRESP(M_AXIMM_86_RRESP),
        .M_AXIMM_86_RLAST(M_AXIMM_86_RLAST),
        .M_AXIMM_86_RVALID(M_AXIMM_86_RVALID),
        .M_AXIMM_86_RREADY(M_AXIMM_86_RREADY),
        .AP_AXIMM_87_AWADDR(AP_AXIMM_87_AWADDR),
        .AP_AXIMM_87_AWLEN(AP_AXIMM_87_AWLEN),
        .AP_AXIMM_87_AWSIZE(AP_AXIMM_87_AWSIZE),
        .AP_AXIMM_87_AWBURST(AP_AXIMM_87_AWBURST),
        .AP_AXIMM_87_AWLOCK(AP_AXIMM_87_AWLOCK),
        .AP_AXIMM_87_AWCACHE(AP_AXIMM_87_AWCACHE),
        .AP_AXIMM_87_AWPROT(AP_AXIMM_87_AWPROT),
        .AP_AXIMM_87_AWREGION(AP_AXIMM_87_AWREGION),
        .AP_AXIMM_87_AWQOS(AP_AXIMM_87_AWQOS),
        .AP_AXIMM_87_AWVALID(AP_AXIMM_87_AWVALID),
        .AP_AXIMM_87_AWREADY(AP_AXIMM_87_AWREADY),
        .AP_AXIMM_87_WDATA(AP_AXIMM_87_WDATA),
        .AP_AXIMM_87_WSTRB(AP_AXIMM_87_WSTRB),
        .AP_AXIMM_87_WLAST(AP_AXIMM_87_WLAST),
        .AP_AXIMM_87_WVALID(AP_AXIMM_87_WVALID),
        .AP_AXIMM_87_WREADY(AP_AXIMM_87_WREADY),
        .AP_AXIMM_87_BRESP(AP_AXIMM_87_BRESP),
        .AP_AXIMM_87_BVALID(AP_AXIMM_87_BVALID),
        .AP_AXIMM_87_BREADY(AP_AXIMM_87_BREADY),
        .AP_AXIMM_87_ARADDR(AP_AXIMM_87_ARADDR),
        .AP_AXIMM_87_ARLEN(AP_AXIMM_87_ARLEN),
        .AP_AXIMM_87_ARSIZE(AP_AXIMM_87_ARSIZE),
        .AP_AXIMM_87_ARBURST(AP_AXIMM_87_ARBURST),
        .AP_AXIMM_87_ARLOCK(AP_AXIMM_87_ARLOCK),
        .AP_AXIMM_87_ARCACHE(AP_AXIMM_87_ARCACHE),
        .AP_AXIMM_87_ARPROT(AP_AXIMM_87_ARPROT),
        .AP_AXIMM_87_ARREGION(AP_AXIMM_87_ARREGION),
        .AP_AXIMM_87_ARQOS(AP_AXIMM_87_ARQOS),
        .AP_AXIMM_87_ARVALID(AP_AXIMM_87_ARVALID),
        .AP_AXIMM_87_ARREADY(AP_AXIMM_87_ARREADY),
        .AP_AXIMM_87_RDATA(AP_AXIMM_87_RDATA),
        .AP_AXIMM_87_RRESP(AP_AXIMM_87_RRESP),
        .AP_AXIMM_87_RLAST(AP_AXIMM_87_RLAST),
        .AP_AXIMM_87_RVALID(AP_AXIMM_87_RVALID),
        .AP_AXIMM_87_RREADY(AP_AXIMM_87_RREADY),
        .M_AXIMM_87_AWADDR(M_AXIMM_87_AWADDR),
        .M_AXIMM_87_AWLEN(M_AXIMM_87_AWLEN),
        .M_AXIMM_87_AWSIZE(M_AXIMM_87_AWSIZE),
        .M_AXIMM_87_AWBURST(M_AXIMM_87_AWBURST),
        .M_AXIMM_87_AWLOCK(M_AXIMM_87_AWLOCK),
        .M_AXIMM_87_AWCACHE(M_AXIMM_87_AWCACHE),
        .M_AXIMM_87_AWPROT(M_AXIMM_87_AWPROT),
        .M_AXIMM_87_AWREGION(M_AXIMM_87_AWREGION),
        .M_AXIMM_87_AWQOS(M_AXIMM_87_AWQOS),
        .M_AXIMM_87_AWVALID(M_AXIMM_87_AWVALID),
        .M_AXIMM_87_AWREADY(M_AXIMM_87_AWREADY),
        .M_AXIMM_87_WDATA(M_AXIMM_87_WDATA),
        .M_AXIMM_87_WSTRB(M_AXIMM_87_WSTRB),
        .M_AXIMM_87_WLAST(M_AXIMM_87_WLAST),
        .M_AXIMM_87_WVALID(M_AXIMM_87_WVALID),
        .M_AXIMM_87_WREADY(M_AXIMM_87_WREADY),
        .M_AXIMM_87_BRESP(M_AXIMM_87_BRESP),
        .M_AXIMM_87_BVALID(M_AXIMM_87_BVALID),
        .M_AXIMM_87_BREADY(M_AXIMM_87_BREADY),
        .M_AXIMM_87_ARADDR(M_AXIMM_87_ARADDR),
        .M_AXIMM_87_ARLEN(M_AXIMM_87_ARLEN),
        .M_AXIMM_87_ARSIZE(M_AXIMM_87_ARSIZE),
        .M_AXIMM_87_ARBURST(M_AXIMM_87_ARBURST),
        .M_AXIMM_87_ARLOCK(M_AXIMM_87_ARLOCK),
        .M_AXIMM_87_ARCACHE(M_AXIMM_87_ARCACHE),
        .M_AXIMM_87_ARPROT(M_AXIMM_87_ARPROT),
        .M_AXIMM_87_ARREGION(M_AXIMM_87_ARREGION),
        .M_AXIMM_87_ARQOS(M_AXIMM_87_ARQOS),
        .M_AXIMM_87_ARVALID(M_AXIMM_87_ARVALID),
        .M_AXIMM_87_ARREADY(M_AXIMM_87_ARREADY),
        .M_AXIMM_87_RDATA(M_AXIMM_87_RDATA),
        .M_AXIMM_87_RRESP(M_AXIMM_87_RRESP),
        .M_AXIMM_87_RLAST(M_AXIMM_87_RLAST),
        .M_AXIMM_87_RVALID(M_AXIMM_87_RVALID),
        .M_AXIMM_87_RREADY(M_AXIMM_87_RREADY),
        .AP_AXIMM_88_AWADDR(AP_AXIMM_88_AWADDR),
        .AP_AXIMM_88_AWLEN(AP_AXIMM_88_AWLEN),
        .AP_AXIMM_88_AWSIZE(AP_AXIMM_88_AWSIZE),
        .AP_AXIMM_88_AWBURST(AP_AXIMM_88_AWBURST),
        .AP_AXIMM_88_AWLOCK(AP_AXIMM_88_AWLOCK),
        .AP_AXIMM_88_AWCACHE(AP_AXIMM_88_AWCACHE),
        .AP_AXIMM_88_AWPROT(AP_AXIMM_88_AWPROT),
        .AP_AXIMM_88_AWREGION(AP_AXIMM_88_AWREGION),
        .AP_AXIMM_88_AWQOS(AP_AXIMM_88_AWQOS),
        .AP_AXIMM_88_AWVALID(AP_AXIMM_88_AWVALID),
        .AP_AXIMM_88_AWREADY(AP_AXIMM_88_AWREADY),
        .AP_AXIMM_88_WDATA(AP_AXIMM_88_WDATA),
        .AP_AXIMM_88_WSTRB(AP_AXIMM_88_WSTRB),
        .AP_AXIMM_88_WLAST(AP_AXIMM_88_WLAST),
        .AP_AXIMM_88_WVALID(AP_AXIMM_88_WVALID),
        .AP_AXIMM_88_WREADY(AP_AXIMM_88_WREADY),
        .AP_AXIMM_88_BRESP(AP_AXIMM_88_BRESP),
        .AP_AXIMM_88_BVALID(AP_AXIMM_88_BVALID),
        .AP_AXIMM_88_BREADY(AP_AXIMM_88_BREADY),
        .AP_AXIMM_88_ARADDR(AP_AXIMM_88_ARADDR),
        .AP_AXIMM_88_ARLEN(AP_AXIMM_88_ARLEN),
        .AP_AXIMM_88_ARSIZE(AP_AXIMM_88_ARSIZE),
        .AP_AXIMM_88_ARBURST(AP_AXIMM_88_ARBURST),
        .AP_AXIMM_88_ARLOCK(AP_AXIMM_88_ARLOCK),
        .AP_AXIMM_88_ARCACHE(AP_AXIMM_88_ARCACHE),
        .AP_AXIMM_88_ARPROT(AP_AXIMM_88_ARPROT),
        .AP_AXIMM_88_ARREGION(AP_AXIMM_88_ARREGION),
        .AP_AXIMM_88_ARQOS(AP_AXIMM_88_ARQOS),
        .AP_AXIMM_88_ARVALID(AP_AXIMM_88_ARVALID),
        .AP_AXIMM_88_ARREADY(AP_AXIMM_88_ARREADY),
        .AP_AXIMM_88_RDATA(AP_AXIMM_88_RDATA),
        .AP_AXIMM_88_RRESP(AP_AXIMM_88_RRESP),
        .AP_AXIMM_88_RLAST(AP_AXIMM_88_RLAST),
        .AP_AXIMM_88_RVALID(AP_AXIMM_88_RVALID),
        .AP_AXIMM_88_RREADY(AP_AXIMM_88_RREADY),
        .M_AXIMM_88_AWADDR(M_AXIMM_88_AWADDR),
        .M_AXIMM_88_AWLEN(M_AXIMM_88_AWLEN),
        .M_AXIMM_88_AWSIZE(M_AXIMM_88_AWSIZE),
        .M_AXIMM_88_AWBURST(M_AXIMM_88_AWBURST),
        .M_AXIMM_88_AWLOCK(M_AXIMM_88_AWLOCK),
        .M_AXIMM_88_AWCACHE(M_AXIMM_88_AWCACHE),
        .M_AXIMM_88_AWPROT(M_AXIMM_88_AWPROT),
        .M_AXIMM_88_AWREGION(M_AXIMM_88_AWREGION),
        .M_AXIMM_88_AWQOS(M_AXIMM_88_AWQOS),
        .M_AXIMM_88_AWVALID(M_AXIMM_88_AWVALID),
        .M_AXIMM_88_AWREADY(M_AXIMM_88_AWREADY),
        .M_AXIMM_88_WDATA(M_AXIMM_88_WDATA),
        .M_AXIMM_88_WSTRB(M_AXIMM_88_WSTRB),
        .M_AXIMM_88_WLAST(M_AXIMM_88_WLAST),
        .M_AXIMM_88_WVALID(M_AXIMM_88_WVALID),
        .M_AXIMM_88_WREADY(M_AXIMM_88_WREADY),
        .M_AXIMM_88_BRESP(M_AXIMM_88_BRESP),
        .M_AXIMM_88_BVALID(M_AXIMM_88_BVALID),
        .M_AXIMM_88_BREADY(M_AXIMM_88_BREADY),
        .M_AXIMM_88_ARADDR(M_AXIMM_88_ARADDR),
        .M_AXIMM_88_ARLEN(M_AXIMM_88_ARLEN),
        .M_AXIMM_88_ARSIZE(M_AXIMM_88_ARSIZE),
        .M_AXIMM_88_ARBURST(M_AXIMM_88_ARBURST),
        .M_AXIMM_88_ARLOCK(M_AXIMM_88_ARLOCK),
        .M_AXIMM_88_ARCACHE(M_AXIMM_88_ARCACHE),
        .M_AXIMM_88_ARPROT(M_AXIMM_88_ARPROT),
        .M_AXIMM_88_ARREGION(M_AXIMM_88_ARREGION),
        .M_AXIMM_88_ARQOS(M_AXIMM_88_ARQOS),
        .M_AXIMM_88_ARVALID(M_AXIMM_88_ARVALID),
        .M_AXIMM_88_ARREADY(M_AXIMM_88_ARREADY),
        .M_AXIMM_88_RDATA(M_AXIMM_88_RDATA),
        .M_AXIMM_88_RRESP(M_AXIMM_88_RRESP),
        .M_AXIMM_88_RLAST(M_AXIMM_88_RLAST),
        .M_AXIMM_88_RVALID(M_AXIMM_88_RVALID),
        .M_AXIMM_88_RREADY(M_AXIMM_88_RREADY),
        .AP_AXIMM_89_AWADDR(AP_AXIMM_89_AWADDR),
        .AP_AXIMM_89_AWLEN(AP_AXIMM_89_AWLEN),
        .AP_AXIMM_89_AWSIZE(AP_AXIMM_89_AWSIZE),
        .AP_AXIMM_89_AWBURST(AP_AXIMM_89_AWBURST),
        .AP_AXIMM_89_AWLOCK(AP_AXIMM_89_AWLOCK),
        .AP_AXIMM_89_AWCACHE(AP_AXIMM_89_AWCACHE),
        .AP_AXIMM_89_AWPROT(AP_AXIMM_89_AWPROT),
        .AP_AXIMM_89_AWREGION(AP_AXIMM_89_AWREGION),
        .AP_AXIMM_89_AWQOS(AP_AXIMM_89_AWQOS),
        .AP_AXIMM_89_AWVALID(AP_AXIMM_89_AWVALID),
        .AP_AXIMM_89_AWREADY(AP_AXIMM_89_AWREADY),
        .AP_AXIMM_89_WDATA(AP_AXIMM_89_WDATA),
        .AP_AXIMM_89_WSTRB(AP_AXIMM_89_WSTRB),
        .AP_AXIMM_89_WLAST(AP_AXIMM_89_WLAST),
        .AP_AXIMM_89_WVALID(AP_AXIMM_89_WVALID),
        .AP_AXIMM_89_WREADY(AP_AXIMM_89_WREADY),
        .AP_AXIMM_89_BRESP(AP_AXIMM_89_BRESP),
        .AP_AXIMM_89_BVALID(AP_AXIMM_89_BVALID),
        .AP_AXIMM_89_BREADY(AP_AXIMM_89_BREADY),
        .AP_AXIMM_89_ARADDR(AP_AXIMM_89_ARADDR),
        .AP_AXIMM_89_ARLEN(AP_AXIMM_89_ARLEN),
        .AP_AXIMM_89_ARSIZE(AP_AXIMM_89_ARSIZE),
        .AP_AXIMM_89_ARBURST(AP_AXIMM_89_ARBURST),
        .AP_AXIMM_89_ARLOCK(AP_AXIMM_89_ARLOCK),
        .AP_AXIMM_89_ARCACHE(AP_AXIMM_89_ARCACHE),
        .AP_AXIMM_89_ARPROT(AP_AXIMM_89_ARPROT),
        .AP_AXIMM_89_ARREGION(AP_AXIMM_89_ARREGION),
        .AP_AXIMM_89_ARQOS(AP_AXIMM_89_ARQOS),
        .AP_AXIMM_89_ARVALID(AP_AXIMM_89_ARVALID),
        .AP_AXIMM_89_ARREADY(AP_AXIMM_89_ARREADY),
        .AP_AXIMM_89_RDATA(AP_AXIMM_89_RDATA),
        .AP_AXIMM_89_RRESP(AP_AXIMM_89_RRESP),
        .AP_AXIMM_89_RLAST(AP_AXIMM_89_RLAST),
        .AP_AXIMM_89_RVALID(AP_AXIMM_89_RVALID),
        .AP_AXIMM_89_RREADY(AP_AXIMM_89_RREADY),
        .M_AXIMM_89_AWADDR(M_AXIMM_89_AWADDR),
        .M_AXIMM_89_AWLEN(M_AXIMM_89_AWLEN),
        .M_AXIMM_89_AWSIZE(M_AXIMM_89_AWSIZE),
        .M_AXIMM_89_AWBURST(M_AXIMM_89_AWBURST),
        .M_AXIMM_89_AWLOCK(M_AXIMM_89_AWLOCK),
        .M_AXIMM_89_AWCACHE(M_AXIMM_89_AWCACHE),
        .M_AXIMM_89_AWPROT(M_AXIMM_89_AWPROT),
        .M_AXIMM_89_AWREGION(M_AXIMM_89_AWREGION),
        .M_AXIMM_89_AWQOS(M_AXIMM_89_AWQOS),
        .M_AXIMM_89_AWVALID(M_AXIMM_89_AWVALID),
        .M_AXIMM_89_AWREADY(M_AXIMM_89_AWREADY),
        .M_AXIMM_89_WDATA(M_AXIMM_89_WDATA),
        .M_AXIMM_89_WSTRB(M_AXIMM_89_WSTRB),
        .M_AXIMM_89_WLAST(M_AXIMM_89_WLAST),
        .M_AXIMM_89_WVALID(M_AXIMM_89_WVALID),
        .M_AXIMM_89_WREADY(M_AXIMM_89_WREADY),
        .M_AXIMM_89_BRESP(M_AXIMM_89_BRESP),
        .M_AXIMM_89_BVALID(M_AXIMM_89_BVALID),
        .M_AXIMM_89_BREADY(M_AXIMM_89_BREADY),
        .M_AXIMM_89_ARADDR(M_AXIMM_89_ARADDR),
        .M_AXIMM_89_ARLEN(M_AXIMM_89_ARLEN),
        .M_AXIMM_89_ARSIZE(M_AXIMM_89_ARSIZE),
        .M_AXIMM_89_ARBURST(M_AXIMM_89_ARBURST),
        .M_AXIMM_89_ARLOCK(M_AXIMM_89_ARLOCK),
        .M_AXIMM_89_ARCACHE(M_AXIMM_89_ARCACHE),
        .M_AXIMM_89_ARPROT(M_AXIMM_89_ARPROT),
        .M_AXIMM_89_ARREGION(M_AXIMM_89_ARREGION),
        .M_AXIMM_89_ARQOS(M_AXIMM_89_ARQOS),
        .M_AXIMM_89_ARVALID(M_AXIMM_89_ARVALID),
        .M_AXIMM_89_ARREADY(M_AXIMM_89_ARREADY),
        .M_AXIMM_89_RDATA(M_AXIMM_89_RDATA),
        .M_AXIMM_89_RRESP(M_AXIMM_89_RRESP),
        .M_AXIMM_89_RLAST(M_AXIMM_89_RLAST),
        .M_AXIMM_89_RVALID(M_AXIMM_89_RVALID),
        .M_AXIMM_89_RREADY(M_AXIMM_89_RREADY),
        .AP_AXIMM_90_AWADDR(AP_AXIMM_90_AWADDR),
        .AP_AXIMM_90_AWLEN(AP_AXIMM_90_AWLEN),
        .AP_AXIMM_90_AWSIZE(AP_AXIMM_90_AWSIZE),
        .AP_AXIMM_90_AWBURST(AP_AXIMM_90_AWBURST),
        .AP_AXIMM_90_AWLOCK(AP_AXIMM_90_AWLOCK),
        .AP_AXIMM_90_AWCACHE(AP_AXIMM_90_AWCACHE),
        .AP_AXIMM_90_AWPROT(AP_AXIMM_90_AWPROT),
        .AP_AXIMM_90_AWREGION(AP_AXIMM_90_AWREGION),
        .AP_AXIMM_90_AWQOS(AP_AXIMM_90_AWQOS),
        .AP_AXIMM_90_AWVALID(AP_AXIMM_90_AWVALID),
        .AP_AXIMM_90_AWREADY(AP_AXIMM_90_AWREADY),
        .AP_AXIMM_90_WDATA(AP_AXIMM_90_WDATA),
        .AP_AXIMM_90_WSTRB(AP_AXIMM_90_WSTRB),
        .AP_AXIMM_90_WLAST(AP_AXIMM_90_WLAST),
        .AP_AXIMM_90_WVALID(AP_AXIMM_90_WVALID),
        .AP_AXIMM_90_WREADY(AP_AXIMM_90_WREADY),
        .AP_AXIMM_90_BRESP(AP_AXIMM_90_BRESP),
        .AP_AXIMM_90_BVALID(AP_AXIMM_90_BVALID),
        .AP_AXIMM_90_BREADY(AP_AXIMM_90_BREADY),
        .AP_AXIMM_90_ARADDR(AP_AXIMM_90_ARADDR),
        .AP_AXIMM_90_ARLEN(AP_AXIMM_90_ARLEN),
        .AP_AXIMM_90_ARSIZE(AP_AXIMM_90_ARSIZE),
        .AP_AXIMM_90_ARBURST(AP_AXIMM_90_ARBURST),
        .AP_AXIMM_90_ARLOCK(AP_AXIMM_90_ARLOCK),
        .AP_AXIMM_90_ARCACHE(AP_AXIMM_90_ARCACHE),
        .AP_AXIMM_90_ARPROT(AP_AXIMM_90_ARPROT),
        .AP_AXIMM_90_ARREGION(AP_AXIMM_90_ARREGION),
        .AP_AXIMM_90_ARQOS(AP_AXIMM_90_ARQOS),
        .AP_AXIMM_90_ARVALID(AP_AXIMM_90_ARVALID),
        .AP_AXIMM_90_ARREADY(AP_AXIMM_90_ARREADY),
        .AP_AXIMM_90_RDATA(AP_AXIMM_90_RDATA),
        .AP_AXIMM_90_RRESP(AP_AXIMM_90_RRESP),
        .AP_AXIMM_90_RLAST(AP_AXIMM_90_RLAST),
        .AP_AXIMM_90_RVALID(AP_AXIMM_90_RVALID),
        .AP_AXIMM_90_RREADY(AP_AXIMM_90_RREADY),
        .M_AXIMM_90_AWADDR(M_AXIMM_90_AWADDR),
        .M_AXIMM_90_AWLEN(M_AXIMM_90_AWLEN),
        .M_AXIMM_90_AWSIZE(M_AXIMM_90_AWSIZE),
        .M_AXIMM_90_AWBURST(M_AXIMM_90_AWBURST),
        .M_AXIMM_90_AWLOCK(M_AXIMM_90_AWLOCK),
        .M_AXIMM_90_AWCACHE(M_AXIMM_90_AWCACHE),
        .M_AXIMM_90_AWPROT(M_AXIMM_90_AWPROT),
        .M_AXIMM_90_AWREGION(M_AXIMM_90_AWREGION),
        .M_AXIMM_90_AWQOS(M_AXIMM_90_AWQOS),
        .M_AXIMM_90_AWVALID(M_AXIMM_90_AWVALID),
        .M_AXIMM_90_AWREADY(M_AXIMM_90_AWREADY),
        .M_AXIMM_90_WDATA(M_AXIMM_90_WDATA),
        .M_AXIMM_90_WSTRB(M_AXIMM_90_WSTRB),
        .M_AXIMM_90_WLAST(M_AXIMM_90_WLAST),
        .M_AXIMM_90_WVALID(M_AXIMM_90_WVALID),
        .M_AXIMM_90_WREADY(M_AXIMM_90_WREADY),
        .M_AXIMM_90_BRESP(M_AXIMM_90_BRESP),
        .M_AXIMM_90_BVALID(M_AXIMM_90_BVALID),
        .M_AXIMM_90_BREADY(M_AXIMM_90_BREADY),
        .M_AXIMM_90_ARADDR(M_AXIMM_90_ARADDR),
        .M_AXIMM_90_ARLEN(M_AXIMM_90_ARLEN),
        .M_AXIMM_90_ARSIZE(M_AXIMM_90_ARSIZE),
        .M_AXIMM_90_ARBURST(M_AXIMM_90_ARBURST),
        .M_AXIMM_90_ARLOCK(M_AXIMM_90_ARLOCK),
        .M_AXIMM_90_ARCACHE(M_AXIMM_90_ARCACHE),
        .M_AXIMM_90_ARPROT(M_AXIMM_90_ARPROT),
        .M_AXIMM_90_ARREGION(M_AXIMM_90_ARREGION),
        .M_AXIMM_90_ARQOS(M_AXIMM_90_ARQOS),
        .M_AXIMM_90_ARVALID(M_AXIMM_90_ARVALID),
        .M_AXIMM_90_ARREADY(M_AXIMM_90_ARREADY),
        .M_AXIMM_90_RDATA(M_AXIMM_90_RDATA),
        .M_AXIMM_90_RRESP(M_AXIMM_90_RRESP),
        .M_AXIMM_90_RLAST(M_AXIMM_90_RLAST),
        .M_AXIMM_90_RVALID(M_AXIMM_90_RVALID),
        .M_AXIMM_90_RREADY(M_AXIMM_90_RREADY),
        .AP_AXIMM_91_AWADDR(AP_AXIMM_91_AWADDR),
        .AP_AXIMM_91_AWLEN(AP_AXIMM_91_AWLEN),
        .AP_AXIMM_91_AWSIZE(AP_AXIMM_91_AWSIZE),
        .AP_AXIMM_91_AWBURST(AP_AXIMM_91_AWBURST),
        .AP_AXIMM_91_AWLOCK(AP_AXIMM_91_AWLOCK),
        .AP_AXIMM_91_AWCACHE(AP_AXIMM_91_AWCACHE),
        .AP_AXIMM_91_AWPROT(AP_AXIMM_91_AWPROT),
        .AP_AXIMM_91_AWREGION(AP_AXIMM_91_AWREGION),
        .AP_AXIMM_91_AWQOS(AP_AXIMM_91_AWQOS),
        .AP_AXIMM_91_AWVALID(AP_AXIMM_91_AWVALID),
        .AP_AXIMM_91_AWREADY(AP_AXIMM_91_AWREADY),
        .AP_AXIMM_91_WDATA(AP_AXIMM_91_WDATA),
        .AP_AXIMM_91_WSTRB(AP_AXIMM_91_WSTRB),
        .AP_AXIMM_91_WLAST(AP_AXIMM_91_WLAST),
        .AP_AXIMM_91_WVALID(AP_AXIMM_91_WVALID),
        .AP_AXIMM_91_WREADY(AP_AXIMM_91_WREADY),
        .AP_AXIMM_91_BRESP(AP_AXIMM_91_BRESP),
        .AP_AXIMM_91_BVALID(AP_AXIMM_91_BVALID),
        .AP_AXIMM_91_BREADY(AP_AXIMM_91_BREADY),
        .AP_AXIMM_91_ARADDR(AP_AXIMM_91_ARADDR),
        .AP_AXIMM_91_ARLEN(AP_AXIMM_91_ARLEN),
        .AP_AXIMM_91_ARSIZE(AP_AXIMM_91_ARSIZE),
        .AP_AXIMM_91_ARBURST(AP_AXIMM_91_ARBURST),
        .AP_AXIMM_91_ARLOCK(AP_AXIMM_91_ARLOCK),
        .AP_AXIMM_91_ARCACHE(AP_AXIMM_91_ARCACHE),
        .AP_AXIMM_91_ARPROT(AP_AXIMM_91_ARPROT),
        .AP_AXIMM_91_ARREGION(AP_AXIMM_91_ARREGION),
        .AP_AXIMM_91_ARQOS(AP_AXIMM_91_ARQOS),
        .AP_AXIMM_91_ARVALID(AP_AXIMM_91_ARVALID),
        .AP_AXIMM_91_ARREADY(AP_AXIMM_91_ARREADY),
        .AP_AXIMM_91_RDATA(AP_AXIMM_91_RDATA),
        .AP_AXIMM_91_RRESP(AP_AXIMM_91_RRESP),
        .AP_AXIMM_91_RLAST(AP_AXIMM_91_RLAST),
        .AP_AXIMM_91_RVALID(AP_AXIMM_91_RVALID),
        .AP_AXIMM_91_RREADY(AP_AXIMM_91_RREADY),
        .M_AXIMM_91_AWADDR(M_AXIMM_91_AWADDR),
        .M_AXIMM_91_AWLEN(M_AXIMM_91_AWLEN),
        .M_AXIMM_91_AWSIZE(M_AXIMM_91_AWSIZE),
        .M_AXIMM_91_AWBURST(M_AXIMM_91_AWBURST),
        .M_AXIMM_91_AWLOCK(M_AXIMM_91_AWLOCK),
        .M_AXIMM_91_AWCACHE(M_AXIMM_91_AWCACHE),
        .M_AXIMM_91_AWPROT(M_AXIMM_91_AWPROT),
        .M_AXIMM_91_AWREGION(M_AXIMM_91_AWREGION),
        .M_AXIMM_91_AWQOS(M_AXIMM_91_AWQOS),
        .M_AXIMM_91_AWVALID(M_AXIMM_91_AWVALID),
        .M_AXIMM_91_AWREADY(M_AXIMM_91_AWREADY),
        .M_AXIMM_91_WDATA(M_AXIMM_91_WDATA),
        .M_AXIMM_91_WSTRB(M_AXIMM_91_WSTRB),
        .M_AXIMM_91_WLAST(M_AXIMM_91_WLAST),
        .M_AXIMM_91_WVALID(M_AXIMM_91_WVALID),
        .M_AXIMM_91_WREADY(M_AXIMM_91_WREADY),
        .M_AXIMM_91_BRESP(M_AXIMM_91_BRESP),
        .M_AXIMM_91_BVALID(M_AXIMM_91_BVALID),
        .M_AXIMM_91_BREADY(M_AXIMM_91_BREADY),
        .M_AXIMM_91_ARADDR(M_AXIMM_91_ARADDR),
        .M_AXIMM_91_ARLEN(M_AXIMM_91_ARLEN),
        .M_AXIMM_91_ARSIZE(M_AXIMM_91_ARSIZE),
        .M_AXIMM_91_ARBURST(M_AXIMM_91_ARBURST),
        .M_AXIMM_91_ARLOCK(M_AXIMM_91_ARLOCK),
        .M_AXIMM_91_ARCACHE(M_AXIMM_91_ARCACHE),
        .M_AXIMM_91_ARPROT(M_AXIMM_91_ARPROT),
        .M_AXIMM_91_ARREGION(M_AXIMM_91_ARREGION),
        .M_AXIMM_91_ARQOS(M_AXIMM_91_ARQOS),
        .M_AXIMM_91_ARVALID(M_AXIMM_91_ARVALID),
        .M_AXIMM_91_ARREADY(M_AXIMM_91_ARREADY),
        .M_AXIMM_91_RDATA(M_AXIMM_91_RDATA),
        .M_AXIMM_91_RRESP(M_AXIMM_91_RRESP),
        .M_AXIMM_91_RLAST(M_AXIMM_91_RLAST),
        .M_AXIMM_91_RVALID(M_AXIMM_91_RVALID),
        .M_AXIMM_91_RREADY(M_AXIMM_91_RREADY),
        .AP_AXIMM_92_AWADDR(AP_AXIMM_92_AWADDR),
        .AP_AXIMM_92_AWLEN(AP_AXIMM_92_AWLEN),
        .AP_AXIMM_92_AWSIZE(AP_AXIMM_92_AWSIZE),
        .AP_AXIMM_92_AWBURST(AP_AXIMM_92_AWBURST),
        .AP_AXIMM_92_AWLOCK(AP_AXIMM_92_AWLOCK),
        .AP_AXIMM_92_AWCACHE(AP_AXIMM_92_AWCACHE),
        .AP_AXIMM_92_AWPROT(AP_AXIMM_92_AWPROT),
        .AP_AXIMM_92_AWREGION(AP_AXIMM_92_AWREGION),
        .AP_AXIMM_92_AWQOS(AP_AXIMM_92_AWQOS),
        .AP_AXIMM_92_AWVALID(AP_AXIMM_92_AWVALID),
        .AP_AXIMM_92_AWREADY(AP_AXIMM_92_AWREADY),
        .AP_AXIMM_92_WDATA(AP_AXIMM_92_WDATA),
        .AP_AXIMM_92_WSTRB(AP_AXIMM_92_WSTRB),
        .AP_AXIMM_92_WLAST(AP_AXIMM_92_WLAST),
        .AP_AXIMM_92_WVALID(AP_AXIMM_92_WVALID),
        .AP_AXIMM_92_WREADY(AP_AXIMM_92_WREADY),
        .AP_AXIMM_92_BRESP(AP_AXIMM_92_BRESP),
        .AP_AXIMM_92_BVALID(AP_AXIMM_92_BVALID),
        .AP_AXIMM_92_BREADY(AP_AXIMM_92_BREADY),
        .AP_AXIMM_92_ARADDR(AP_AXIMM_92_ARADDR),
        .AP_AXIMM_92_ARLEN(AP_AXIMM_92_ARLEN),
        .AP_AXIMM_92_ARSIZE(AP_AXIMM_92_ARSIZE),
        .AP_AXIMM_92_ARBURST(AP_AXIMM_92_ARBURST),
        .AP_AXIMM_92_ARLOCK(AP_AXIMM_92_ARLOCK),
        .AP_AXIMM_92_ARCACHE(AP_AXIMM_92_ARCACHE),
        .AP_AXIMM_92_ARPROT(AP_AXIMM_92_ARPROT),
        .AP_AXIMM_92_ARREGION(AP_AXIMM_92_ARREGION),
        .AP_AXIMM_92_ARQOS(AP_AXIMM_92_ARQOS),
        .AP_AXIMM_92_ARVALID(AP_AXIMM_92_ARVALID),
        .AP_AXIMM_92_ARREADY(AP_AXIMM_92_ARREADY),
        .AP_AXIMM_92_RDATA(AP_AXIMM_92_RDATA),
        .AP_AXIMM_92_RRESP(AP_AXIMM_92_RRESP),
        .AP_AXIMM_92_RLAST(AP_AXIMM_92_RLAST),
        .AP_AXIMM_92_RVALID(AP_AXIMM_92_RVALID),
        .AP_AXIMM_92_RREADY(AP_AXIMM_92_RREADY),
        .M_AXIMM_92_AWADDR(M_AXIMM_92_AWADDR),
        .M_AXIMM_92_AWLEN(M_AXIMM_92_AWLEN),
        .M_AXIMM_92_AWSIZE(M_AXIMM_92_AWSIZE),
        .M_AXIMM_92_AWBURST(M_AXIMM_92_AWBURST),
        .M_AXIMM_92_AWLOCK(M_AXIMM_92_AWLOCK),
        .M_AXIMM_92_AWCACHE(M_AXIMM_92_AWCACHE),
        .M_AXIMM_92_AWPROT(M_AXIMM_92_AWPROT),
        .M_AXIMM_92_AWREGION(M_AXIMM_92_AWREGION),
        .M_AXIMM_92_AWQOS(M_AXIMM_92_AWQOS),
        .M_AXIMM_92_AWVALID(M_AXIMM_92_AWVALID),
        .M_AXIMM_92_AWREADY(M_AXIMM_92_AWREADY),
        .M_AXIMM_92_WDATA(M_AXIMM_92_WDATA),
        .M_AXIMM_92_WSTRB(M_AXIMM_92_WSTRB),
        .M_AXIMM_92_WLAST(M_AXIMM_92_WLAST),
        .M_AXIMM_92_WVALID(M_AXIMM_92_WVALID),
        .M_AXIMM_92_WREADY(M_AXIMM_92_WREADY),
        .M_AXIMM_92_BRESP(M_AXIMM_92_BRESP),
        .M_AXIMM_92_BVALID(M_AXIMM_92_BVALID),
        .M_AXIMM_92_BREADY(M_AXIMM_92_BREADY),
        .M_AXIMM_92_ARADDR(M_AXIMM_92_ARADDR),
        .M_AXIMM_92_ARLEN(M_AXIMM_92_ARLEN),
        .M_AXIMM_92_ARSIZE(M_AXIMM_92_ARSIZE),
        .M_AXIMM_92_ARBURST(M_AXIMM_92_ARBURST),
        .M_AXIMM_92_ARLOCK(M_AXIMM_92_ARLOCK),
        .M_AXIMM_92_ARCACHE(M_AXIMM_92_ARCACHE),
        .M_AXIMM_92_ARPROT(M_AXIMM_92_ARPROT),
        .M_AXIMM_92_ARREGION(M_AXIMM_92_ARREGION),
        .M_AXIMM_92_ARQOS(M_AXIMM_92_ARQOS),
        .M_AXIMM_92_ARVALID(M_AXIMM_92_ARVALID),
        .M_AXIMM_92_ARREADY(M_AXIMM_92_ARREADY),
        .M_AXIMM_92_RDATA(M_AXIMM_92_RDATA),
        .M_AXIMM_92_RRESP(M_AXIMM_92_RRESP),
        .M_AXIMM_92_RLAST(M_AXIMM_92_RLAST),
        .M_AXIMM_92_RVALID(M_AXIMM_92_RVALID),
        .M_AXIMM_92_RREADY(M_AXIMM_92_RREADY),
        .AP_AXIMM_93_AWADDR(AP_AXIMM_93_AWADDR),
        .AP_AXIMM_93_AWLEN(AP_AXIMM_93_AWLEN),
        .AP_AXIMM_93_AWSIZE(AP_AXIMM_93_AWSIZE),
        .AP_AXIMM_93_AWBURST(AP_AXIMM_93_AWBURST),
        .AP_AXIMM_93_AWLOCK(AP_AXIMM_93_AWLOCK),
        .AP_AXIMM_93_AWCACHE(AP_AXIMM_93_AWCACHE),
        .AP_AXIMM_93_AWPROT(AP_AXIMM_93_AWPROT),
        .AP_AXIMM_93_AWREGION(AP_AXIMM_93_AWREGION),
        .AP_AXIMM_93_AWQOS(AP_AXIMM_93_AWQOS),
        .AP_AXIMM_93_AWVALID(AP_AXIMM_93_AWVALID),
        .AP_AXIMM_93_AWREADY(AP_AXIMM_93_AWREADY),
        .AP_AXIMM_93_WDATA(AP_AXIMM_93_WDATA),
        .AP_AXIMM_93_WSTRB(AP_AXIMM_93_WSTRB),
        .AP_AXIMM_93_WLAST(AP_AXIMM_93_WLAST),
        .AP_AXIMM_93_WVALID(AP_AXIMM_93_WVALID),
        .AP_AXIMM_93_WREADY(AP_AXIMM_93_WREADY),
        .AP_AXIMM_93_BRESP(AP_AXIMM_93_BRESP),
        .AP_AXIMM_93_BVALID(AP_AXIMM_93_BVALID),
        .AP_AXIMM_93_BREADY(AP_AXIMM_93_BREADY),
        .AP_AXIMM_93_ARADDR(AP_AXIMM_93_ARADDR),
        .AP_AXIMM_93_ARLEN(AP_AXIMM_93_ARLEN),
        .AP_AXIMM_93_ARSIZE(AP_AXIMM_93_ARSIZE),
        .AP_AXIMM_93_ARBURST(AP_AXIMM_93_ARBURST),
        .AP_AXIMM_93_ARLOCK(AP_AXIMM_93_ARLOCK),
        .AP_AXIMM_93_ARCACHE(AP_AXIMM_93_ARCACHE),
        .AP_AXIMM_93_ARPROT(AP_AXIMM_93_ARPROT),
        .AP_AXIMM_93_ARREGION(AP_AXIMM_93_ARREGION),
        .AP_AXIMM_93_ARQOS(AP_AXIMM_93_ARQOS),
        .AP_AXIMM_93_ARVALID(AP_AXIMM_93_ARVALID),
        .AP_AXIMM_93_ARREADY(AP_AXIMM_93_ARREADY),
        .AP_AXIMM_93_RDATA(AP_AXIMM_93_RDATA),
        .AP_AXIMM_93_RRESP(AP_AXIMM_93_RRESP),
        .AP_AXIMM_93_RLAST(AP_AXIMM_93_RLAST),
        .AP_AXIMM_93_RVALID(AP_AXIMM_93_RVALID),
        .AP_AXIMM_93_RREADY(AP_AXIMM_93_RREADY),
        .M_AXIMM_93_AWADDR(M_AXIMM_93_AWADDR),
        .M_AXIMM_93_AWLEN(M_AXIMM_93_AWLEN),
        .M_AXIMM_93_AWSIZE(M_AXIMM_93_AWSIZE),
        .M_AXIMM_93_AWBURST(M_AXIMM_93_AWBURST),
        .M_AXIMM_93_AWLOCK(M_AXIMM_93_AWLOCK),
        .M_AXIMM_93_AWCACHE(M_AXIMM_93_AWCACHE),
        .M_AXIMM_93_AWPROT(M_AXIMM_93_AWPROT),
        .M_AXIMM_93_AWREGION(M_AXIMM_93_AWREGION),
        .M_AXIMM_93_AWQOS(M_AXIMM_93_AWQOS),
        .M_AXIMM_93_AWVALID(M_AXIMM_93_AWVALID),
        .M_AXIMM_93_AWREADY(M_AXIMM_93_AWREADY),
        .M_AXIMM_93_WDATA(M_AXIMM_93_WDATA),
        .M_AXIMM_93_WSTRB(M_AXIMM_93_WSTRB),
        .M_AXIMM_93_WLAST(M_AXIMM_93_WLAST),
        .M_AXIMM_93_WVALID(M_AXIMM_93_WVALID),
        .M_AXIMM_93_WREADY(M_AXIMM_93_WREADY),
        .M_AXIMM_93_BRESP(M_AXIMM_93_BRESP),
        .M_AXIMM_93_BVALID(M_AXIMM_93_BVALID),
        .M_AXIMM_93_BREADY(M_AXIMM_93_BREADY),
        .M_AXIMM_93_ARADDR(M_AXIMM_93_ARADDR),
        .M_AXIMM_93_ARLEN(M_AXIMM_93_ARLEN),
        .M_AXIMM_93_ARSIZE(M_AXIMM_93_ARSIZE),
        .M_AXIMM_93_ARBURST(M_AXIMM_93_ARBURST),
        .M_AXIMM_93_ARLOCK(M_AXIMM_93_ARLOCK),
        .M_AXIMM_93_ARCACHE(M_AXIMM_93_ARCACHE),
        .M_AXIMM_93_ARPROT(M_AXIMM_93_ARPROT),
        .M_AXIMM_93_ARREGION(M_AXIMM_93_ARREGION),
        .M_AXIMM_93_ARQOS(M_AXIMM_93_ARQOS),
        .M_AXIMM_93_ARVALID(M_AXIMM_93_ARVALID),
        .M_AXIMM_93_ARREADY(M_AXIMM_93_ARREADY),
        .M_AXIMM_93_RDATA(M_AXIMM_93_RDATA),
        .M_AXIMM_93_RRESP(M_AXIMM_93_RRESP),
        .M_AXIMM_93_RLAST(M_AXIMM_93_RLAST),
        .M_AXIMM_93_RVALID(M_AXIMM_93_RVALID),
        .M_AXIMM_93_RREADY(M_AXIMM_93_RREADY),
        .AP_AXIMM_94_AWADDR(AP_AXIMM_94_AWADDR),
        .AP_AXIMM_94_AWLEN(AP_AXIMM_94_AWLEN),
        .AP_AXIMM_94_AWSIZE(AP_AXIMM_94_AWSIZE),
        .AP_AXIMM_94_AWBURST(AP_AXIMM_94_AWBURST),
        .AP_AXIMM_94_AWLOCK(AP_AXIMM_94_AWLOCK),
        .AP_AXIMM_94_AWCACHE(AP_AXIMM_94_AWCACHE),
        .AP_AXIMM_94_AWPROT(AP_AXIMM_94_AWPROT),
        .AP_AXIMM_94_AWREGION(AP_AXIMM_94_AWREGION),
        .AP_AXIMM_94_AWQOS(AP_AXIMM_94_AWQOS),
        .AP_AXIMM_94_AWVALID(AP_AXIMM_94_AWVALID),
        .AP_AXIMM_94_AWREADY(AP_AXIMM_94_AWREADY),
        .AP_AXIMM_94_WDATA(AP_AXIMM_94_WDATA),
        .AP_AXIMM_94_WSTRB(AP_AXIMM_94_WSTRB),
        .AP_AXIMM_94_WLAST(AP_AXIMM_94_WLAST),
        .AP_AXIMM_94_WVALID(AP_AXIMM_94_WVALID),
        .AP_AXIMM_94_WREADY(AP_AXIMM_94_WREADY),
        .AP_AXIMM_94_BRESP(AP_AXIMM_94_BRESP),
        .AP_AXIMM_94_BVALID(AP_AXIMM_94_BVALID),
        .AP_AXIMM_94_BREADY(AP_AXIMM_94_BREADY),
        .AP_AXIMM_94_ARADDR(AP_AXIMM_94_ARADDR),
        .AP_AXIMM_94_ARLEN(AP_AXIMM_94_ARLEN),
        .AP_AXIMM_94_ARSIZE(AP_AXIMM_94_ARSIZE),
        .AP_AXIMM_94_ARBURST(AP_AXIMM_94_ARBURST),
        .AP_AXIMM_94_ARLOCK(AP_AXIMM_94_ARLOCK),
        .AP_AXIMM_94_ARCACHE(AP_AXIMM_94_ARCACHE),
        .AP_AXIMM_94_ARPROT(AP_AXIMM_94_ARPROT),
        .AP_AXIMM_94_ARREGION(AP_AXIMM_94_ARREGION),
        .AP_AXIMM_94_ARQOS(AP_AXIMM_94_ARQOS),
        .AP_AXIMM_94_ARVALID(AP_AXIMM_94_ARVALID),
        .AP_AXIMM_94_ARREADY(AP_AXIMM_94_ARREADY),
        .AP_AXIMM_94_RDATA(AP_AXIMM_94_RDATA),
        .AP_AXIMM_94_RRESP(AP_AXIMM_94_RRESP),
        .AP_AXIMM_94_RLAST(AP_AXIMM_94_RLAST),
        .AP_AXIMM_94_RVALID(AP_AXIMM_94_RVALID),
        .AP_AXIMM_94_RREADY(AP_AXIMM_94_RREADY),
        .M_AXIMM_94_AWADDR(M_AXIMM_94_AWADDR),
        .M_AXIMM_94_AWLEN(M_AXIMM_94_AWLEN),
        .M_AXIMM_94_AWSIZE(M_AXIMM_94_AWSIZE),
        .M_AXIMM_94_AWBURST(M_AXIMM_94_AWBURST),
        .M_AXIMM_94_AWLOCK(M_AXIMM_94_AWLOCK),
        .M_AXIMM_94_AWCACHE(M_AXIMM_94_AWCACHE),
        .M_AXIMM_94_AWPROT(M_AXIMM_94_AWPROT),
        .M_AXIMM_94_AWREGION(M_AXIMM_94_AWREGION),
        .M_AXIMM_94_AWQOS(M_AXIMM_94_AWQOS),
        .M_AXIMM_94_AWVALID(M_AXIMM_94_AWVALID),
        .M_AXIMM_94_AWREADY(M_AXIMM_94_AWREADY),
        .M_AXIMM_94_WDATA(M_AXIMM_94_WDATA),
        .M_AXIMM_94_WSTRB(M_AXIMM_94_WSTRB),
        .M_AXIMM_94_WLAST(M_AXIMM_94_WLAST),
        .M_AXIMM_94_WVALID(M_AXIMM_94_WVALID),
        .M_AXIMM_94_WREADY(M_AXIMM_94_WREADY),
        .M_AXIMM_94_BRESP(M_AXIMM_94_BRESP),
        .M_AXIMM_94_BVALID(M_AXIMM_94_BVALID),
        .M_AXIMM_94_BREADY(M_AXIMM_94_BREADY),
        .M_AXIMM_94_ARADDR(M_AXIMM_94_ARADDR),
        .M_AXIMM_94_ARLEN(M_AXIMM_94_ARLEN),
        .M_AXIMM_94_ARSIZE(M_AXIMM_94_ARSIZE),
        .M_AXIMM_94_ARBURST(M_AXIMM_94_ARBURST),
        .M_AXIMM_94_ARLOCK(M_AXIMM_94_ARLOCK),
        .M_AXIMM_94_ARCACHE(M_AXIMM_94_ARCACHE),
        .M_AXIMM_94_ARPROT(M_AXIMM_94_ARPROT),
        .M_AXIMM_94_ARREGION(M_AXIMM_94_ARREGION),
        .M_AXIMM_94_ARQOS(M_AXIMM_94_ARQOS),
        .M_AXIMM_94_ARVALID(M_AXIMM_94_ARVALID),
        .M_AXIMM_94_ARREADY(M_AXIMM_94_ARREADY),
        .M_AXIMM_94_RDATA(M_AXIMM_94_RDATA),
        .M_AXIMM_94_RRESP(M_AXIMM_94_RRESP),
        .M_AXIMM_94_RLAST(M_AXIMM_94_RLAST),
        .M_AXIMM_94_RVALID(M_AXIMM_94_RVALID),
        .M_AXIMM_94_RREADY(M_AXIMM_94_RREADY),
        .AP_AXIMM_95_AWADDR(AP_AXIMM_95_AWADDR),
        .AP_AXIMM_95_AWLEN(AP_AXIMM_95_AWLEN),
        .AP_AXIMM_95_AWSIZE(AP_AXIMM_95_AWSIZE),
        .AP_AXIMM_95_AWBURST(AP_AXIMM_95_AWBURST),
        .AP_AXIMM_95_AWLOCK(AP_AXIMM_95_AWLOCK),
        .AP_AXIMM_95_AWCACHE(AP_AXIMM_95_AWCACHE),
        .AP_AXIMM_95_AWPROT(AP_AXIMM_95_AWPROT),
        .AP_AXIMM_95_AWREGION(AP_AXIMM_95_AWREGION),
        .AP_AXIMM_95_AWQOS(AP_AXIMM_95_AWQOS),
        .AP_AXIMM_95_AWVALID(AP_AXIMM_95_AWVALID),
        .AP_AXIMM_95_AWREADY(AP_AXIMM_95_AWREADY),
        .AP_AXIMM_95_WDATA(AP_AXIMM_95_WDATA),
        .AP_AXIMM_95_WSTRB(AP_AXIMM_95_WSTRB),
        .AP_AXIMM_95_WLAST(AP_AXIMM_95_WLAST),
        .AP_AXIMM_95_WVALID(AP_AXIMM_95_WVALID),
        .AP_AXIMM_95_WREADY(AP_AXIMM_95_WREADY),
        .AP_AXIMM_95_BRESP(AP_AXIMM_95_BRESP),
        .AP_AXIMM_95_BVALID(AP_AXIMM_95_BVALID),
        .AP_AXIMM_95_BREADY(AP_AXIMM_95_BREADY),
        .AP_AXIMM_95_ARADDR(AP_AXIMM_95_ARADDR),
        .AP_AXIMM_95_ARLEN(AP_AXIMM_95_ARLEN),
        .AP_AXIMM_95_ARSIZE(AP_AXIMM_95_ARSIZE),
        .AP_AXIMM_95_ARBURST(AP_AXIMM_95_ARBURST),
        .AP_AXIMM_95_ARLOCK(AP_AXIMM_95_ARLOCK),
        .AP_AXIMM_95_ARCACHE(AP_AXIMM_95_ARCACHE),
        .AP_AXIMM_95_ARPROT(AP_AXIMM_95_ARPROT),
        .AP_AXIMM_95_ARREGION(AP_AXIMM_95_ARREGION),
        .AP_AXIMM_95_ARQOS(AP_AXIMM_95_ARQOS),
        .AP_AXIMM_95_ARVALID(AP_AXIMM_95_ARVALID),
        .AP_AXIMM_95_ARREADY(AP_AXIMM_95_ARREADY),
        .AP_AXIMM_95_RDATA(AP_AXIMM_95_RDATA),
        .AP_AXIMM_95_RRESP(AP_AXIMM_95_RRESP),
        .AP_AXIMM_95_RLAST(AP_AXIMM_95_RLAST),
        .AP_AXIMM_95_RVALID(AP_AXIMM_95_RVALID),
        .AP_AXIMM_95_RREADY(AP_AXIMM_95_RREADY),
        .M_AXIMM_95_AWADDR(M_AXIMM_95_AWADDR),
        .M_AXIMM_95_AWLEN(M_AXIMM_95_AWLEN),
        .M_AXIMM_95_AWSIZE(M_AXIMM_95_AWSIZE),
        .M_AXIMM_95_AWBURST(M_AXIMM_95_AWBURST),
        .M_AXIMM_95_AWLOCK(M_AXIMM_95_AWLOCK),
        .M_AXIMM_95_AWCACHE(M_AXIMM_95_AWCACHE),
        .M_AXIMM_95_AWPROT(M_AXIMM_95_AWPROT),
        .M_AXIMM_95_AWREGION(M_AXIMM_95_AWREGION),
        .M_AXIMM_95_AWQOS(M_AXIMM_95_AWQOS),
        .M_AXIMM_95_AWVALID(M_AXIMM_95_AWVALID),
        .M_AXIMM_95_AWREADY(M_AXIMM_95_AWREADY),
        .M_AXIMM_95_WDATA(M_AXIMM_95_WDATA),
        .M_AXIMM_95_WSTRB(M_AXIMM_95_WSTRB),
        .M_AXIMM_95_WLAST(M_AXIMM_95_WLAST),
        .M_AXIMM_95_WVALID(M_AXIMM_95_WVALID),
        .M_AXIMM_95_WREADY(M_AXIMM_95_WREADY),
        .M_AXIMM_95_BRESP(M_AXIMM_95_BRESP),
        .M_AXIMM_95_BVALID(M_AXIMM_95_BVALID),
        .M_AXIMM_95_BREADY(M_AXIMM_95_BREADY),
        .M_AXIMM_95_ARADDR(M_AXIMM_95_ARADDR),
        .M_AXIMM_95_ARLEN(M_AXIMM_95_ARLEN),
        .M_AXIMM_95_ARSIZE(M_AXIMM_95_ARSIZE),
        .M_AXIMM_95_ARBURST(M_AXIMM_95_ARBURST),
        .M_AXIMM_95_ARLOCK(M_AXIMM_95_ARLOCK),
        .M_AXIMM_95_ARCACHE(M_AXIMM_95_ARCACHE),
        .M_AXIMM_95_ARPROT(M_AXIMM_95_ARPROT),
        .M_AXIMM_95_ARREGION(M_AXIMM_95_ARREGION),
        .M_AXIMM_95_ARQOS(M_AXIMM_95_ARQOS),
        .M_AXIMM_95_ARVALID(M_AXIMM_95_ARVALID),
        .M_AXIMM_95_ARREADY(M_AXIMM_95_ARREADY),
        .M_AXIMM_95_RDATA(M_AXIMM_95_RDATA),
        .M_AXIMM_95_RRESP(M_AXIMM_95_RRESP),
        .M_AXIMM_95_RLAST(M_AXIMM_95_RLAST),
        .M_AXIMM_95_RVALID(M_AXIMM_95_RVALID),
        .M_AXIMM_95_RREADY(M_AXIMM_95_RREADY),
        .AP_AXIMM_96_AWADDR(AP_AXIMM_96_AWADDR),
        .AP_AXIMM_96_AWLEN(AP_AXIMM_96_AWLEN),
        .AP_AXIMM_96_AWSIZE(AP_AXIMM_96_AWSIZE),
        .AP_AXIMM_96_AWBURST(AP_AXIMM_96_AWBURST),
        .AP_AXIMM_96_AWLOCK(AP_AXIMM_96_AWLOCK),
        .AP_AXIMM_96_AWCACHE(AP_AXIMM_96_AWCACHE),
        .AP_AXIMM_96_AWPROT(AP_AXIMM_96_AWPROT),
        .AP_AXIMM_96_AWREGION(AP_AXIMM_96_AWREGION),
        .AP_AXIMM_96_AWQOS(AP_AXIMM_96_AWQOS),
        .AP_AXIMM_96_AWVALID(AP_AXIMM_96_AWVALID),
        .AP_AXIMM_96_AWREADY(AP_AXIMM_96_AWREADY),
        .AP_AXIMM_96_WDATA(AP_AXIMM_96_WDATA),
        .AP_AXIMM_96_WSTRB(AP_AXIMM_96_WSTRB),
        .AP_AXIMM_96_WLAST(AP_AXIMM_96_WLAST),
        .AP_AXIMM_96_WVALID(AP_AXIMM_96_WVALID),
        .AP_AXIMM_96_WREADY(AP_AXIMM_96_WREADY),
        .AP_AXIMM_96_BRESP(AP_AXIMM_96_BRESP),
        .AP_AXIMM_96_BVALID(AP_AXIMM_96_BVALID),
        .AP_AXIMM_96_BREADY(AP_AXIMM_96_BREADY),
        .AP_AXIMM_96_ARADDR(AP_AXIMM_96_ARADDR),
        .AP_AXIMM_96_ARLEN(AP_AXIMM_96_ARLEN),
        .AP_AXIMM_96_ARSIZE(AP_AXIMM_96_ARSIZE),
        .AP_AXIMM_96_ARBURST(AP_AXIMM_96_ARBURST),
        .AP_AXIMM_96_ARLOCK(AP_AXIMM_96_ARLOCK),
        .AP_AXIMM_96_ARCACHE(AP_AXIMM_96_ARCACHE),
        .AP_AXIMM_96_ARPROT(AP_AXIMM_96_ARPROT),
        .AP_AXIMM_96_ARREGION(AP_AXIMM_96_ARREGION),
        .AP_AXIMM_96_ARQOS(AP_AXIMM_96_ARQOS),
        .AP_AXIMM_96_ARVALID(AP_AXIMM_96_ARVALID),
        .AP_AXIMM_96_ARREADY(AP_AXIMM_96_ARREADY),
        .AP_AXIMM_96_RDATA(AP_AXIMM_96_RDATA),
        .AP_AXIMM_96_RRESP(AP_AXIMM_96_RRESP),
        .AP_AXIMM_96_RLAST(AP_AXIMM_96_RLAST),
        .AP_AXIMM_96_RVALID(AP_AXIMM_96_RVALID),
        .AP_AXIMM_96_RREADY(AP_AXIMM_96_RREADY),
        .M_AXIMM_96_AWADDR(M_AXIMM_96_AWADDR),
        .M_AXIMM_96_AWLEN(M_AXIMM_96_AWLEN),
        .M_AXIMM_96_AWSIZE(M_AXIMM_96_AWSIZE),
        .M_AXIMM_96_AWBURST(M_AXIMM_96_AWBURST),
        .M_AXIMM_96_AWLOCK(M_AXIMM_96_AWLOCK),
        .M_AXIMM_96_AWCACHE(M_AXIMM_96_AWCACHE),
        .M_AXIMM_96_AWPROT(M_AXIMM_96_AWPROT),
        .M_AXIMM_96_AWREGION(M_AXIMM_96_AWREGION),
        .M_AXIMM_96_AWQOS(M_AXIMM_96_AWQOS),
        .M_AXIMM_96_AWVALID(M_AXIMM_96_AWVALID),
        .M_AXIMM_96_AWREADY(M_AXIMM_96_AWREADY),
        .M_AXIMM_96_WDATA(M_AXIMM_96_WDATA),
        .M_AXIMM_96_WSTRB(M_AXIMM_96_WSTRB),
        .M_AXIMM_96_WLAST(M_AXIMM_96_WLAST),
        .M_AXIMM_96_WVALID(M_AXIMM_96_WVALID),
        .M_AXIMM_96_WREADY(M_AXIMM_96_WREADY),
        .M_AXIMM_96_BRESP(M_AXIMM_96_BRESP),
        .M_AXIMM_96_BVALID(M_AXIMM_96_BVALID),
        .M_AXIMM_96_BREADY(M_AXIMM_96_BREADY),
        .M_AXIMM_96_ARADDR(M_AXIMM_96_ARADDR),
        .M_AXIMM_96_ARLEN(M_AXIMM_96_ARLEN),
        .M_AXIMM_96_ARSIZE(M_AXIMM_96_ARSIZE),
        .M_AXIMM_96_ARBURST(M_AXIMM_96_ARBURST),
        .M_AXIMM_96_ARLOCK(M_AXIMM_96_ARLOCK),
        .M_AXIMM_96_ARCACHE(M_AXIMM_96_ARCACHE),
        .M_AXIMM_96_ARPROT(M_AXIMM_96_ARPROT),
        .M_AXIMM_96_ARREGION(M_AXIMM_96_ARREGION),
        .M_AXIMM_96_ARQOS(M_AXIMM_96_ARQOS),
        .M_AXIMM_96_ARVALID(M_AXIMM_96_ARVALID),
        .M_AXIMM_96_ARREADY(M_AXIMM_96_ARREADY),
        .M_AXIMM_96_RDATA(M_AXIMM_96_RDATA),
        .M_AXIMM_96_RRESP(M_AXIMM_96_RRESP),
        .M_AXIMM_96_RLAST(M_AXIMM_96_RLAST),
        .M_AXIMM_96_RVALID(M_AXIMM_96_RVALID),
        .M_AXIMM_96_RREADY(M_AXIMM_96_RREADY),
        .AP_AXIMM_97_AWADDR(AP_AXIMM_97_AWADDR),
        .AP_AXIMM_97_AWLEN(AP_AXIMM_97_AWLEN),
        .AP_AXIMM_97_AWSIZE(AP_AXIMM_97_AWSIZE),
        .AP_AXIMM_97_AWBURST(AP_AXIMM_97_AWBURST),
        .AP_AXIMM_97_AWLOCK(AP_AXIMM_97_AWLOCK),
        .AP_AXIMM_97_AWCACHE(AP_AXIMM_97_AWCACHE),
        .AP_AXIMM_97_AWPROT(AP_AXIMM_97_AWPROT),
        .AP_AXIMM_97_AWREGION(AP_AXIMM_97_AWREGION),
        .AP_AXIMM_97_AWQOS(AP_AXIMM_97_AWQOS),
        .AP_AXIMM_97_AWVALID(AP_AXIMM_97_AWVALID),
        .AP_AXIMM_97_AWREADY(AP_AXIMM_97_AWREADY),
        .AP_AXIMM_97_WDATA(AP_AXIMM_97_WDATA),
        .AP_AXIMM_97_WSTRB(AP_AXIMM_97_WSTRB),
        .AP_AXIMM_97_WLAST(AP_AXIMM_97_WLAST),
        .AP_AXIMM_97_WVALID(AP_AXIMM_97_WVALID),
        .AP_AXIMM_97_WREADY(AP_AXIMM_97_WREADY),
        .AP_AXIMM_97_BRESP(AP_AXIMM_97_BRESP),
        .AP_AXIMM_97_BVALID(AP_AXIMM_97_BVALID),
        .AP_AXIMM_97_BREADY(AP_AXIMM_97_BREADY),
        .AP_AXIMM_97_ARADDR(AP_AXIMM_97_ARADDR),
        .AP_AXIMM_97_ARLEN(AP_AXIMM_97_ARLEN),
        .AP_AXIMM_97_ARSIZE(AP_AXIMM_97_ARSIZE),
        .AP_AXIMM_97_ARBURST(AP_AXIMM_97_ARBURST),
        .AP_AXIMM_97_ARLOCK(AP_AXIMM_97_ARLOCK),
        .AP_AXIMM_97_ARCACHE(AP_AXIMM_97_ARCACHE),
        .AP_AXIMM_97_ARPROT(AP_AXIMM_97_ARPROT),
        .AP_AXIMM_97_ARREGION(AP_AXIMM_97_ARREGION),
        .AP_AXIMM_97_ARQOS(AP_AXIMM_97_ARQOS),
        .AP_AXIMM_97_ARVALID(AP_AXIMM_97_ARVALID),
        .AP_AXIMM_97_ARREADY(AP_AXIMM_97_ARREADY),
        .AP_AXIMM_97_RDATA(AP_AXIMM_97_RDATA),
        .AP_AXIMM_97_RRESP(AP_AXIMM_97_RRESP),
        .AP_AXIMM_97_RLAST(AP_AXIMM_97_RLAST),
        .AP_AXIMM_97_RVALID(AP_AXIMM_97_RVALID),
        .AP_AXIMM_97_RREADY(AP_AXIMM_97_RREADY),
        .M_AXIMM_97_AWADDR(M_AXIMM_97_AWADDR),
        .M_AXIMM_97_AWLEN(M_AXIMM_97_AWLEN),
        .M_AXIMM_97_AWSIZE(M_AXIMM_97_AWSIZE),
        .M_AXIMM_97_AWBURST(M_AXIMM_97_AWBURST),
        .M_AXIMM_97_AWLOCK(M_AXIMM_97_AWLOCK),
        .M_AXIMM_97_AWCACHE(M_AXIMM_97_AWCACHE),
        .M_AXIMM_97_AWPROT(M_AXIMM_97_AWPROT),
        .M_AXIMM_97_AWREGION(M_AXIMM_97_AWREGION),
        .M_AXIMM_97_AWQOS(M_AXIMM_97_AWQOS),
        .M_AXIMM_97_AWVALID(M_AXIMM_97_AWVALID),
        .M_AXIMM_97_AWREADY(M_AXIMM_97_AWREADY),
        .M_AXIMM_97_WDATA(M_AXIMM_97_WDATA),
        .M_AXIMM_97_WSTRB(M_AXIMM_97_WSTRB),
        .M_AXIMM_97_WLAST(M_AXIMM_97_WLAST),
        .M_AXIMM_97_WVALID(M_AXIMM_97_WVALID),
        .M_AXIMM_97_WREADY(M_AXIMM_97_WREADY),
        .M_AXIMM_97_BRESP(M_AXIMM_97_BRESP),
        .M_AXIMM_97_BVALID(M_AXIMM_97_BVALID),
        .M_AXIMM_97_BREADY(M_AXIMM_97_BREADY),
        .M_AXIMM_97_ARADDR(M_AXIMM_97_ARADDR),
        .M_AXIMM_97_ARLEN(M_AXIMM_97_ARLEN),
        .M_AXIMM_97_ARSIZE(M_AXIMM_97_ARSIZE),
        .M_AXIMM_97_ARBURST(M_AXIMM_97_ARBURST),
        .M_AXIMM_97_ARLOCK(M_AXIMM_97_ARLOCK),
        .M_AXIMM_97_ARCACHE(M_AXIMM_97_ARCACHE),
        .M_AXIMM_97_ARPROT(M_AXIMM_97_ARPROT),
        .M_AXIMM_97_ARREGION(M_AXIMM_97_ARREGION),
        .M_AXIMM_97_ARQOS(M_AXIMM_97_ARQOS),
        .M_AXIMM_97_ARVALID(M_AXIMM_97_ARVALID),
        .M_AXIMM_97_ARREADY(M_AXIMM_97_ARREADY),
        .M_AXIMM_97_RDATA(M_AXIMM_97_RDATA),
        .M_AXIMM_97_RRESP(M_AXIMM_97_RRESP),
        .M_AXIMM_97_RLAST(M_AXIMM_97_RLAST),
        .M_AXIMM_97_RVALID(M_AXIMM_97_RVALID),
        .M_AXIMM_97_RREADY(M_AXIMM_97_RREADY),
        .AP_AXIMM_98_AWADDR(AP_AXIMM_98_AWADDR),
        .AP_AXIMM_98_AWLEN(AP_AXIMM_98_AWLEN),
        .AP_AXIMM_98_AWSIZE(AP_AXIMM_98_AWSIZE),
        .AP_AXIMM_98_AWBURST(AP_AXIMM_98_AWBURST),
        .AP_AXIMM_98_AWLOCK(AP_AXIMM_98_AWLOCK),
        .AP_AXIMM_98_AWCACHE(AP_AXIMM_98_AWCACHE),
        .AP_AXIMM_98_AWPROT(AP_AXIMM_98_AWPROT),
        .AP_AXIMM_98_AWREGION(AP_AXIMM_98_AWREGION),
        .AP_AXIMM_98_AWQOS(AP_AXIMM_98_AWQOS),
        .AP_AXIMM_98_AWVALID(AP_AXIMM_98_AWVALID),
        .AP_AXIMM_98_AWREADY(AP_AXIMM_98_AWREADY),
        .AP_AXIMM_98_WDATA(AP_AXIMM_98_WDATA),
        .AP_AXIMM_98_WSTRB(AP_AXIMM_98_WSTRB),
        .AP_AXIMM_98_WLAST(AP_AXIMM_98_WLAST),
        .AP_AXIMM_98_WVALID(AP_AXIMM_98_WVALID),
        .AP_AXIMM_98_WREADY(AP_AXIMM_98_WREADY),
        .AP_AXIMM_98_BRESP(AP_AXIMM_98_BRESP),
        .AP_AXIMM_98_BVALID(AP_AXIMM_98_BVALID),
        .AP_AXIMM_98_BREADY(AP_AXIMM_98_BREADY),
        .AP_AXIMM_98_ARADDR(AP_AXIMM_98_ARADDR),
        .AP_AXIMM_98_ARLEN(AP_AXIMM_98_ARLEN),
        .AP_AXIMM_98_ARSIZE(AP_AXIMM_98_ARSIZE),
        .AP_AXIMM_98_ARBURST(AP_AXIMM_98_ARBURST),
        .AP_AXIMM_98_ARLOCK(AP_AXIMM_98_ARLOCK),
        .AP_AXIMM_98_ARCACHE(AP_AXIMM_98_ARCACHE),
        .AP_AXIMM_98_ARPROT(AP_AXIMM_98_ARPROT),
        .AP_AXIMM_98_ARREGION(AP_AXIMM_98_ARREGION),
        .AP_AXIMM_98_ARQOS(AP_AXIMM_98_ARQOS),
        .AP_AXIMM_98_ARVALID(AP_AXIMM_98_ARVALID),
        .AP_AXIMM_98_ARREADY(AP_AXIMM_98_ARREADY),
        .AP_AXIMM_98_RDATA(AP_AXIMM_98_RDATA),
        .AP_AXIMM_98_RRESP(AP_AXIMM_98_RRESP),
        .AP_AXIMM_98_RLAST(AP_AXIMM_98_RLAST),
        .AP_AXIMM_98_RVALID(AP_AXIMM_98_RVALID),
        .AP_AXIMM_98_RREADY(AP_AXIMM_98_RREADY),
        .M_AXIMM_98_AWADDR(M_AXIMM_98_AWADDR),
        .M_AXIMM_98_AWLEN(M_AXIMM_98_AWLEN),
        .M_AXIMM_98_AWSIZE(M_AXIMM_98_AWSIZE),
        .M_AXIMM_98_AWBURST(M_AXIMM_98_AWBURST),
        .M_AXIMM_98_AWLOCK(M_AXIMM_98_AWLOCK),
        .M_AXIMM_98_AWCACHE(M_AXIMM_98_AWCACHE),
        .M_AXIMM_98_AWPROT(M_AXIMM_98_AWPROT),
        .M_AXIMM_98_AWREGION(M_AXIMM_98_AWREGION),
        .M_AXIMM_98_AWQOS(M_AXIMM_98_AWQOS),
        .M_AXIMM_98_AWVALID(M_AXIMM_98_AWVALID),
        .M_AXIMM_98_AWREADY(M_AXIMM_98_AWREADY),
        .M_AXIMM_98_WDATA(M_AXIMM_98_WDATA),
        .M_AXIMM_98_WSTRB(M_AXIMM_98_WSTRB),
        .M_AXIMM_98_WLAST(M_AXIMM_98_WLAST),
        .M_AXIMM_98_WVALID(M_AXIMM_98_WVALID),
        .M_AXIMM_98_WREADY(M_AXIMM_98_WREADY),
        .M_AXIMM_98_BRESP(M_AXIMM_98_BRESP),
        .M_AXIMM_98_BVALID(M_AXIMM_98_BVALID),
        .M_AXIMM_98_BREADY(M_AXIMM_98_BREADY),
        .M_AXIMM_98_ARADDR(M_AXIMM_98_ARADDR),
        .M_AXIMM_98_ARLEN(M_AXIMM_98_ARLEN),
        .M_AXIMM_98_ARSIZE(M_AXIMM_98_ARSIZE),
        .M_AXIMM_98_ARBURST(M_AXIMM_98_ARBURST),
        .M_AXIMM_98_ARLOCK(M_AXIMM_98_ARLOCK),
        .M_AXIMM_98_ARCACHE(M_AXIMM_98_ARCACHE),
        .M_AXIMM_98_ARPROT(M_AXIMM_98_ARPROT),
        .M_AXIMM_98_ARREGION(M_AXIMM_98_ARREGION),
        .M_AXIMM_98_ARQOS(M_AXIMM_98_ARQOS),
        .M_AXIMM_98_ARVALID(M_AXIMM_98_ARVALID),
        .M_AXIMM_98_ARREADY(M_AXIMM_98_ARREADY),
        .M_AXIMM_98_RDATA(M_AXIMM_98_RDATA),
        .M_AXIMM_98_RRESP(M_AXIMM_98_RRESP),
        .M_AXIMM_98_RLAST(M_AXIMM_98_RLAST),
        .M_AXIMM_98_RVALID(M_AXIMM_98_RVALID),
        .M_AXIMM_98_RREADY(M_AXIMM_98_RREADY),
        .AP_AXIMM_99_AWADDR(AP_AXIMM_99_AWADDR),
        .AP_AXIMM_99_AWLEN(AP_AXIMM_99_AWLEN),
        .AP_AXIMM_99_AWSIZE(AP_AXIMM_99_AWSIZE),
        .AP_AXIMM_99_AWBURST(AP_AXIMM_99_AWBURST),
        .AP_AXIMM_99_AWLOCK(AP_AXIMM_99_AWLOCK),
        .AP_AXIMM_99_AWCACHE(AP_AXIMM_99_AWCACHE),
        .AP_AXIMM_99_AWPROT(AP_AXIMM_99_AWPROT),
        .AP_AXIMM_99_AWREGION(AP_AXIMM_99_AWREGION),
        .AP_AXIMM_99_AWQOS(AP_AXIMM_99_AWQOS),
        .AP_AXIMM_99_AWVALID(AP_AXIMM_99_AWVALID),
        .AP_AXIMM_99_AWREADY(AP_AXIMM_99_AWREADY),
        .AP_AXIMM_99_WDATA(AP_AXIMM_99_WDATA),
        .AP_AXIMM_99_WSTRB(AP_AXIMM_99_WSTRB),
        .AP_AXIMM_99_WLAST(AP_AXIMM_99_WLAST),
        .AP_AXIMM_99_WVALID(AP_AXIMM_99_WVALID),
        .AP_AXIMM_99_WREADY(AP_AXIMM_99_WREADY),
        .AP_AXIMM_99_BRESP(AP_AXIMM_99_BRESP),
        .AP_AXIMM_99_BVALID(AP_AXIMM_99_BVALID),
        .AP_AXIMM_99_BREADY(AP_AXIMM_99_BREADY),
        .AP_AXIMM_99_ARADDR(AP_AXIMM_99_ARADDR),
        .AP_AXIMM_99_ARLEN(AP_AXIMM_99_ARLEN),
        .AP_AXIMM_99_ARSIZE(AP_AXIMM_99_ARSIZE),
        .AP_AXIMM_99_ARBURST(AP_AXIMM_99_ARBURST),
        .AP_AXIMM_99_ARLOCK(AP_AXIMM_99_ARLOCK),
        .AP_AXIMM_99_ARCACHE(AP_AXIMM_99_ARCACHE),
        .AP_AXIMM_99_ARPROT(AP_AXIMM_99_ARPROT),
        .AP_AXIMM_99_ARREGION(AP_AXIMM_99_ARREGION),
        .AP_AXIMM_99_ARQOS(AP_AXIMM_99_ARQOS),
        .AP_AXIMM_99_ARVALID(AP_AXIMM_99_ARVALID),
        .AP_AXIMM_99_ARREADY(AP_AXIMM_99_ARREADY),
        .AP_AXIMM_99_RDATA(AP_AXIMM_99_RDATA),
        .AP_AXIMM_99_RRESP(AP_AXIMM_99_RRESP),
        .AP_AXIMM_99_RLAST(AP_AXIMM_99_RLAST),
        .AP_AXIMM_99_RVALID(AP_AXIMM_99_RVALID),
        .AP_AXIMM_99_RREADY(AP_AXIMM_99_RREADY),
        .M_AXIMM_99_AWADDR(M_AXIMM_99_AWADDR),
        .M_AXIMM_99_AWLEN(M_AXIMM_99_AWLEN),
        .M_AXIMM_99_AWSIZE(M_AXIMM_99_AWSIZE),
        .M_AXIMM_99_AWBURST(M_AXIMM_99_AWBURST),
        .M_AXIMM_99_AWLOCK(M_AXIMM_99_AWLOCK),
        .M_AXIMM_99_AWCACHE(M_AXIMM_99_AWCACHE),
        .M_AXIMM_99_AWPROT(M_AXIMM_99_AWPROT),
        .M_AXIMM_99_AWREGION(M_AXIMM_99_AWREGION),
        .M_AXIMM_99_AWQOS(M_AXIMM_99_AWQOS),
        .M_AXIMM_99_AWVALID(M_AXIMM_99_AWVALID),
        .M_AXIMM_99_AWREADY(M_AXIMM_99_AWREADY),
        .M_AXIMM_99_WDATA(M_AXIMM_99_WDATA),
        .M_AXIMM_99_WSTRB(M_AXIMM_99_WSTRB),
        .M_AXIMM_99_WLAST(M_AXIMM_99_WLAST),
        .M_AXIMM_99_WVALID(M_AXIMM_99_WVALID),
        .M_AXIMM_99_WREADY(M_AXIMM_99_WREADY),
        .M_AXIMM_99_BRESP(M_AXIMM_99_BRESP),
        .M_AXIMM_99_BVALID(M_AXIMM_99_BVALID),
        .M_AXIMM_99_BREADY(M_AXIMM_99_BREADY),
        .M_AXIMM_99_ARADDR(M_AXIMM_99_ARADDR),
        .M_AXIMM_99_ARLEN(M_AXIMM_99_ARLEN),
        .M_AXIMM_99_ARSIZE(M_AXIMM_99_ARSIZE),
        .M_AXIMM_99_ARBURST(M_AXIMM_99_ARBURST),
        .M_AXIMM_99_ARLOCK(M_AXIMM_99_ARLOCK),
        .M_AXIMM_99_ARCACHE(M_AXIMM_99_ARCACHE),
        .M_AXIMM_99_ARPROT(M_AXIMM_99_ARPROT),
        .M_AXIMM_99_ARREGION(M_AXIMM_99_ARREGION),
        .M_AXIMM_99_ARQOS(M_AXIMM_99_ARQOS),
        .M_AXIMM_99_ARVALID(M_AXIMM_99_ARVALID),
        .M_AXIMM_99_ARREADY(M_AXIMM_99_ARREADY),
        .M_AXIMM_99_RDATA(M_AXIMM_99_RDATA),
        .M_AXIMM_99_RRESP(M_AXIMM_99_RRESP),
        .M_AXIMM_99_RLAST(M_AXIMM_99_RLAST),
        .M_AXIMM_99_RVALID(M_AXIMM_99_RVALID),
        .M_AXIMM_99_RREADY(M_AXIMM_99_RREADY),
        .AP_AXIMM_100_AWADDR(AP_AXIMM_100_AWADDR),
        .AP_AXIMM_100_AWLEN(AP_AXIMM_100_AWLEN),
        .AP_AXIMM_100_AWSIZE(AP_AXIMM_100_AWSIZE),
        .AP_AXIMM_100_AWBURST(AP_AXIMM_100_AWBURST),
        .AP_AXIMM_100_AWLOCK(AP_AXIMM_100_AWLOCK),
        .AP_AXIMM_100_AWCACHE(AP_AXIMM_100_AWCACHE),
        .AP_AXIMM_100_AWPROT(AP_AXIMM_100_AWPROT),
        .AP_AXIMM_100_AWREGION(AP_AXIMM_100_AWREGION),
        .AP_AXIMM_100_AWQOS(AP_AXIMM_100_AWQOS),
        .AP_AXIMM_100_AWVALID(AP_AXIMM_100_AWVALID),
        .AP_AXIMM_100_AWREADY(AP_AXIMM_100_AWREADY),
        .AP_AXIMM_100_WDATA(AP_AXIMM_100_WDATA),
        .AP_AXIMM_100_WSTRB(AP_AXIMM_100_WSTRB),
        .AP_AXIMM_100_WLAST(AP_AXIMM_100_WLAST),
        .AP_AXIMM_100_WVALID(AP_AXIMM_100_WVALID),
        .AP_AXIMM_100_WREADY(AP_AXIMM_100_WREADY),
        .AP_AXIMM_100_BRESP(AP_AXIMM_100_BRESP),
        .AP_AXIMM_100_BVALID(AP_AXIMM_100_BVALID),
        .AP_AXIMM_100_BREADY(AP_AXIMM_100_BREADY),
        .AP_AXIMM_100_ARADDR(AP_AXIMM_100_ARADDR),
        .AP_AXIMM_100_ARLEN(AP_AXIMM_100_ARLEN),
        .AP_AXIMM_100_ARSIZE(AP_AXIMM_100_ARSIZE),
        .AP_AXIMM_100_ARBURST(AP_AXIMM_100_ARBURST),
        .AP_AXIMM_100_ARLOCK(AP_AXIMM_100_ARLOCK),
        .AP_AXIMM_100_ARCACHE(AP_AXIMM_100_ARCACHE),
        .AP_AXIMM_100_ARPROT(AP_AXIMM_100_ARPROT),
        .AP_AXIMM_100_ARREGION(AP_AXIMM_100_ARREGION),
        .AP_AXIMM_100_ARQOS(AP_AXIMM_100_ARQOS),
        .AP_AXIMM_100_ARVALID(AP_AXIMM_100_ARVALID),
        .AP_AXIMM_100_ARREADY(AP_AXIMM_100_ARREADY),
        .AP_AXIMM_100_RDATA(AP_AXIMM_100_RDATA),
        .AP_AXIMM_100_RRESP(AP_AXIMM_100_RRESP),
        .AP_AXIMM_100_RLAST(AP_AXIMM_100_RLAST),
        .AP_AXIMM_100_RVALID(AP_AXIMM_100_RVALID),
        .AP_AXIMM_100_RREADY(AP_AXIMM_100_RREADY),
        .M_AXIMM_100_AWADDR(M_AXIMM_100_AWADDR),
        .M_AXIMM_100_AWLEN(M_AXIMM_100_AWLEN),
        .M_AXIMM_100_AWSIZE(M_AXIMM_100_AWSIZE),
        .M_AXIMM_100_AWBURST(M_AXIMM_100_AWBURST),
        .M_AXIMM_100_AWLOCK(M_AXIMM_100_AWLOCK),
        .M_AXIMM_100_AWCACHE(M_AXIMM_100_AWCACHE),
        .M_AXIMM_100_AWPROT(M_AXIMM_100_AWPROT),
        .M_AXIMM_100_AWREGION(M_AXIMM_100_AWREGION),
        .M_AXIMM_100_AWQOS(M_AXIMM_100_AWQOS),
        .M_AXIMM_100_AWVALID(M_AXIMM_100_AWVALID),
        .M_AXIMM_100_AWREADY(M_AXIMM_100_AWREADY),
        .M_AXIMM_100_WDATA(M_AXIMM_100_WDATA),
        .M_AXIMM_100_WSTRB(M_AXIMM_100_WSTRB),
        .M_AXIMM_100_WLAST(M_AXIMM_100_WLAST),
        .M_AXIMM_100_WVALID(M_AXIMM_100_WVALID),
        .M_AXIMM_100_WREADY(M_AXIMM_100_WREADY),
        .M_AXIMM_100_BRESP(M_AXIMM_100_BRESP),
        .M_AXIMM_100_BVALID(M_AXIMM_100_BVALID),
        .M_AXIMM_100_BREADY(M_AXIMM_100_BREADY),
        .M_AXIMM_100_ARADDR(M_AXIMM_100_ARADDR),
        .M_AXIMM_100_ARLEN(M_AXIMM_100_ARLEN),
        .M_AXIMM_100_ARSIZE(M_AXIMM_100_ARSIZE),
        .M_AXIMM_100_ARBURST(M_AXIMM_100_ARBURST),
        .M_AXIMM_100_ARLOCK(M_AXIMM_100_ARLOCK),
        .M_AXIMM_100_ARCACHE(M_AXIMM_100_ARCACHE),
        .M_AXIMM_100_ARPROT(M_AXIMM_100_ARPROT),
        .M_AXIMM_100_ARREGION(M_AXIMM_100_ARREGION),
        .M_AXIMM_100_ARQOS(M_AXIMM_100_ARQOS),
        .M_AXIMM_100_ARVALID(M_AXIMM_100_ARVALID),
        .M_AXIMM_100_ARREADY(M_AXIMM_100_ARREADY),
        .M_AXIMM_100_RDATA(M_AXIMM_100_RDATA),
        .M_AXIMM_100_RRESP(M_AXIMM_100_RRESP),
        .M_AXIMM_100_RLAST(M_AXIMM_100_RLAST),
        .M_AXIMM_100_RVALID(M_AXIMM_100_RVALID),
        .M_AXIMM_100_RREADY(M_AXIMM_100_RREADY),
        .AP_AXIMM_101_AWADDR(AP_AXIMM_101_AWADDR),
        .AP_AXIMM_101_AWLEN(AP_AXIMM_101_AWLEN),
        .AP_AXIMM_101_AWSIZE(AP_AXIMM_101_AWSIZE),
        .AP_AXIMM_101_AWBURST(AP_AXIMM_101_AWBURST),
        .AP_AXIMM_101_AWLOCK(AP_AXIMM_101_AWLOCK),
        .AP_AXIMM_101_AWCACHE(AP_AXIMM_101_AWCACHE),
        .AP_AXIMM_101_AWPROT(AP_AXIMM_101_AWPROT),
        .AP_AXIMM_101_AWREGION(AP_AXIMM_101_AWREGION),
        .AP_AXIMM_101_AWQOS(AP_AXIMM_101_AWQOS),
        .AP_AXIMM_101_AWVALID(AP_AXIMM_101_AWVALID),
        .AP_AXIMM_101_AWREADY(AP_AXIMM_101_AWREADY),
        .AP_AXIMM_101_WDATA(AP_AXIMM_101_WDATA),
        .AP_AXIMM_101_WSTRB(AP_AXIMM_101_WSTRB),
        .AP_AXIMM_101_WLAST(AP_AXIMM_101_WLAST),
        .AP_AXIMM_101_WVALID(AP_AXIMM_101_WVALID),
        .AP_AXIMM_101_WREADY(AP_AXIMM_101_WREADY),
        .AP_AXIMM_101_BRESP(AP_AXIMM_101_BRESP),
        .AP_AXIMM_101_BVALID(AP_AXIMM_101_BVALID),
        .AP_AXIMM_101_BREADY(AP_AXIMM_101_BREADY),
        .AP_AXIMM_101_ARADDR(AP_AXIMM_101_ARADDR),
        .AP_AXIMM_101_ARLEN(AP_AXIMM_101_ARLEN),
        .AP_AXIMM_101_ARSIZE(AP_AXIMM_101_ARSIZE),
        .AP_AXIMM_101_ARBURST(AP_AXIMM_101_ARBURST),
        .AP_AXIMM_101_ARLOCK(AP_AXIMM_101_ARLOCK),
        .AP_AXIMM_101_ARCACHE(AP_AXIMM_101_ARCACHE),
        .AP_AXIMM_101_ARPROT(AP_AXIMM_101_ARPROT),
        .AP_AXIMM_101_ARREGION(AP_AXIMM_101_ARREGION),
        .AP_AXIMM_101_ARQOS(AP_AXIMM_101_ARQOS),
        .AP_AXIMM_101_ARVALID(AP_AXIMM_101_ARVALID),
        .AP_AXIMM_101_ARREADY(AP_AXIMM_101_ARREADY),
        .AP_AXIMM_101_RDATA(AP_AXIMM_101_RDATA),
        .AP_AXIMM_101_RRESP(AP_AXIMM_101_RRESP),
        .AP_AXIMM_101_RLAST(AP_AXIMM_101_RLAST),
        .AP_AXIMM_101_RVALID(AP_AXIMM_101_RVALID),
        .AP_AXIMM_101_RREADY(AP_AXIMM_101_RREADY),
        .M_AXIMM_101_AWADDR(M_AXIMM_101_AWADDR),
        .M_AXIMM_101_AWLEN(M_AXIMM_101_AWLEN),
        .M_AXIMM_101_AWSIZE(M_AXIMM_101_AWSIZE),
        .M_AXIMM_101_AWBURST(M_AXIMM_101_AWBURST),
        .M_AXIMM_101_AWLOCK(M_AXIMM_101_AWLOCK),
        .M_AXIMM_101_AWCACHE(M_AXIMM_101_AWCACHE),
        .M_AXIMM_101_AWPROT(M_AXIMM_101_AWPROT),
        .M_AXIMM_101_AWREGION(M_AXIMM_101_AWREGION),
        .M_AXIMM_101_AWQOS(M_AXIMM_101_AWQOS),
        .M_AXIMM_101_AWVALID(M_AXIMM_101_AWVALID),
        .M_AXIMM_101_AWREADY(M_AXIMM_101_AWREADY),
        .M_AXIMM_101_WDATA(M_AXIMM_101_WDATA),
        .M_AXIMM_101_WSTRB(M_AXIMM_101_WSTRB),
        .M_AXIMM_101_WLAST(M_AXIMM_101_WLAST),
        .M_AXIMM_101_WVALID(M_AXIMM_101_WVALID),
        .M_AXIMM_101_WREADY(M_AXIMM_101_WREADY),
        .M_AXIMM_101_BRESP(M_AXIMM_101_BRESP),
        .M_AXIMM_101_BVALID(M_AXIMM_101_BVALID),
        .M_AXIMM_101_BREADY(M_AXIMM_101_BREADY),
        .M_AXIMM_101_ARADDR(M_AXIMM_101_ARADDR),
        .M_AXIMM_101_ARLEN(M_AXIMM_101_ARLEN),
        .M_AXIMM_101_ARSIZE(M_AXIMM_101_ARSIZE),
        .M_AXIMM_101_ARBURST(M_AXIMM_101_ARBURST),
        .M_AXIMM_101_ARLOCK(M_AXIMM_101_ARLOCK),
        .M_AXIMM_101_ARCACHE(M_AXIMM_101_ARCACHE),
        .M_AXIMM_101_ARPROT(M_AXIMM_101_ARPROT),
        .M_AXIMM_101_ARREGION(M_AXIMM_101_ARREGION),
        .M_AXIMM_101_ARQOS(M_AXIMM_101_ARQOS),
        .M_AXIMM_101_ARVALID(M_AXIMM_101_ARVALID),
        .M_AXIMM_101_ARREADY(M_AXIMM_101_ARREADY),
        .M_AXIMM_101_RDATA(M_AXIMM_101_RDATA),
        .M_AXIMM_101_RRESP(M_AXIMM_101_RRESP),
        .M_AXIMM_101_RLAST(M_AXIMM_101_RLAST),
        .M_AXIMM_101_RVALID(M_AXIMM_101_RVALID),
        .M_AXIMM_101_RREADY(M_AXIMM_101_RREADY),
        .AP_AXIMM_102_AWADDR(AP_AXIMM_102_AWADDR),
        .AP_AXIMM_102_AWLEN(AP_AXIMM_102_AWLEN),
        .AP_AXIMM_102_AWSIZE(AP_AXIMM_102_AWSIZE),
        .AP_AXIMM_102_AWBURST(AP_AXIMM_102_AWBURST),
        .AP_AXIMM_102_AWLOCK(AP_AXIMM_102_AWLOCK),
        .AP_AXIMM_102_AWCACHE(AP_AXIMM_102_AWCACHE),
        .AP_AXIMM_102_AWPROT(AP_AXIMM_102_AWPROT),
        .AP_AXIMM_102_AWREGION(AP_AXIMM_102_AWREGION),
        .AP_AXIMM_102_AWQOS(AP_AXIMM_102_AWQOS),
        .AP_AXIMM_102_AWVALID(AP_AXIMM_102_AWVALID),
        .AP_AXIMM_102_AWREADY(AP_AXIMM_102_AWREADY),
        .AP_AXIMM_102_WDATA(AP_AXIMM_102_WDATA),
        .AP_AXIMM_102_WSTRB(AP_AXIMM_102_WSTRB),
        .AP_AXIMM_102_WLAST(AP_AXIMM_102_WLAST),
        .AP_AXIMM_102_WVALID(AP_AXIMM_102_WVALID),
        .AP_AXIMM_102_WREADY(AP_AXIMM_102_WREADY),
        .AP_AXIMM_102_BRESP(AP_AXIMM_102_BRESP),
        .AP_AXIMM_102_BVALID(AP_AXIMM_102_BVALID),
        .AP_AXIMM_102_BREADY(AP_AXIMM_102_BREADY),
        .AP_AXIMM_102_ARADDR(AP_AXIMM_102_ARADDR),
        .AP_AXIMM_102_ARLEN(AP_AXIMM_102_ARLEN),
        .AP_AXIMM_102_ARSIZE(AP_AXIMM_102_ARSIZE),
        .AP_AXIMM_102_ARBURST(AP_AXIMM_102_ARBURST),
        .AP_AXIMM_102_ARLOCK(AP_AXIMM_102_ARLOCK),
        .AP_AXIMM_102_ARCACHE(AP_AXIMM_102_ARCACHE),
        .AP_AXIMM_102_ARPROT(AP_AXIMM_102_ARPROT),
        .AP_AXIMM_102_ARREGION(AP_AXIMM_102_ARREGION),
        .AP_AXIMM_102_ARQOS(AP_AXIMM_102_ARQOS),
        .AP_AXIMM_102_ARVALID(AP_AXIMM_102_ARVALID),
        .AP_AXIMM_102_ARREADY(AP_AXIMM_102_ARREADY),
        .AP_AXIMM_102_RDATA(AP_AXIMM_102_RDATA),
        .AP_AXIMM_102_RRESP(AP_AXIMM_102_RRESP),
        .AP_AXIMM_102_RLAST(AP_AXIMM_102_RLAST),
        .AP_AXIMM_102_RVALID(AP_AXIMM_102_RVALID),
        .AP_AXIMM_102_RREADY(AP_AXIMM_102_RREADY),
        .M_AXIMM_102_AWADDR(M_AXIMM_102_AWADDR),
        .M_AXIMM_102_AWLEN(M_AXIMM_102_AWLEN),
        .M_AXIMM_102_AWSIZE(M_AXIMM_102_AWSIZE),
        .M_AXIMM_102_AWBURST(M_AXIMM_102_AWBURST),
        .M_AXIMM_102_AWLOCK(M_AXIMM_102_AWLOCK),
        .M_AXIMM_102_AWCACHE(M_AXIMM_102_AWCACHE),
        .M_AXIMM_102_AWPROT(M_AXIMM_102_AWPROT),
        .M_AXIMM_102_AWREGION(M_AXIMM_102_AWREGION),
        .M_AXIMM_102_AWQOS(M_AXIMM_102_AWQOS),
        .M_AXIMM_102_AWVALID(M_AXIMM_102_AWVALID),
        .M_AXIMM_102_AWREADY(M_AXIMM_102_AWREADY),
        .M_AXIMM_102_WDATA(M_AXIMM_102_WDATA),
        .M_AXIMM_102_WSTRB(M_AXIMM_102_WSTRB),
        .M_AXIMM_102_WLAST(M_AXIMM_102_WLAST),
        .M_AXIMM_102_WVALID(M_AXIMM_102_WVALID),
        .M_AXIMM_102_WREADY(M_AXIMM_102_WREADY),
        .M_AXIMM_102_BRESP(M_AXIMM_102_BRESP),
        .M_AXIMM_102_BVALID(M_AXIMM_102_BVALID),
        .M_AXIMM_102_BREADY(M_AXIMM_102_BREADY),
        .M_AXIMM_102_ARADDR(M_AXIMM_102_ARADDR),
        .M_AXIMM_102_ARLEN(M_AXIMM_102_ARLEN),
        .M_AXIMM_102_ARSIZE(M_AXIMM_102_ARSIZE),
        .M_AXIMM_102_ARBURST(M_AXIMM_102_ARBURST),
        .M_AXIMM_102_ARLOCK(M_AXIMM_102_ARLOCK),
        .M_AXIMM_102_ARCACHE(M_AXIMM_102_ARCACHE),
        .M_AXIMM_102_ARPROT(M_AXIMM_102_ARPROT),
        .M_AXIMM_102_ARREGION(M_AXIMM_102_ARREGION),
        .M_AXIMM_102_ARQOS(M_AXIMM_102_ARQOS),
        .M_AXIMM_102_ARVALID(M_AXIMM_102_ARVALID),
        .M_AXIMM_102_ARREADY(M_AXIMM_102_ARREADY),
        .M_AXIMM_102_RDATA(M_AXIMM_102_RDATA),
        .M_AXIMM_102_RRESP(M_AXIMM_102_RRESP),
        .M_AXIMM_102_RLAST(M_AXIMM_102_RLAST),
        .M_AXIMM_102_RVALID(M_AXIMM_102_RVALID),
        .M_AXIMM_102_RREADY(M_AXIMM_102_RREADY),
        .AP_AXIMM_103_AWADDR(AP_AXIMM_103_AWADDR),
        .AP_AXIMM_103_AWLEN(AP_AXIMM_103_AWLEN),
        .AP_AXIMM_103_AWSIZE(AP_AXIMM_103_AWSIZE),
        .AP_AXIMM_103_AWBURST(AP_AXIMM_103_AWBURST),
        .AP_AXIMM_103_AWLOCK(AP_AXIMM_103_AWLOCK),
        .AP_AXIMM_103_AWCACHE(AP_AXIMM_103_AWCACHE),
        .AP_AXIMM_103_AWPROT(AP_AXIMM_103_AWPROT),
        .AP_AXIMM_103_AWREGION(AP_AXIMM_103_AWREGION),
        .AP_AXIMM_103_AWQOS(AP_AXIMM_103_AWQOS),
        .AP_AXIMM_103_AWVALID(AP_AXIMM_103_AWVALID),
        .AP_AXIMM_103_AWREADY(AP_AXIMM_103_AWREADY),
        .AP_AXIMM_103_WDATA(AP_AXIMM_103_WDATA),
        .AP_AXIMM_103_WSTRB(AP_AXIMM_103_WSTRB),
        .AP_AXIMM_103_WLAST(AP_AXIMM_103_WLAST),
        .AP_AXIMM_103_WVALID(AP_AXIMM_103_WVALID),
        .AP_AXIMM_103_WREADY(AP_AXIMM_103_WREADY),
        .AP_AXIMM_103_BRESP(AP_AXIMM_103_BRESP),
        .AP_AXIMM_103_BVALID(AP_AXIMM_103_BVALID),
        .AP_AXIMM_103_BREADY(AP_AXIMM_103_BREADY),
        .AP_AXIMM_103_ARADDR(AP_AXIMM_103_ARADDR),
        .AP_AXIMM_103_ARLEN(AP_AXIMM_103_ARLEN),
        .AP_AXIMM_103_ARSIZE(AP_AXIMM_103_ARSIZE),
        .AP_AXIMM_103_ARBURST(AP_AXIMM_103_ARBURST),
        .AP_AXIMM_103_ARLOCK(AP_AXIMM_103_ARLOCK),
        .AP_AXIMM_103_ARCACHE(AP_AXIMM_103_ARCACHE),
        .AP_AXIMM_103_ARPROT(AP_AXIMM_103_ARPROT),
        .AP_AXIMM_103_ARREGION(AP_AXIMM_103_ARREGION),
        .AP_AXIMM_103_ARQOS(AP_AXIMM_103_ARQOS),
        .AP_AXIMM_103_ARVALID(AP_AXIMM_103_ARVALID),
        .AP_AXIMM_103_ARREADY(AP_AXIMM_103_ARREADY),
        .AP_AXIMM_103_RDATA(AP_AXIMM_103_RDATA),
        .AP_AXIMM_103_RRESP(AP_AXIMM_103_RRESP),
        .AP_AXIMM_103_RLAST(AP_AXIMM_103_RLAST),
        .AP_AXIMM_103_RVALID(AP_AXIMM_103_RVALID),
        .AP_AXIMM_103_RREADY(AP_AXIMM_103_RREADY),
        .M_AXIMM_103_AWADDR(M_AXIMM_103_AWADDR),
        .M_AXIMM_103_AWLEN(M_AXIMM_103_AWLEN),
        .M_AXIMM_103_AWSIZE(M_AXIMM_103_AWSIZE),
        .M_AXIMM_103_AWBURST(M_AXIMM_103_AWBURST),
        .M_AXIMM_103_AWLOCK(M_AXIMM_103_AWLOCK),
        .M_AXIMM_103_AWCACHE(M_AXIMM_103_AWCACHE),
        .M_AXIMM_103_AWPROT(M_AXIMM_103_AWPROT),
        .M_AXIMM_103_AWREGION(M_AXIMM_103_AWREGION),
        .M_AXIMM_103_AWQOS(M_AXIMM_103_AWQOS),
        .M_AXIMM_103_AWVALID(M_AXIMM_103_AWVALID),
        .M_AXIMM_103_AWREADY(M_AXIMM_103_AWREADY),
        .M_AXIMM_103_WDATA(M_AXIMM_103_WDATA),
        .M_AXIMM_103_WSTRB(M_AXIMM_103_WSTRB),
        .M_AXIMM_103_WLAST(M_AXIMM_103_WLAST),
        .M_AXIMM_103_WVALID(M_AXIMM_103_WVALID),
        .M_AXIMM_103_WREADY(M_AXIMM_103_WREADY),
        .M_AXIMM_103_BRESP(M_AXIMM_103_BRESP),
        .M_AXIMM_103_BVALID(M_AXIMM_103_BVALID),
        .M_AXIMM_103_BREADY(M_AXIMM_103_BREADY),
        .M_AXIMM_103_ARADDR(M_AXIMM_103_ARADDR),
        .M_AXIMM_103_ARLEN(M_AXIMM_103_ARLEN),
        .M_AXIMM_103_ARSIZE(M_AXIMM_103_ARSIZE),
        .M_AXIMM_103_ARBURST(M_AXIMM_103_ARBURST),
        .M_AXIMM_103_ARLOCK(M_AXIMM_103_ARLOCK),
        .M_AXIMM_103_ARCACHE(M_AXIMM_103_ARCACHE),
        .M_AXIMM_103_ARPROT(M_AXIMM_103_ARPROT),
        .M_AXIMM_103_ARREGION(M_AXIMM_103_ARREGION),
        .M_AXIMM_103_ARQOS(M_AXIMM_103_ARQOS),
        .M_AXIMM_103_ARVALID(M_AXIMM_103_ARVALID),
        .M_AXIMM_103_ARREADY(M_AXIMM_103_ARREADY),
        .M_AXIMM_103_RDATA(M_AXIMM_103_RDATA),
        .M_AXIMM_103_RRESP(M_AXIMM_103_RRESP),
        .M_AXIMM_103_RLAST(M_AXIMM_103_RLAST),
        .M_AXIMM_103_RVALID(M_AXIMM_103_RVALID),
        .M_AXIMM_103_RREADY(M_AXIMM_103_RREADY),
        .AP_AXIMM_104_AWADDR(AP_AXIMM_104_AWADDR),
        .AP_AXIMM_104_AWLEN(AP_AXIMM_104_AWLEN),
        .AP_AXIMM_104_AWSIZE(AP_AXIMM_104_AWSIZE),
        .AP_AXIMM_104_AWBURST(AP_AXIMM_104_AWBURST),
        .AP_AXIMM_104_AWLOCK(AP_AXIMM_104_AWLOCK),
        .AP_AXIMM_104_AWCACHE(AP_AXIMM_104_AWCACHE),
        .AP_AXIMM_104_AWPROT(AP_AXIMM_104_AWPROT),
        .AP_AXIMM_104_AWREGION(AP_AXIMM_104_AWREGION),
        .AP_AXIMM_104_AWQOS(AP_AXIMM_104_AWQOS),
        .AP_AXIMM_104_AWVALID(AP_AXIMM_104_AWVALID),
        .AP_AXIMM_104_AWREADY(AP_AXIMM_104_AWREADY),
        .AP_AXIMM_104_WDATA(AP_AXIMM_104_WDATA),
        .AP_AXIMM_104_WSTRB(AP_AXIMM_104_WSTRB),
        .AP_AXIMM_104_WLAST(AP_AXIMM_104_WLAST),
        .AP_AXIMM_104_WVALID(AP_AXIMM_104_WVALID),
        .AP_AXIMM_104_WREADY(AP_AXIMM_104_WREADY),
        .AP_AXIMM_104_BRESP(AP_AXIMM_104_BRESP),
        .AP_AXIMM_104_BVALID(AP_AXIMM_104_BVALID),
        .AP_AXIMM_104_BREADY(AP_AXIMM_104_BREADY),
        .AP_AXIMM_104_ARADDR(AP_AXIMM_104_ARADDR),
        .AP_AXIMM_104_ARLEN(AP_AXIMM_104_ARLEN),
        .AP_AXIMM_104_ARSIZE(AP_AXIMM_104_ARSIZE),
        .AP_AXIMM_104_ARBURST(AP_AXIMM_104_ARBURST),
        .AP_AXIMM_104_ARLOCK(AP_AXIMM_104_ARLOCK),
        .AP_AXIMM_104_ARCACHE(AP_AXIMM_104_ARCACHE),
        .AP_AXIMM_104_ARPROT(AP_AXIMM_104_ARPROT),
        .AP_AXIMM_104_ARREGION(AP_AXIMM_104_ARREGION),
        .AP_AXIMM_104_ARQOS(AP_AXIMM_104_ARQOS),
        .AP_AXIMM_104_ARVALID(AP_AXIMM_104_ARVALID),
        .AP_AXIMM_104_ARREADY(AP_AXIMM_104_ARREADY),
        .AP_AXIMM_104_RDATA(AP_AXIMM_104_RDATA),
        .AP_AXIMM_104_RRESP(AP_AXIMM_104_RRESP),
        .AP_AXIMM_104_RLAST(AP_AXIMM_104_RLAST),
        .AP_AXIMM_104_RVALID(AP_AXIMM_104_RVALID),
        .AP_AXIMM_104_RREADY(AP_AXIMM_104_RREADY),
        .M_AXIMM_104_AWADDR(M_AXIMM_104_AWADDR),
        .M_AXIMM_104_AWLEN(M_AXIMM_104_AWLEN),
        .M_AXIMM_104_AWSIZE(M_AXIMM_104_AWSIZE),
        .M_AXIMM_104_AWBURST(M_AXIMM_104_AWBURST),
        .M_AXIMM_104_AWLOCK(M_AXIMM_104_AWLOCK),
        .M_AXIMM_104_AWCACHE(M_AXIMM_104_AWCACHE),
        .M_AXIMM_104_AWPROT(M_AXIMM_104_AWPROT),
        .M_AXIMM_104_AWREGION(M_AXIMM_104_AWREGION),
        .M_AXIMM_104_AWQOS(M_AXIMM_104_AWQOS),
        .M_AXIMM_104_AWVALID(M_AXIMM_104_AWVALID),
        .M_AXIMM_104_AWREADY(M_AXIMM_104_AWREADY),
        .M_AXIMM_104_WDATA(M_AXIMM_104_WDATA),
        .M_AXIMM_104_WSTRB(M_AXIMM_104_WSTRB),
        .M_AXIMM_104_WLAST(M_AXIMM_104_WLAST),
        .M_AXIMM_104_WVALID(M_AXIMM_104_WVALID),
        .M_AXIMM_104_WREADY(M_AXIMM_104_WREADY),
        .M_AXIMM_104_BRESP(M_AXIMM_104_BRESP),
        .M_AXIMM_104_BVALID(M_AXIMM_104_BVALID),
        .M_AXIMM_104_BREADY(M_AXIMM_104_BREADY),
        .M_AXIMM_104_ARADDR(M_AXIMM_104_ARADDR),
        .M_AXIMM_104_ARLEN(M_AXIMM_104_ARLEN),
        .M_AXIMM_104_ARSIZE(M_AXIMM_104_ARSIZE),
        .M_AXIMM_104_ARBURST(M_AXIMM_104_ARBURST),
        .M_AXIMM_104_ARLOCK(M_AXIMM_104_ARLOCK),
        .M_AXIMM_104_ARCACHE(M_AXIMM_104_ARCACHE),
        .M_AXIMM_104_ARPROT(M_AXIMM_104_ARPROT),
        .M_AXIMM_104_ARREGION(M_AXIMM_104_ARREGION),
        .M_AXIMM_104_ARQOS(M_AXIMM_104_ARQOS),
        .M_AXIMM_104_ARVALID(M_AXIMM_104_ARVALID),
        .M_AXIMM_104_ARREADY(M_AXIMM_104_ARREADY),
        .M_AXIMM_104_RDATA(M_AXIMM_104_RDATA),
        .M_AXIMM_104_RRESP(M_AXIMM_104_RRESP),
        .M_AXIMM_104_RLAST(M_AXIMM_104_RLAST),
        .M_AXIMM_104_RVALID(M_AXIMM_104_RVALID),
        .M_AXIMM_104_RREADY(M_AXIMM_104_RREADY),
        .AP_AXIMM_105_AWADDR(AP_AXIMM_105_AWADDR),
        .AP_AXIMM_105_AWLEN(AP_AXIMM_105_AWLEN),
        .AP_AXIMM_105_AWSIZE(AP_AXIMM_105_AWSIZE),
        .AP_AXIMM_105_AWBURST(AP_AXIMM_105_AWBURST),
        .AP_AXIMM_105_AWLOCK(AP_AXIMM_105_AWLOCK),
        .AP_AXIMM_105_AWCACHE(AP_AXIMM_105_AWCACHE),
        .AP_AXIMM_105_AWPROT(AP_AXIMM_105_AWPROT),
        .AP_AXIMM_105_AWREGION(AP_AXIMM_105_AWREGION),
        .AP_AXIMM_105_AWQOS(AP_AXIMM_105_AWQOS),
        .AP_AXIMM_105_AWVALID(AP_AXIMM_105_AWVALID),
        .AP_AXIMM_105_AWREADY(AP_AXIMM_105_AWREADY),
        .AP_AXIMM_105_WDATA(AP_AXIMM_105_WDATA),
        .AP_AXIMM_105_WSTRB(AP_AXIMM_105_WSTRB),
        .AP_AXIMM_105_WLAST(AP_AXIMM_105_WLAST),
        .AP_AXIMM_105_WVALID(AP_AXIMM_105_WVALID),
        .AP_AXIMM_105_WREADY(AP_AXIMM_105_WREADY),
        .AP_AXIMM_105_BRESP(AP_AXIMM_105_BRESP),
        .AP_AXIMM_105_BVALID(AP_AXIMM_105_BVALID),
        .AP_AXIMM_105_BREADY(AP_AXIMM_105_BREADY),
        .AP_AXIMM_105_ARADDR(AP_AXIMM_105_ARADDR),
        .AP_AXIMM_105_ARLEN(AP_AXIMM_105_ARLEN),
        .AP_AXIMM_105_ARSIZE(AP_AXIMM_105_ARSIZE),
        .AP_AXIMM_105_ARBURST(AP_AXIMM_105_ARBURST),
        .AP_AXIMM_105_ARLOCK(AP_AXIMM_105_ARLOCK),
        .AP_AXIMM_105_ARCACHE(AP_AXIMM_105_ARCACHE),
        .AP_AXIMM_105_ARPROT(AP_AXIMM_105_ARPROT),
        .AP_AXIMM_105_ARREGION(AP_AXIMM_105_ARREGION),
        .AP_AXIMM_105_ARQOS(AP_AXIMM_105_ARQOS),
        .AP_AXIMM_105_ARVALID(AP_AXIMM_105_ARVALID),
        .AP_AXIMM_105_ARREADY(AP_AXIMM_105_ARREADY),
        .AP_AXIMM_105_RDATA(AP_AXIMM_105_RDATA),
        .AP_AXIMM_105_RRESP(AP_AXIMM_105_RRESP),
        .AP_AXIMM_105_RLAST(AP_AXIMM_105_RLAST),
        .AP_AXIMM_105_RVALID(AP_AXIMM_105_RVALID),
        .AP_AXIMM_105_RREADY(AP_AXIMM_105_RREADY),
        .M_AXIMM_105_AWADDR(M_AXIMM_105_AWADDR),
        .M_AXIMM_105_AWLEN(M_AXIMM_105_AWLEN),
        .M_AXIMM_105_AWSIZE(M_AXIMM_105_AWSIZE),
        .M_AXIMM_105_AWBURST(M_AXIMM_105_AWBURST),
        .M_AXIMM_105_AWLOCK(M_AXIMM_105_AWLOCK),
        .M_AXIMM_105_AWCACHE(M_AXIMM_105_AWCACHE),
        .M_AXIMM_105_AWPROT(M_AXIMM_105_AWPROT),
        .M_AXIMM_105_AWREGION(M_AXIMM_105_AWREGION),
        .M_AXIMM_105_AWQOS(M_AXIMM_105_AWQOS),
        .M_AXIMM_105_AWVALID(M_AXIMM_105_AWVALID),
        .M_AXIMM_105_AWREADY(M_AXIMM_105_AWREADY),
        .M_AXIMM_105_WDATA(M_AXIMM_105_WDATA),
        .M_AXIMM_105_WSTRB(M_AXIMM_105_WSTRB),
        .M_AXIMM_105_WLAST(M_AXIMM_105_WLAST),
        .M_AXIMM_105_WVALID(M_AXIMM_105_WVALID),
        .M_AXIMM_105_WREADY(M_AXIMM_105_WREADY),
        .M_AXIMM_105_BRESP(M_AXIMM_105_BRESP),
        .M_AXIMM_105_BVALID(M_AXIMM_105_BVALID),
        .M_AXIMM_105_BREADY(M_AXIMM_105_BREADY),
        .M_AXIMM_105_ARADDR(M_AXIMM_105_ARADDR),
        .M_AXIMM_105_ARLEN(M_AXIMM_105_ARLEN),
        .M_AXIMM_105_ARSIZE(M_AXIMM_105_ARSIZE),
        .M_AXIMM_105_ARBURST(M_AXIMM_105_ARBURST),
        .M_AXIMM_105_ARLOCK(M_AXIMM_105_ARLOCK),
        .M_AXIMM_105_ARCACHE(M_AXIMM_105_ARCACHE),
        .M_AXIMM_105_ARPROT(M_AXIMM_105_ARPROT),
        .M_AXIMM_105_ARREGION(M_AXIMM_105_ARREGION),
        .M_AXIMM_105_ARQOS(M_AXIMM_105_ARQOS),
        .M_AXIMM_105_ARVALID(M_AXIMM_105_ARVALID),
        .M_AXIMM_105_ARREADY(M_AXIMM_105_ARREADY),
        .M_AXIMM_105_RDATA(M_AXIMM_105_RDATA),
        .M_AXIMM_105_RRESP(M_AXIMM_105_RRESP),
        .M_AXIMM_105_RLAST(M_AXIMM_105_RLAST),
        .M_AXIMM_105_RVALID(M_AXIMM_105_RVALID),
        .M_AXIMM_105_RREADY(M_AXIMM_105_RREADY),
        .AP_AXIMM_106_AWADDR(AP_AXIMM_106_AWADDR),
        .AP_AXIMM_106_AWLEN(AP_AXIMM_106_AWLEN),
        .AP_AXIMM_106_AWSIZE(AP_AXIMM_106_AWSIZE),
        .AP_AXIMM_106_AWBURST(AP_AXIMM_106_AWBURST),
        .AP_AXIMM_106_AWLOCK(AP_AXIMM_106_AWLOCK),
        .AP_AXIMM_106_AWCACHE(AP_AXIMM_106_AWCACHE),
        .AP_AXIMM_106_AWPROT(AP_AXIMM_106_AWPROT),
        .AP_AXIMM_106_AWREGION(AP_AXIMM_106_AWREGION),
        .AP_AXIMM_106_AWQOS(AP_AXIMM_106_AWQOS),
        .AP_AXIMM_106_AWVALID(AP_AXIMM_106_AWVALID),
        .AP_AXIMM_106_AWREADY(AP_AXIMM_106_AWREADY),
        .AP_AXIMM_106_WDATA(AP_AXIMM_106_WDATA),
        .AP_AXIMM_106_WSTRB(AP_AXIMM_106_WSTRB),
        .AP_AXIMM_106_WLAST(AP_AXIMM_106_WLAST),
        .AP_AXIMM_106_WVALID(AP_AXIMM_106_WVALID),
        .AP_AXIMM_106_WREADY(AP_AXIMM_106_WREADY),
        .AP_AXIMM_106_BRESP(AP_AXIMM_106_BRESP),
        .AP_AXIMM_106_BVALID(AP_AXIMM_106_BVALID),
        .AP_AXIMM_106_BREADY(AP_AXIMM_106_BREADY),
        .AP_AXIMM_106_ARADDR(AP_AXIMM_106_ARADDR),
        .AP_AXIMM_106_ARLEN(AP_AXIMM_106_ARLEN),
        .AP_AXIMM_106_ARSIZE(AP_AXIMM_106_ARSIZE),
        .AP_AXIMM_106_ARBURST(AP_AXIMM_106_ARBURST),
        .AP_AXIMM_106_ARLOCK(AP_AXIMM_106_ARLOCK),
        .AP_AXIMM_106_ARCACHE(AP_AXIMM_106_ARCACHE),
        .AP_AXIMM_106_ARPROT(AP_AXIMM_106_ARPROT),
        .AP_AXIMM_106_ARREGION(AP_AXIMM_106_ARREGION),
        .AP_AXIMM_106_ARQOS(AP_AXIMM_106_ARQOS),
        .AP_AXIMM_106_ARVALID(AP_AXIMM_106_ARVALID),
        .AP_AXIMM_106_ARREADY(AP_AXIMM_106_ARREADY),
        .AP_AXIMM_106_RDATA(AP_AXIMM_106_RDATA),
        .AP_AXIMM_106_RRESP(AP_AXIMM_106_RRESP),
        .AP_AXIMM_106_RLAST(AP_AXIMM_106_RLAST),
        .AP_AXIMM_106_RVALID(AP_AXIMM_106_RVALID),
        .AP_AXIMM_106_RREADY(AP_AXIMM_106_RREADY),
        .M_AXIMM_106_AWADDR(M_AXIMM_106_AWADDR),
        .M_AXIMM_106_AWLEN(M_AXIMM_106_AWLEN),
        .M_AXIMM_106_AWSIZE(M_AXIMM_106_AWSIZE),
        .M_AXIMM_106_AWBURST(M_AXIMM_106_AWBURST),
        .M_AXIMM_106_AWLOCK(M_AXIMM_106_AWLOCK),
        .M_AXIMM_106_AWCACHE(M_AXIMM_106_AWCACHE),
        .M_AXIMM_106_AWPROT(M_AXIMM_106_AWPROT),
        .M_AXIMM_106_AWREGION(M_AXIMM_106_AWREGION),
        .M_AXIMM_106_AWQOS(M_AXIMM_106_AWQOS),
        .M_AXIMM_106_AWVALID(M_AXIMM_106_AWVALID),
        .M_AXIMM_106_AWREADY(M_AXIMM_106_AWREADY),
        .M_AXIMM_106_WDATA(M_AXIMM_106_WDATA),
        .M_AXIMM_106_WSTRB(M_AXIMM_106_WSTRB),
        .M_AXIMM_106_WLAST(M_AXIMM_106_WLAST),
        .M_AXIMM_106_WVALID(M_AXIMM_106_WVALID),
        .M_AXIMM_106_WREADY(M_AXIMM_106_WREADY),
        .M_AXIMM_106_BRESP(M_AXIMM_106_BRESP),
        .M_AXIMM_106_BVALID(M_AXIMM_106_BVALID),
        .M_AXIMM_106_BREADY(M_AXIMM_106_BREADY),
        .M_AXIMM_106_ARADDR(M_AXIMM_106_ARADDR),
        .M_AXIMM_106_ARLEN(M_AXIMM_106_ARLEN),
        .M_AXIMM_106_ARSIZE(M_AXIMM_106_ARSIZE),
        .M_AXIMM_106_ARBURST(M_AXIMM_106_ARBURST),
        .M_AXIMM_106_ARLOCK(M_AXIMM_106_ARLOCK),
        .M_AXIMM_106_ARCACHE(M_AXIMM_106_ARCACHE),
        .M_AXIMM_106_ARPROT(M_AXIMM_106_ARPROT),
        .M_AXIMM_106_ARREGION(M_AXIMM_106_ARREGION),
        .M_AXIMM_106_ARQOS(M_AXIMM_106_ARQOS),
        .M_AXIMM_106_ARVALID(M_AXIMM_106_ARVALID),
        .M_AXIMM_106_ARREADY(M_AXIMM_106_ARREADY),
        .M_AXIMM_106_RDATA(M_AXIMM_106_RDATA),
        .M_AXIMM_106_RRESP(M_AXIMM_106_RRESP),
        .M_AXIMM_106_RLAST(M_AXIMM_106_RLAST),
        .M_AXIMM_106_RVALID(M_AXIMM_106_RVALID),
        .M_AXIMM_106_RREADY(M_AXIMM_106_RREADY),
        .AP_AXIMM_107_AWADDR(AP_AXIMM_107_AWADDR),
        .AP_AXIMM_107_AWLEN(AP_AXIMM_107_AWLEN),
        .AP_AXIMM_107_AWSIZE(AP_AXIMM_107_AWSIZE),
        .AP_AXIMM_107_AWBURST(AP_AXIMM_107_AWBURST),
        .AP_AXIMM_107_AWLOCK(AP_AXIMM_107_AWLOCK),
        .AP_AXIMM_107_AWCACHE(AP_AXIMM_107_AWCACHE),
        .AP_AXIMM_107_AWPROT(AP_AXIMM_107_AWPROT),
        .AP_AXIMM_107_AWREGION(AP_AXIMM_107_AWREGION),
        .AP_AXIMM_107_AWQOS(AP_AXIMM_107_AWQOS),
        .AP_AXIMM_107_AWVALID(AP_AXIMM_107_AWVALID),
        .AP_AXIMM_107_AWREADY(AP_AXIMM_107_AWREADY),
        .AP_AXIMM_107_WDATA(AP_AXIMM_107_WDATA),
        .AP_AXIMM_107_WSTRB(AP_AXIMM_107_WSTRB),
        .AP_AXIMM_107_WLAST(AP_AXIMM_107_WLAST),
        .AP_AXIMM_107_WVALID(AP_AXIMM_107_WVALID),
        .AP_AXIMM_107_WREADY(AP_AXIMM_107_WREADY),
        .AP_AXIMM_107_BRESP(AP_AXIMM_107_BRESP),
        .AP_AXIMM_107_BVALID(AP_AXIMM_107_BVALID),
        .AP_AXIMM_107_BREADY(AP_AXIMM_107_BREADY),
        .AP_AXIMM_107_ARADDR(AP_AXIMM_107_ARADDR),
        .AP_AXIMM_107_ARLEN(AP_AXIMM_107_ARLEN),
        .AP_AXIMM_107_ARSIZE(AP_AXIMM_107_ARSIZE),
        .AP_AXIMM_107_ARBURST(AP_AXIMM_107_ARBURST),
        .AP_AXIMM_107_ARLOCK(AP_AXIMM_107_ARLOCK),
        .AP_AXIMM_107_ARCACHE(AP_AXIMM_107_ARCACHE),
        .AP_AXIMM_107_ARPROT(AP_AXIMM_107_ARPROT),
        .AP_AXIMM_107_ARREGION(AP_AXIMM_107_ARREGION),
        .AP_AXIMM_107_ARQOS(AP_AXIMM_107_ARQOS),
        .AP_AXIMM_107_ARVALID(AP_AXIMM_107_ARVALID),
        .AP_AXIMM_107_ARREADY(AP_AXIMM_107_ARREADY),
        .AP_AXIMM_107_RDATA(AP_AXIMM_107_RDATA),
        .AP_AXIMM_107_RRESP(AP_AXIMM_107_RRESP),
        .AP_AXIMM_107_RLAST(AP_AXIMM_107_RLAST),
        .AP_AXIMM_107_RVALID(AP_AXIMM_107_RVALID),
        .AP_AXIMM_107_RREADY(AP_AXIMM_107_RREADY),
        .M_AXIMM_107_AWADDR(M_AXIMM_107_AWADDR),
        .M_AXIMM_107_AWLEN(M_AXIMM_107_AWLEN),
        .M_AXIMM_107_AWSIZE(M_AXIMM_107_AWSIZE),
        .M_AXIMM_107_AWBURST(M_AXIMM_107_AWBURST),
        .M_AXIMM_107_AWLOCK(M_AXIMM_107_AWLOCK),
        .M_AXIMM_107_AWCACHE(M_AXIMM_107_AWCACHE),
        .M_AXIMM_107_AWPROT(M_AXIMM_107_AWPROT),
        .M_AXIMM_107_AWREGION(M_AXIMM_107_AWREGION),
        .M_AXIMM_107_AWQOS(M_AXIMM_107_AWQOS),
        .M_AXIMM_107_AWVALID(M_AXIMM_107_AWVALID),
        .M_AXIMM_107_AWREADY(M_AXIMM_107_AWREADY),
        .M_AXIMM_107_WDATA(M_AXIMM_107_WDATA),
        .M_AXIMM_107_WSTRB(M_AXIMM_107_WSTRB),
        .M_AXIMM_107_WLAST(M_AXIMM_107_WLAST),
        .M_AXIMM_107_WVALID(M_AXIMM_107_WVALID),
        .M_AXIMM_107_WREADY(M_AXIMM_107_WREADY),
        .M_AXIMM_107_BRESP(M_AXIMM_107_BRESP),
        .M_AXIMM_107_BVALID(M_AXIMM_107_BVALID),
        .M_AXIMM_107_BREADY(M_AXIMM_107_BREADY),
        .M_AXIMM_107_ARADDR(M_AXIMM_107_ARADDR),
        .M_AXIMM_107_ARLEN(M_AXIMM_107_ARLEN),
        .M_AXIMM_107_ARSIZE(M_AXIMM_107_ARSIZE),
        .M_AXIMM_107_ARBURST(M_AXIMM_107_ARBURST),
        .M_AXIMM_107_ARLOCK(M_AXIMM_107_ARLOCK),
        .M_AXIMM_107_ARCACHE(M_AXIMM_107_ARCACHE),
        .M_AXIMM_107_ARPROT(M_AXIMM_107_ARPROT),
        .M_AXIMM_107_ARREGION(M_AXIMM_107_ARREGION),
        .M_AXIMM_107_ARQOS(M_AXIMM_107_ARQOS),
        .M_AXIMM_107_ARVALID(M_AXIMM_107_ARVALID),
        .M_AXIMM_107_ARREADY(M_AXIMM_107_ARREADY),
        .M_AXIMM_107_RDATA(M_AXIMM_107_RDATA),
        .M_AXIMM_107_RRESP(M_AXIMM_107_RRESP),
        .M_AXIMM_107_RLAST(M_AXIMM_107_RLAST),
        .M_AXIMM_107_RVALID(M_AXIMM_107_RVALID),
        .M_AXIMM_107_RREADY(M_AXIMM_107_RREADY),
        .AP_AXIMM_108_AWADDR(AP_AXIMM_108_AWADDR),
        .AP_AXIMM_108_AWLEN(AP_AXIMM_108_AWLEN),
        .AP_AXIMM_108_AWSIZE(AP_AXIMM_108_AWSIZE),
        .AP_AXIMM_108_AWBURST(AP_AXIMM_108_AWBURST),
        .AP_AXIMM_108_AWLOCK(AP_AXIMM_108_AWLOCK),
        .AP_AXIMM_108_AWCACHE(AP_AXIMM_108_AWCACHE),
        .AP_AXIMM_108_AWPROT(AP_AXIMM_108_AWPROT),
        .AP_AXIMM_108_AWREGION(AP_AXIMM_108_AWREGION),
        .AP_AXIMM_108_AWQOS(AP_AXIMM_108_AWQOS),
        .AP_AXIMM_108_AWVALID(AP_AXIMM_108_AWVALID),
        .AP_AXIMM_108_AWREADY(AP_AXIMM_108_AWREADY),
        .AP_AXIMM_108_WDATA(AP_AXIMM_108_WDATA),
        .AP_AXIMM_108_WSTRB(AP_AXIMM_108_WSTRB),
        .AP_AXIMM_108_WLAST(AP_AXIMM_108_WLAST),
        .AP_AXIMM_108_WVALID(AP_AXIMM_108_WVALID),
        .AP_AXIMM_108_WREADY(AP_AXIMM_108_WREADY),
        .AP_AXIMM_108_BRESP(AP_AXIMM_108_BRESP),
        .AP_AXIMM_108_BVALID(AP_AXIMM_108_BVALID),
        .AP_AXIMM_108_BREADY(AP_AXIMM_108_BREADY),
        .AP_AXIMM_108_ARADDR(AP_AXIMM_108_ARADDR),
        .AP_AXIMM_108_ARLEN(AP_AXIMM_108_ARLEN),
        .AP_AXIMM_108_ARSIZE(AP_AXIMM_108_ARSIZE),
        .AP_AXIMM_108_ARBURST(AP_AXIMM_108_ARBURST),
        .AP_AXIMM_108_ARLOCK(AP_AXIMM_108_ARLOCK),
        .AP_AXIMM_108_ARCACHE(AP_AXIMM_108_ARCACHE),
        .AP_AXIMM_108_ARPROT(AP_AXIMM_108_ARPROT),
        .AP_AXIMM_108_ARREGION(AP_AXIMM_108_ARREGION),
        .AP_AXIMM_108_ARQOS(AP_AXIMM_108_ARQOS),
        .AP_AXIMM_108_ARVALID(AP_AXIMM_108_ARVALID),
        .AP_AXIMM_108_ARREADY(AP_AXIMM_108_ARREADY),
        .AP_AXIMM_108_RDATA(AP_AXIMM_108_RDATA),
        .AP_AXIMM_108_RRESP(AP_AXIMM_108_RRESP),
        .AP_AXIMM_108_RLAST(AP_AXIMM_108_RLAST),
        .AP_AXIMM_108_RVALID(AP_AXIMM_108_RVALID),
        .AP_AXIMM_108_RREADY(AP_AXIMM_108_RREADY),
        .M_AXIMM_108_AWADDR(M_AXIMM_108_AWADDR),
        .M_AXIMM_108_AWLEN(M_AXIMM_108_AWLEN),
        .M_AXIMM_108_AWSIZE(M_AXIMM_108_AWSIZE),
        .M_AXIMM_108_AWBURST(M_AXIMM_108_AWBURST),
        .M_AXIMM_108_AWLOCK(M_AXIMM_108_AWLOCK),
        .M_AXIMM_108_AWCACHE(M_AXIMM_108_AWCACHE),
        .M_AXIMM_108_AWPROT(M_AXIMM_108_AWPROT),
        .M_AXIMM_108_AWREGION(M_AXIMM_108_AWREGION),
        .M_AXIMM_108_AWQOS(M_AXIMM_108_AWQOS),
        .M_AXIMM_108_AWVALID(M_AXIMM_108_AWVALID),
        .M_AXIMM_108_AWREADY(M_AXIMM_108_AWREADY),
        .M_AXIMM_108_WDATA(M_AXIMM_108_WDATA),
        .M_AXIMM_108_WSTRB(M_AXIMM_108_WSTRB),
        .M_AXIMM_108_WLAST(M_AXIMM_108_WLAST),
        .M_AXIMM_108_WVALID(M_AXIMM_108_WVALID),
        .M_AXIMM_108_WREADY(M_AXIMM_108_WREADY),
        .M_AXIMM_108_BRESP(M_AXIMM_108_BRESP),
        .M_AXIMM_108_BVALID(M_AXIMM_108_BVALID),
        .M_AXIMM_108_BREADY(M_AXIMM_108_BREADY),
        .M_AXIMM_108_ARADDR(M_AXIMM_108_ARADDR),
        .M_AXIMM_108_ARLEN(M_AXIMM_108_ARLEN),
        .M_AXIMM_108_ARSIZE(M_AXIMM_108_ARSIZE),
        .M_AXIMM_108_ARBURST(M_AXIMM_108_ARBURST),
        .M_AXIMM_108_ARLOCK(M_AXIMM_108_ARLOCK),
        .M_AXIMM_108_ARCACHE(M_AXIMM_108_ARCACHE),
        .M_AXIMM_108_ARPROT(M_AXIMM_108_ARPROT),
        .M_AXIMM_108_ARREGION(M_AXIMM_108_ARREGION),
        .M_AXIMM_108_ARQOS(M_AXIMM_108_ARQOS),
        .M_AXIMM_108_ARVALID(M_AXIMM_108_ARVALID),
        .M_AXIMM_108_ARREADY(M_AXIMM_108_ARREADY),
        .M_AXIMM_108_RDATA(M_AXIMM_108_RDATA),
        .M_AXIMM_108_RRESP(M_AXIMM_108_RRESP),
        .M_AXIMM_108_RLAST(M_AXIMM_108_RLAST),
        .M_AXIMM_108_RVALID(M_AXIMM_108_RVALID),
        .M_AXIMM_108_RREADY(M_AXIMM_108_RREADY),
        .AP_AXIMM_109_AWADDR(AP_AXIMM_109_AWADDR),
        .AP_AXIMM_109_AWLEN(AP_AXIMM_109_AWLEN),
        .AP_AXIMM_109_AWSIZE(AP_AXIMM_109_AWSIZE),
        .AP_AXIMM_109_AWBURST(AP_AXIMM_109_AWBURST),
        .AP_AXIMM_109_AWLOCK(AP_AXIMM_109_AWLOCK),
        .AP_AXIMM_109_AWCACHE(AP_AXIMM_109_AWCACHE),
        .AP_AXIMM_109_AWPROT(AP_AXIMM_109_AWPROT),
        .AP_AXIMM_109_AWREGION(AP_AXIMM_109_AWREGION),
        .AP_AXIMM_109_AWQOS(AP_AXIMM_109_AWQOS),
        .AP_AXIMM_109_AWVALID(AP_AXIMM_109_AWVALID),
        .AP_AXIMM_109_AWREADY(AP_AXIMM_109_AWREADY),
        .AP_AXIMM_109_WDATA(AP_AXIMM_109_WDATA),
        .AP_AXIMM_109_WSTRB(AP_AXIMM_109_WSTRB),
        .AP_AXIMM_109_WLAST(AP_AXIMM_109_WLAST),
        .AP_AXIMM_109_WVALID(AP_AXIMM_109_WVALID),
        .AP_AXIMM_109_WREADY(AP_AXIMM_109_WREADY),
        .AP_AXIMM_109_BRESP(AP_AXIMM_109_BRESP),
        .AP_AXIMM_109_BVALID(AP_AXIMM_109_BVALID),
        .AP_AXIMM_109_BREADY(AP_AXIMM_109_BREADY),
        .AP_AXIMM_109_ARADDR(AP_AXIMM_109_ARADDR),
        .AP_AXIMM_109_ARLEN(AP_AXIMM_109_ARLEN),
        .AP_AXIMM_109_ARSIZE(AP_AXIMM_109_ARSIZE),
        .AP_AXIMM_109_ARBURST(AP_AXIMM_109_ARBURST),
        .AP_AXIMM_109_ARLOCK(AP_AXIMM_109_ARLOCK),
        .AP_AXIMM_109_ARCACHE(AP_AXIMM_109_ARCACHE),
        .AP_AXIMM_109_ARPROT(AP_AXIMM_109_ARPROT),
        .AP_AXIMM_109_ARREGION(AP_AXIMM_109_ARREGION),
        .AP_AXIMM_109_ARQOS(AP_AXIMM_109_ARQOS),
        .AP_AXIMM_109_ARVALID(AP_AXIMM_109_ARVALID),
        .AP_AXIMM_109_ARREADY(AP_AXIMM_109_ARREADY),
        .AP_AXIMM_109_RDATA(AP_AXIMM_109_RDATA),
        .AP_AXIMM_109_RRESP(AP_AXIMM_109_RRESP),
        .AP_AXIMM_109_RLAST(AP_AXIMM_109_RLAST),
        .AP_AXIMM_109_RVALID(AP_AXIMM_109_RVALID),
        .AP_AXIMM_109_RREADY(AP_AXIMM_109_RREADY),
        .M_AXIMM_109_AWADDR(M_AXIMM_109_AWADDR),
        .M_AXIMM_109_AWLEN(M_AXIMM_109_AWLEN),
        .M_AXIMM_109_AWSIZE(M_AXIMM_109_AWSIZE),
        .M_AXIMM_109_AWBURST(M_AXIMM_109_AWBURST),
        .M_AXIMM_109_AWLOCK(M_AXIMM_109_AWLOCK),
        .M_AXIMM_109_AWCACHE(M_AXIMM_109_AWCACHE),
        .M_AXIMM_109_AWPROT(M_AXIMM_109_AWPROT),
        .M_AXIMM_109_AWREGION(M_AXIMM_109_AWREGION),
        .M_AXIMM_109_AWQOS(M_AXIMM_109_AWQOS),
        .M_AXIMM_109_AWVALID(M_AXIMM_109_AWVALID),
        .M_AXIMM_109_AWREADY(M_AXIMM_109_AWREADY),
        .M_AXIMM_109_WDATA(M_AXIMM_109_WDATA),
        .M_AXIMM_109_WSTRB(M_AXIMM_109_WSTRB),
        .M_AXIMM_109_WLAST(M_AXIMM_109_WLAST),
        .M_AXIMM_109_WVALID(M_AXIMM_109_WVALID),
        .M_AXIMM_109_WREADY(M_AXIMM_109_WREADY),
        .M_AXIMM_109_BRESP(M_AXIMM_109_BRESP),
        .M_AXIMM_109_BVALID(M_AXIMM_109_BVALID),
        .M_AXIMM_109_BREADY(M_AXIMM_109_BREADY),
        .M_AXIMM_109_ARADDR(M_AXIMM_109_ARADDR),
        .M_AXIMM_109_ARLEN(M_AXIMM_109_ARLEN),
        .M_AXIMM_109_ARSIZE(M_AXIMM_109_ARSIZE),
        .M_AXIMM_109_ARBURST(M_AXIMM_109_ARBURST),
        .M_AXIMM_109_ARLOCK(M_AXIMM_109_ARLOCK),
        .M_AXIMM_109_ARCACHE(M_AXIMM_109_ARCACHE),
        .M_AXIMM_109_ARPROT(M_AXIMM_109_ARPROT),
        .M_AXIMM_109_ARREGION(M_AXIMM_109_ARREGION),
        .M_AXIMM_109_ARQOS(M_AXIMM_109_ARQOS),
        .M_AXIMM_109_ARVALID(M_AXIMM_109_ARVALID),
        .M_AXIMM_109_ARREADY(M_AXIMM_109_ARREADY),
        .M_AXIMM_109_RDATA(M_AXIMM_109_RDATA),
        .M_AXIMM_109_RRESP(M_AXIMM_109_RRESP),
        .M_AXIMM_109_RLAST(M_AXIMM_109_RLAST),
        .M_AXIMM_109_RVALID(M_AXIMM_109_RVALID),
        .M_AXIMM_109_RREADY(M_AXIMM_109_RREADY),
        .AP_AXIMM_110_AWADDR(AP_AXIMM_110_AWADDR),
        .AP_AXIMM_110_AWLEN(AP_AXIMM_110_AWLEN),
        .AP_AXIMM_110_AWSIZE(AP_AXIMM_110_AWSIZE),
        .AP_AXIMM_110_AWBURST(AP_AXIMM_110_AWBURST),
        .AP_AXIMM_110_AWLOCK(AP_AXIMM_110_AWLOCK),
        .AP_AXIMM_110_AWCACHE(AP_AXIMM_110_AWCACHE),
        .AP_AXIMM_110_AWPROT(AP_AXIMM_110_AWPROT),
        .AP_AXIMM_110_AWREGION(AP_AXIMM_110_AWREGION),
        .AP_AXIMM_110_AWQOS(AP_AXIMM_110_AWQOS),
        .AP_AXIMM_110_AWVALID(AP_AXIMM_110_AWVALID),
        .AP_AXIMM_110_AWREADY(AP_AXIMM_110_AWREADY),
        .AP_AXIMM_110_WDATA(AP_AXIMM_110_WDATA),
        .AP_AXIMM_110_WSTRB(AP_AXIMM_110_WSTRB),
        .AP_AXIMM_110_WLAST(AP_AXIMM_110_WLAST),
        .AP_AXIMM_110_WVALID(AP_AXIMM_110_WVALID),
        .AP_AXIMM_110_WREADY(AP_AXIMM_110_WREADY),
        .AP_AXIMM_110_BRESP(AP_AXIMM_110_BRESP),
        .AP_AXIMM_110_BVALID(AP_AXIMM_110_BVALID),
        .AP_AXIMM_110_BREADY(AP_AXIMM_110_BREADY),
        .AP_AXIMM_110_ARADDR(AP_AXIMM_110_ARADDR),
        .AP_AXIMM_110_ARLEN(AP_AXIMM_110_ARLEN),
        .AP_AXIMM_110_ARSIZE(AP_AXIMM_110_ARSIZE),
        .AP_AXIMM_110_ARBURST(AP_AXIMM_110_ARBURST),
        .AP_AXIMM_110_ARLOCK(AP_AXIMM_110_ARLOCK),
        .AP_AXIMM_110_ARCACHE(AP_AXIMM_110_ARCACHE),
        .AP_AXIMM_110_ARPROT(AP_AXIMM_110_ARPROT),
        .AP_AXIMM_110_ARREGION(AP_AXIMM_110_ARREGION),
        .AP_AXIMM_110_ARQOS(AP_AXIMM_110_ARQOS),
        .AP_AXIMM_110_ARVALID(AP_AXIMM_110_ARVALID),
        .AP_AXIMM_110_ARREADY(AP_AXIMM_110_ARREADY),
        .AP_AXIMM_110_RDATA(AP_AXIMM_110_RDATA),
        .AP_AXIMM_110_RRESP(AP_AXIMM_110_RRESP),
        .AP_AXIMM_110_RLAST(AP_AXIMM_110_RLAST),
        .AP_AXIMM_110_RVALID(AP_AXIMM_110_RVALID),
        .AP_AXIMM_110_RREADY(AP_AXIMM_110_RREADY),
        .M_AXIMM_110_AWADDR(M_AXIMM_110_AWADDR),
        .M_AXIMM_110_AWLEN(M_AXIMM_110_AWLEN),
        .M_AXIMM_110_AWSIZE(M_AXIMM_110_AWSIZE),
        .M_AXIMM_110_AWBURST(M_AXIMM_110_AWBURST),
        .M_AXIMM_110_AWLOCK(M_AXIMM_110_AWLOCK),
        .M_AXIMM_110_AWCACHE(M_AXIMM_110_AWCACHE),
        .M_AXIMM_110_AWPROT(M_AXIMM_110_AWPROT),
        .M_AXIMM_110_AWREGION(M_AXIMM_110_AWREGION),
        .M_AXIMM_110_AWQOS(M_AXIMM_110_AWQOS),
        .M_AXIMM_110_AWVALID(M_AXIMM_110_AWVALID),
        .M_AXIMM_110_AWREADY(M_AXIMM_110_AWREADY),
        .M_AXIMM_110_WDATA(M_AXIMM_110_WDATA),
        .M_AXIMM_110_WSTRB(M_AXIMM_110_WSTRB),
        .M_AXIMM_110_WLAST(M_AXIMM_110_WLAST),
        .M_AXIMM_110_WVALID(M_AXIMM_110_WVALID),
        .M_AXIMM_110_WREADY(M_AXIMM_110_WREADY),
        .M_AXIMM_110_BRESP(M_AXIMM_110_BRESP),
        .M_AXIMM_110_BVALID(M_AXIMM_110_BVALID),
        .M_AXIMM_110_BREADY(M_AXIMM_110_BREADY),
        .M_AXIMM_110_ARADDR(M_AXIMM_110_ARADDR),
        .M_AXIMM_110_ARLEN(M_AXIMM_110_ARLEN),
        .M_AXIMM_110_ARSIZE(M_AXIMM_110_ARSIZE),
        .M_AXIMM_110_ARBURST(M_AXIMM_110_ARBURST),
        .M_AXIMM_110_ARLOCK(M_AXIMM_110_ARLOCK),
        .M_AXIMM_110_ARCACHE(M_AXIMM_110_ARCACHE),
        .M_AXIMM_110_ARPROT(M_AXIMM_110_ARPROT),
        .M_AXIMM_110_ARREGION(M_AXIMM_110_ARREGION),
        .M_AXIMM_110_ARQOS(M_AXIMM_110_ARQOS),
        .M_AXIMM_110_ARVALID(M_AXIMM_110_ARVALID),
        .M_AXIMM_110_ARREADY(M_AXIMM_110_ARREADY),
        .M_AXIMM_110_RDATA(M_AXIMM_110_RDATA),
        .M_AXIMM_110_RRESP(M_AXIMM_110_RRESP),
        .M_AXIMM_110_RLAST(M_AXIMM_110_RLAST),
        .M_AXIMM_110_RVALID(M_AXIMM_110_RVALID),
        .M_AXIMM_110_RREADY(M_AXIMM_110_RREADY),
        .AP_AXIMM_111_AWADDR(AP_AXIMM_111_AWADDR),
        .AP_AXIMM_111_AWLEN(AP_AXIMM_111_AWLEN),
        .AP_AXIMM_111_AWSIZE(AP_AXIMM_111_AWSIZE),
        .AP_AXIMM_111_AWBURST(AP_AXIMM_111_AWBURST),
        .AP_AXIMM_111_AWLOCK(AP_AXIMM_111_AWLOCK),
        .AP_AXIMM_111_AWCACHE(AP_AXIMM_111_AWCACHE),
        .AP_AXIMM_111_AWPROT(AP_AXIMM_111_AWPROT),
        .AP_AXIMM_111_AWREGION(AP_AXIMM_111_AWREGION),
        .AP_AXIMM_111_AWQOS(AP_AXIMM_111_AWQOS),
        .AP_AXIMM_111_AWVALID(AP_AXIMM_111_AWVALID),
        .AP_AXIMM_111_AWREADY(AP_AXIMM_111_AWREADY),
        .AP_AXIMM_111_WDATA(AP_AXIMM_111_WDATA),
        .AP_AXIMM_111_WSTRB(AP_AXIMM_111_WSTRB),
        .AP_AXIMM_111_WLAST(AP_AXIMM_111_WLAST),
        .AP_AXIMM_111_WVALID(AP_AXIMM_111_WVALID),
        .AP_AXIMM_111_WREADY(AP_AXIMM_111_WREADY),
        .AP_AXIMM_111_BRESP(AP_AXIMM_111_BRESP),
        .AP_AXIMM_111_BVALID(AP_AXIMM_111_BVALID),
        .AP_AXIMM_111_BREADY(AP_AXIMM_111_BREADY),
        .AP_AXIMM_111_ARADDR(AP_AXIMM_111_ARADDR),
        .AP_AXIMM_111_ARLEN(AP_AXIMM_111_ARLEN),
        .AP_AXIMM_111_ARSIZE(AP_AXIMM_111_ARSIZE),
        .AP_AXIMM_111_ARBURST(AP_AXIMM_111_ARBURST),
        .AP_AXIMM_111_ARLOCK(AP_AXIMM_111_ARLOCK),
        .AP_AXIMM_111_ARCACHE(AP_AXIMM_111_ARCACHE),
        .AP_AXIMM_111_ARPROT(AP_AXIMM_111_ARPROT),
        .AP_AXIMM_111_ARREGION(AP_AXIMM_111_ARREGION),
        .AP_AXIMM_111_ARQOS(AP_AXIMM_111_ARQOS),
        .AP_AXIMM_111_ARVALID(AP_AXIMM_111_ARVALID),
        .AP_AXIMM_111_ARREADY(AP_AXIMM_111_ARREADY),
        .AP_AXIMM_111_RDATA(AP_AXIMM_111_RDATA),
        .AP_AXIMM_111_RRESP(AP_AXIMM_111_RRESP),
        .AP_AXIMM_111_RLAST(AP_AXIMM_111_RLAST),
        .AP_AXIMM_111_RVALID(AP_AXIMM_111_RVALID),
        .AP_AXIMM_111_RREADY(AP_AXIMM_111_RREADY),
        .M_AXIMM_111_AWADDR(M_AXIMM_111_AWADDR),
        .M_AXIMM_111_AWLEN(M_AXIMM_111_AWLEN),
        .M_AXIMM_111_AWSIZE(M_AXIMM_111_AWSIZE),
        .M_AXIMM_111_AWBURST(M_AXIMM_111_AWBURST),
        .M_AXIMM_111_AWLOCK(M_AXIMM_111_AWLOCK),
        .M_AXIMM_111_AWCACHE(M_AXIMM_111_AWCACHE),
        .M_AXIMM_111_AWPROT(M_AXIMM_111_AWPROT),
        .M_AXIMM_111_AWREGION(M_AXIMM_111_AWREGION),
        .M_AXIMM_111_AWQOS(M_AXIMM_111_AWQOS),
        .M_AXIMM_111_AWVALID(M_AXIMM_111_AWVALID),
        .M_AXIMM_111_AWREADY(M_AXIMM_111_AWREADY),
        .M_AXIMM_111_WDATA(M_AXIMM_111_WDATA),
        .M_AXIMM_111_WSTRB(M_AXIMM_111_WSTRB),
        .M_AXIMM_111_WLAST(M_AXIMM_111_WLAST),
        .M_AXIMM_111_WVALID(M_AXIMM_111_WVALID),
        .M_AXIMM_111_WREADY(M_AXIMM_111_WREADY),
        .M_AXIMM_111_BRESP(M_AXIMM_111_BRESP),
        .M_AXIMM_111_BVALID(M_AXIMM_111_BVALID),
        .M_AXIMM_111_BREADY(M_AXIMM_111_BREADY),
        .M_AXIMM_111_ARADDR(M_AXIMM_111_ARADDR),
        .M_AXIMM_111_ARLEN(M_AXIMM_111_ARLEN),
        .M_AXIMM_111_ARSIZE(M_AXIMM_111_ARSIZE),
        .M_AXIMM_111_ARBURST(M_AXIMM_111_ARBURST),
        .M_AXIMM_111_ARLOCK(M_AXIMM_111_ARLOCK),
        .M_AXIMM_111_ARCACHE(M_AXIMM_111_ARCACHE),
        .M_AXIMM_111_ARPROT(M_AXIMM_111_ARPROT),
        .M_AXIMM_111_ARREGION(M_AXIMM_111_ARREGION),
        .M_AXIMM_111_ARQOS(M_AXIMM_111_ARQOS),
        .M_AXIMM_111_ARVALID(M_AXIMM_111_ARVALID),
        .M_AXIMM_111_ARREADY(M_AXIMM_111_ARREADY),
        .M_AXIMM_111_RDATA(M_AXIMM_111_RDATA),
        .M_AXIMM_111_RRESP(M_AXIMM_111_RRESP),
        .M_AXIMM_111_RLAST(M_AXIMM_111_RLAST),
        .M_AXIMM_111_RVALID(M_AXIMM_111_RVALID),
        .M_AXIMM_111_RREADY(M_AXIMM_111_RREADY),
        .AP_AXIMM_112_AWADDR(AP_AXIMM_112_AWADDR),
        .AP_AXIMM_112_AWLEN(AP_AXIMM_112_AWLEN),
        .AP_AXIMM_112_AWSIZE(AP_AXIMM_112_AWSIZE),
        .AP_AXIMM_112_AWBURST(AP_AXIMM_112_AWBURST),
        .AP_AXIMM_112_AWLOCK(AP_AXIMM_112_AWLOCK),
        .AP_AXIMM_112_AWCACHE(AP_AXIMM_112_AWCACHE),
        .AP_AXIMM_112_AWPROT(AP_AXIMM_112_AWPROT),
        .AP_AXIMM_112_AWREGION(AP_AXIMM_112_AWREGION),
        .AP_AXIMM_112_AWQOS(AP_AXIMM_112_AWQOS),
        .AP_AXIMM_112_AWVALID(AP_AXIMM_112_AWVALID),
        .AP_AXIMM_112_AWREADY(AP_AXIMM_112_AWREADY),
        .AP_AXIMM_112_WDATA(AP_AXIMM_112_WDATA),
        .AP_AXIMM_112_WSTRB(AP_AXIMM_112_WSTRB),
        .AP_AXIMM_112_WLAST(AP_AXIMM_112_WLAST),
        .AP_AXIMM_112_WVALID(AP_AXIMM_112_WVALID),
        .AP_AXIMM_112_WREADY(AP_AXIMM_112_WREADY),
        .AP_AXIMM_112_BRESP(AP_AXIMM_112_BRESP),
        .AP_AXIMM_112_BVALID(AP_AXIMM_112_BVALID),
        .AP_AXIMM_112_BREADY(AP_AXIMM_112_BREADY),
        .AP_AXIMM_112_ARADDR(AP_AXIMM_112_ARADDR),
        .AP_AXIMM_112_ARLEN(AP_AXIMM_112_ARLEN),
        .AP_AXIMM_112_ARSIZE(AP_AXIMM_112_ARSIZE),
        .AP_AXIMM_112_ARBURST(AP_AXIMM_112_ARBURST),
        .AP_AXIMM_112_ARLOCK(AP_AXIMM_112_ARLOCK),
        .AP_AXIMM_112_ARCACHE(AP_AXIMM_112_ARCACHE),
        .AP_AXIMM_112_ARPROT(AP_AXIMM_112_ARPROT),
        .AP_AXIMM_112_ARREGION(AP_AXIMM_112_ARREGION),
        .AP_AXIMM_112_ARQOS(AP_AXIMM_112_ARQOS),
        .AP_AXIMM_112_ARVALID(AP_AXIMM_112_ARVALID),
        .AP_AXIMM_112_ARREADY(AP_AXIMM_112_ARREADY),
        .AP_AXIMM_112_RDATA(AP_AXIMM_112_RDATA),
        .AP_AXIMM_112_RRESP(AP_AXIMM_112_RRESP),
        .AP_AXIMM_112_RLAST(AP_AXIMM_112_RLAST),
        .AP_AXIMM_112_RVALID(AP_AXIMM_112_RVALID),
        .AP_AXIMM_112_RREADY(AP_AXIMM_112_RREADY),
        .M_AXIMM_112_AWADDR(M_AXIMM_112_AWADDR),
        .M_AXIMM_112_AWLEN(M_AXIMM_112_AWLEN),
        .M_AXIMM_112_AWSIZE(M_AXIMM_112_AWSIZE),
        .M_AXIMM_112_AWBURST(M_AXIMM_112_AWBURST),
        .M_AXIMM_112_AWLOCK(M_AXIMM_112_AWLOCK),
        .M_AXIMM_112_AWCACHE(M_AXIMM_112_AWCACHE),
        .M_AXIMM_112_AWPROT(M_AXIMM_112_AWPROT),
        .M_AXIMM_112_AWREGION(M_AXIMM_112_AWREGION),
        .M_AXIMM_112_AWQOS(M_AXIMM_112_AWQOS),
        .M_AXIMM_112_AWVALID(M_AXIMM_112_AWVALID),
        .M_AXIMM_112_AWREADY(M_AXIMM_112_AWREADY),
        .M_AXIMM_112_WDATA(M_AXIMM_112_WDATA),
        .M_AXIMM_112_WSTRB(M_AXIMM_112_WSTRB),
        .M_AXIMM_112_WLAST(M_AXIMM_112_WLAST),
        .M_AXIMM_112_WVALID(M_AXIMM_112_WVALID),
        .M_AXIMM_112_WREADY(M_AXIMM_112_WREADY),
        .M_AXIMM_112_BRESP(M_AXIMM_112_BRESP),
        .M_AXIMM_112_BVALID(M_AXIMM_112_BVALID),
        .M_AXIMM_112_BREADY(M_AXIMM_112_BREADY),
        .M_AXIMM_112_ARADDR(M_AXIMM_112_ARADDR),
        .M_AXIMM_112_ARLEN(M_AXIMM_112_ARLEN),
        .M_AXIMM_112_ARSIZE(M_AXIMM_112_ARSIZE),
        .M_AXIMM_112_ARBURST(M_AXIMM_112_ARBURST),
        .M_AXIMM_112_ARLOCK(M_AXIMM_112_ARLOCK),
        .M_AXIMM_112_ARCACHE(M_AXIMM_112_ARCACHE),
        .M_AXIMM_112_ARPROT(M_AXIMM_112_ARPROT),
        .M_AXIMM_112_ARREGION(M_AXIMM_112_ARREGION),
        .M_AXIMM_112_ARQOS(M_AXIMM_112_ARQOS),
        .M_AXIMM_112_ARVALID(M_AXIMM_112_ARVALID),
        .M_AXIMM_112_ARREADY(M_AXIMM_112_ARREADY),
        .M_AXIMM_112_RDATA(M_AXIMM_112_RDATA),
        .M_AXIMM_112_RRESP(M_AXIMM_112_RRESP),
        .M_AXIMM_112_RLAST(M_AXIMM_112_RLAST),
        .M_AXIMM_112_RVALID(M_AXIMM_112_RVALID),
        .M_AXIMM_112_RREADY(M_AXIMM_112_RREADY),
        .AP_AXIMM_113_AWADDR(AP_AXIMM_113_AWADDR),
        .AP_AXIMM_113_AWLEN(AP_AXIMM_113_AWLEN),
        .AP_AXIMM_113_AWSIZE(AP_AXIMM_113_AWSIZE),
        .AP_AXIMM_113_AWBURST(AP_AXIMM_113_AWBURST),
        .AP_AXIMM_113_AWLOCK(AP_AXIMM_113_AWLOCK),
        .AP_AXIMM_113_AWCACHE(AP_AXIMM_113_AWCACHE),
        .AP_AXIMM_113_AWPROT(AP_AXIMM_113_AWPROT),
        .AP_AXIMM_113_AWREGION(AP_AXIMM_113_AWREGION),
        .AP_AXIMM_113_AWQOS(AP_AXIMM_113_AWQOS),
        .AP_AXIMM_113_AWVALID(AP_AXIMM_113_AWVALID),
        .AP_AXIMM_113_AWREADY(AP_AXIMM_113_AWREADY),
        .AP_AXIMM_113_WDATA(AP_AXIMM_113_WDATA),
        .AP_AXIMM_113_WSTRB(AP_AXIMM_113_WSTRB),
        .AP_AXIMM_113_WLAST(AP_AXIMM_113_WLAST),
        .AP_AXIMM_113_WVALID(AP_AXIMM_113_WVALID),
        .AP_AXIMM_113_WREADY(AP_AXIMM_113_WREADY),
        .AP_AXIMM_113_BRESP(AP_AXIMM_113_BRESP),
        .AP_AXIMM_113_BVALID(AP_AXIMM_113_BVALID),
        .AP_AXIMM_113_BREADY(AP_AXIMM_113_BREADY),
        .AP_AXIMM_113_ARADDR(AP_AXIMM_113_ARADDR),
        .AP_AXIMM_113_ARLEN(AP_AXIMM_113_ARLEN),
        .AP_AXIMM_113_ARSIZE(AP_AXIMM_113_ARSIZE),
        .AP_AXIMM_113_ARBURST(AP_AXIMM_113_ARBURST),
        .AP_AXIMM_113_ARLOCK(AP_AXIMM_113_ARLOCK),
        .AP_AXIMM_113_ARCACHE(AP_AXIMM_113_ARCACHE),
        .AP_AXIMM_113_ARPROT(AP_AXIMM_113_ARPROT),
        .AP_AXIMM_113_ARREGION(AP_AXIMM_113_ARREGION),
        .AP_AXIMM_113_ARQOS(AP_AXIMM_113_ARQOS),
        .AP_AXIMM_113_ARVALID(AP_AXIMM_113_ARVALID),
        .AP_AXIMM_113_ARREADY(AP_AXIMM_113_ARREADY),
        .AP_AXIMM_113_RDATA(AP_AXIMM_113_RDATA),
        .AP_AXIMM_113_RRESP(AP_AXIMM_113_RRESP),
        .AP_AXIMM_113_RLAST(AP_AXIMM_113_RLAST),
        .AP_AXIMM_113_RVALID(AP_AXIMM_113_RVALID),
        .AP_AXIMM_113_RREADY(AP_AXIMM_113_RREADY),
        .M_AXIMM_113_AWADDR(M_AXIMM_113_AWADDR),
        .M_AXIMM_113_AWLEN(M_AXIMM_113_AWLEN),
        .M_AXIMM_113_AWSIZE(M_AXIMM_113_AWSIZE),
        .M_AXIMM_113_AWBURST(M_AXIMM_113_AWBURST),
        .M_AXIMM_113_AWLOCK(M_AXIMM_113_AWLOCK),
        .M_AXIMM_113_AWCACHE(M_AXIMM_113_AWCACHE),
        .M_AXIMM_113_AWPROT(M_AXIMM_113_AWPROT),
        .M_AXIMM_113_AWREGION(M_AXIMM_113_AWREGION),
        .M_AXIMM_113_AWQOS(M_AXIMM_113_AWQOS),
        .M_AXIMM_113_AWVALID(M_AXIMM_113_AWVALID),
        .M_AXIMM_113_AWREADY(M_AXIMM_113_AWREADY),
        .M_AXIMM_113_WDATA(M_AXIMM_113_WDATA),
        .M_AXIMM_113_WSTRB(M_AXIMM_113_WSTRB),
        .M_AXIMM_113_WLAST(M_AXIMM_113_WLAST),
        .M_AXIMM_113_WVALID(M_AXIMM_113_WVALID),
        .M_AXIMM_113_WREADY(M_AXIMM_113_WREADY),
        .M_AXIMM_113_BRESP(M_AXIMM_113_BRESP),
        .M_AXIMM_113_BVALID(M_AXIMM_113_BVALID),
        .M_AXIMM_113_BREADY(M_AXIMM_113_BREADY),
        .M_AXIMM_113_ARADDR(M_AXIMM_113_ARADDR),
        .M_AXIMM_113_ARLEN(M_AXIMM_113_ARLEN),
        .M_AXIMM_113_ARSIZE(M_AXIMM_113_ARSIZE),
        .M_AXIMM_113_ARBURST(M_AXIMM_113_ARBURST),
        .M_AXIMM_113_ARLOCK(M_AXIMM_113_ARLOCK),
        .M_AXIMM_113_ARCACHE(M_AXIMM_113_ARCACHE),
        .M_AXIMM_113_ARPROT(M_AXIMM_113_ARPROT),
        .M_AXIMM_113_ARREGION(M_AXIMM_113_ARREGION),
        .M_AXIMM_113_ARQOS(M_AXIMM_113_ARQOS),
        .M_AXIMM_113_ARVALID(M_AXIMM_113_ARVALID),
        .M_AXIMM_113_ARREADY(M_AXIMM_113_ARREADY),
        .M_AXIMM_113_RDATA(M_AXIMM_113_RDATA),
        .M_AXIMM_113_RRESP(M_AXIMM_113_RRESP),
        .M_AXIMM_113_RLAST(M_AXIMM_113_RLAST),
        .M_AXIMM_113_RVALID(M_AXIMM_113_RVALID),
        .M_AXIMM_113_RREADY(M_AXIMM_113_RREADY),
        .AP_AXIMM_114_AWADDR(AP_AXIMM_114_AWADDR),
        .AP_AXIMM_114_AWLEN(AP_AXIMM_114_AWLEN),
        .AP_AXIMM_114_AWSIZE(AP_AXIMM_114_AWSIZE),
        .AP_AXIMM_114_AWBURST(AP_AXIMM_114_AWBURST),
        .AP_AXIMM_114_AWLOCK(AP_AXIMM_114_AWLOCK),
        .AP_AXIMM_114_AWCACHE(AP_AXIMM_114_AWCACHE),
        .AP_AXIMM_114_AWPROT(AP_AXIMM_114_AWPROT),
        .AP_AXIMM_114_AWREGION(AP_AXIMM_114_AWREGION),
        .AP_AXIMM_114_AWQOS(AP_AXIMM_114_AWQOS),
        .AP_AXIMM_114_AWVALID(AP_AXIMM_114_AWVALID),
        .AP_AXIMM_114_AWREADY(AP_AXIMM_114_AWREADY),
        .AP_AXIMM_114_WDATA(AP_AXIMM_114_WDATA),
        .AP_AXIMM_114_WSTRB(AP_AXIMM_114_WSTRB),
        .AP_AXIMM_114_WLAST(AP_AXIMM_114_WLAST),
        .AP_AXIMM_114_WVALID(AP_AXIMM_114_WVALID),
        .AP_AXIMM_114_WREADY(AP_AXIMM_114_WREADY),
        .AP_AXIMM_114_BRESP(AP_AXIMM_114_BRESP),
        .AP_AXIMM_114_BVALID(AP_AXIMM_114_BVALID),
        .AP_AXIMM_114_BREADY(AP_AXIMM_114_BREADY),
        .AP_AXIMM_114_ARADDR(AP_AXIMM_114_ARADDR),
        .AP_AXIMM_114_ARLEN(AP_AXIMM_114_ARLEN),
        .AP_AXIMM_114_ARSIZE(AP_AXIMM_114_ARSIZE),
        .AP_AXIMM_114_ARBURST(AP_AXIMM_114_ARBURST),
        .AP_AXIMM_114_ARLOCK(AP_AXIMM_114_ARLOCK),
        .AP_AXIMM_114_ARCACHE(AP_AXIMM_114_ARCACHE),
        .AP_AXIMM_114_ARPROT(AP_AXIMM_114_ARPROT),
        .AP_AXIMM_114_ARREGION(AP_AXIMM_114_ARREGION),
        .AP_AXIMM_114_ARQOS(AP_AXIMM_114_ARQOS),
        .AP_AXIMM_114_ARVALID(AP_AXIMM_114_ARVALID),
        .AP_AXIMM_114_ARREADY(AP_AXIMM_114_ARREADY),
        .AP_AXIMM_114_RDATA(AP_AXIMM_114_RDATA),
        .AP_AXIMM_114_RRESP(AP_AXIMM_114_RRESP),
        .AP_AXIMM_114_RLAST(AP_AXIMM_114_RLAST),
        .AP_AXIMM_114_RVALID(AP_AXIMM_114_RVALID),
        .AP_AXIMM_114_RREADY(AP_AXIMM_114_RREADY),
        .M_AXIMM_114_AWADDR(M_AXIMM_114_AWADDR),
        .M_AXIMM_114_AWLEN(M_AXIMM_114_AWLEN),
        .M_AXIMM_114_AWSIZE(M_AXIMM_114_AWSIZE),
        .M_AXIMM_114_AWBURST(M_AXIMM_114_AWBURST),
        .M_AXIMM_114_AWLOCK(M_AXIMM_114_AWLOCK),
        .M_AXIMM_114_AWCACHE(M_AXIMM_114_AWCACHE),
        .M_AXIMM_114_AWPROT(M_AXIMM_114_AWPROT),
        .M_AXIMM_114_AWREGION(M_AXIMM_114_AWREGION),
        .M_AXIMM_114_AWQOS(M_AXIMM_114_AWQOS),
        .M_AXIMM_114_AWVALID(M_AXIMM_114_AWVALID),
        .M_AXIMM_114_AWREADY(M_AXIMM_114_AWREADY),
        .M_AXIMM_114_WDATA(M_AXIMM_114_WDATA),
        .M_AXIMM_114_WSTRB(M_AXIMM_114_WSTRB),
        .M_AXIMM_114_WLAST(M_AXIMM_114_WLAST),
        .M_AXIMM_114_WVALID(M_AXIMM_114_WVALID),
        .M_AXIMM_114_WREADY(M_AXIMM_114_WREADY),
        .M_AXIMM_114_BRESP(M_AXIMM_114_BRESP),
        .M_AXIMM_114_BVALID(M_AXIMM_114_BVALID),
        .M_AXIMM_114_BREADY(M_AXIMM_114_BREADY),
        .M_AXIMM_114_ARADDR(M_AXIMM_114_ARADDR),
        .M_AXIMM_114_ARLEN(M_AXIMM_114_ARLEN),
        .M_AXIMM_114_ARSIZE(M_AXIMM_114_ARSIZE),
        .M_AXIMM_114_ARBURST(M_AXIMM_114_ARBURST),
        .M_AXIMM_114_ARLOCK(M_AXIMM_114_ARLOCK),
        .M_AXIMM_114_ARCACHE(M_AXIMM_114_ARCACHE),
        .M_AXIMM_114_ARPROT(M_AXIMM_114_ARPROT),
        .M_AXIMM_114_ARREGION(M_AXIMM_114_ARREGION),
        .M_AXIMM_114_ARQOS(M_AXIMM_114_ARQOS),
        .M_AXIMM_114_ARVALID(M_AXIMM_114_ARVALID),
        .M_AXIMM_114_ARREADY(M_AXIMM_114_ARREADY),
        .M_AXIMM_114_RDATA(M_AXIMM_114_RDATA),
        .M_AXIMM_114_RRESP(M_AXIMM_114_RRESP),
        .M_AXIMM_114_RLAST(M_AXIMM_114_RLAST),
        .M_AXIMM_114_RVALID(M_AXIMM_114_RVALID),
        .M_AXIMM_114_RREADY(M_AXIMM_114_RREADY),
        .AP_AXIMM_115_AWADDR(AP_AXIMM_115_AWADDR),
        .AP_AXIMM_115_AWLEN(AP_AXIMM_115_AWLEN),
        .AP_AXIMM_115_AWSIZE(AP_AXIMM_115_AWSIZE),
        .AP_AXIMM_115_AWBURST(AP_AXIMM_115_AWBURST),
        .AP_AXIMM_115_AWLOCK(AP_AXIMM_115_AWLOCK),
        .AP_AXIMM_115_AWCACHE(AP_AXIMM_115_AWCACHE),
        .AP_AXIMM_115_AWPROT(AP_AXIMM_115_AWPROT),
        .AP_AXIMM_115_AWREGION(AP_AXIMM_115_AWREGION),
        .AP_AXIMM_115_AWQOS(AP_AXIMM_115_AWQOS),
        .AP_AXIMM_115_AWVALID(AP_AXIMM_115_AWVALID),
        .AP_AXIMM_115_AWREADY(AP_AXIMM_115_AWREADY),
        .AP_AXIMM_115_WDATA(AP_AXIMM_115_WDATA),
        .AP_AXIMM_115_WSTRB(AP_AXIMM_115_WSTRB),
        .AP_AXIMM_115_WLAST(AP_AXIMM_115_WLAST),
        .AP_AXIMM_115_WVALID(AP_AXIMM_115_WVALID),
        .AP_AXIMM_115_WREADY(AP_AXIMM_115_WREADY),
        .AP_AXIMM_115_BRESP(AP_AXIMM_115_BRESP),
        .AP_AXIMM_115_BVALID(AP_AXIMM_115_BVALID),
        .AP_AXIMM_115_BREADY(AP_AXIMM_115_BREADY),
        .AP_AXIMM_115_ARADDR(AP_AXIMM_115_ARADDR),
        .AP_AXIMM_115_ARLEN(AP_AXIMM_115_ARLEN),
        .AP_AXIMM_115_ARSIZE(AP_AXIMM_115_ARSIZE),
        .AP_AXIMM_115_ARBURST(AP_AXIMM_115_ARBURST),
        .AP_AXIMM_115_ARLOCK(AP_AXIMM_115_ARLOCK),
        .AP_AXIMM_115_ARCACHE(AP_AXIMM_115_ARCACHE),
        .AP_AXIMM_115_ARPROT(AP_AXIMM_115_ARPROT),
        .AP_AXIMM_115_ARREGION(AP_AXIMM_115_ARREGION),
        .AP_AXIMM_115_ARQOS(AP_AXIMM_115_ARQOS),
        .AP_AXIMM_115_ARVALID(AP_AXIMM_115_ARVALID),
        .AP_AXIMM_115_ARREADY(AP_AXIMM_115_ARREADY),
        .AP_AXIMM_115_RDATA(AP_AXIMM_115_RDATA),
        .AP_AXIMM_115_RRESP(AP_AXIMM_115_RRESP),
        .AP_AXIMM_115_RLAST(AP_AXIMM_115_RLAST),
        .AP_AXIMM_115_RVALID(AP_AXIMM_115_RVALID),
        .AP_AXIMM_115_RREADY(AP_AXIMM_115_RREADY),
        .M_AXIMM_115_AWADDR(M_AXIMM_115_AWADDR),
        .M_AXIMM_115_AWLEN(M_AXIMM_115_AWLEN),
        .M_AXIMM_115_AWSIZE(M_AXIMM_115_AWSIZE),
        .M_AXIMM_115_AWBURST(M_AXIMM_115_AWBURST),
        .M_AXIMM_115_AWLOCK(M_AXIMM_115_AWLOCK),
        .M_AXIMM_115_AWCACHE(M_AXIMM_115_AWCACHE),
        .M_AXIMM_115_AWPROT(M_AXIMM_115_AWPROT),
        .M_AXIMM_115_AWREGION(M_AXIMM_115_AWREGION),
        .M_AXIMM_115_AWQOS(M_AXIMM_115_AWQOS),
        .M_AXIMM_115_AWVALID(M_AXIMM_115_AWVALID),
        .M_AXIMM_115_AWREADY(M_AXIMM_115_AWREADY),
        .M_AXIMM_115_WDATA(M_AXIMM_115_WDATA),
        .M_AXIMM_115_WSTRB(M_AXIMM_115_WSTRB),
        .M_AXIMM_115_WLAST(M_AXIMM_115_WLAST),
        .M_AXIMM_115_WVALID(M_AXIMM_115_WVALID),
        .M_AXIMM_115_WREADY(M_AXIMM_115_WREADY),
        .M_AXIMM_115_BRESP(M_AXIMM_115_BRESP),
        .M_AXIMM_115_BVALID(M_AXIMM_115_BVALID),
        .M_AXIMM_115_BREADY(M_AXIMM_115_BREADY),
        .M_AXIMM_115_ARADDR(M_AXIMM_115_ARADDR),
        .M_AXIMM_115_ARLEN(M_AXIMM_115_ARLEN),
        .M_AXIMM_115_ARSIZE(M_AXIMM_115_ARSIZE),
        .M_AXIMM_115_ARBURST(M_AXIMM_115_ARBURST),
        .M_AXIMM_115_ARLOCK(M_AXIMM_115_ARLOCK),
        .M_AXIMM_115_ARCACHE(M_AXIMM_115_ARCACHE),
        .M_AXIMM_115_ARPROT(M_AXIMM_115_ARPROT),
        .M_AXIMM_115_ARREGION(M_AXIMM_115_ARREGION),
        .M_AXIMM_115_ARQOS(M_AXIMM_115_ARQOS),
        .M_AXIMM_115_ARVALID(M_AXIMM_115_ARVALID),
        .M_AXIMM_115_ARREADY(M_AXIMM_115_ARREADY),
        .M_AXIMM_115_RDATA(M_AXIMM_115_RDATA),
        .M_AXIMM_115_RRESP(M_AXIMM_115_RRESP),
        .M_AXIMM_115_RLAST(M_AXIMM_115_RLAST),
        .M_AXIMM_115_RVALID(M_AXIMM_115_RVALID),
        .M_AXIMM_115_RREADY(M_AXIMM_115_RREADY),
        .AP_AXIMM_116_AWADDR(AP_AXIMM_116_AWADDR),
        .AP_AXIMM_116_AWLEN(AP_AXIMM_116_AWLEN),
        .AP_AXIMM_116_AWSIZE(AP_AXIMM_116_AWSIZE),
        .AP_AXIMM_116_AWBURST(AP_AXIMM_116_AWBURST),
        .AP_AXIMM_116_AWLOCK(AP_AXIMM_116_AWLOCK),
        .AP_AXIMM_116_AWCACHE(AP_AXIMM_116_AWCACHE),
        .AP_AXIMM_116_AWPROT(AP_AXIMM_116_AWPROT),
        .AP_AXIMM_116_AWREGION(AP_AXIMM_116_AWREGION),
        .AP_AXIMM_116_AWQOS(AP_AXIMM_116_AWQOS),
        .AP_AXIMM_116_AWVALID(AP_AXIMM_116_AWVALID),
        .AP_AXIMM_116_AWREADY(AP_AXIMM_116_AWREADY),
        .AP_AXIMM_116_WDATA(AP_AXIMM_116_WDATA),
        .AP_AXIMM_116_WSTRB(AP_AXIMM_116_WSTRB),
        .AP_AXIMM_116_WLAST(AP_AXIMM_116_WLAST),
        .AP_AXIMM_116_WVALID(AP_AXIMM_116_WVALID),
        .AP_AXIMM_116_WREADY(AP_AXIMM_116_WREADY),
        .AP_AXIMM_116_BRESP(AP_AXIMM_116_BRESP),
        .AP_AXIMM_116_BVALID(AP_AXIMM_116_BVALID),
        .AP_AXIMM_116_BREADY(AP_AXIMM_116_BREADY),
        .AP_AXIMM_116_ARADDR(AP_AXIMM_116_ARADDR),
        .AP_AXIMM_116_ARLEN(AP_AXIMM_116_ARLEN),
        .AP_AXIMM_116_ARSIZE(AP_AXIMM_116_ARSIZE),
        .AP_AXIMM_116_ARBURST(AP_AXIMM_116_ARBURST),
        .AP_AXIMM_116_ARLOCK(AP_AXIMM_116_ARLOCK),
        .AP_AXIMM_116_ARCACHE(AP_AXIMM_116_ARCACHE),
        .AP_AXIMM_116_ARPROT(AP_AXIMM_116_ARPROT),
        .AP_AXIMM_116_ARREGION(AP_AXIMM_116_ARREGION),
        .AP_AXIMM_116_ARQOS(AP_AXIMM_116_ARQOS),
        .AP_AXIMM_116_ARVALID(AP_AXIMM_116_ARVALID),
        .AP_AXIMM_116_ARREADY(AP_AXIMM_116_ARREADY),
        .AP_AXIMM_116_RDATA(AP_AXIMM_116_RDATA),
        .AP_AXIMM_116_RRESP(AP_AXIMM_116_RRESP),
        .AP_AXIMM_116_RLAST(AP_AXIMM_116_RLAST),
        .AP_AXIMM_116_RVALID(AP_AXIMM_116_RVALID),
        .AP_AXIMM_116_RREADY(AP_AXIMM_116_RREADY),
        .M_AXIMM_116_AWADDR(M_AXIMM_116_AWADDR),
        .M_AXIMM_116_AWLEN(M_AXIMM_116_AWLEN),
        .M_AXIMM_116_AWSIZE(M_AXIMM_116_AWSIZE),
        .M_AXIMM_116_AWBURST(M_AXIMM_116_AWBURST),
        .M_AXIMM_116_AWLOCK(M_AXIMM_116_AWLOCK),
        .M_AXIMM_116_AWCACHE(M_AXIMM_116_AWCACHE),
        .M_AXIMM_116_AWPROT(M_AXIMM_116_AWPROT),
        .M_AXIMM_116_AWREGION(M_AXIMM_116_AWREGION),
        .M_AXIMM_116_AWQOS(M_AXIMM_116_AWQOS),
        .M_AXIMM_116_AWVALID(M_AXIMM_116_AWVALID),
        .M_AXIMM_116_AWREADY(M_AXIMM_116_AWREADY),
        .M_AXIMM_116_WDATA(M_AXIMM_116_WDATA),
        .M_AXIMM_116_WSTRB(M_AXIMM_116_WSTRB),
        .M_AXIMM_116_WLAST(M_AXIMM_116_WLAST),
        .M_AXIMM_116_WVALID(M_AXIMM_116_WVALID),
        .M_AXIMM_116_WREADY(M_AXIMM_116_WREADY),
        .M_AXIMM_116_BRESP(M_AXIMM_116_BRESP),
        .M_AXIMM_116_BVALID(M_AXIMM_116_BVALID),
        .M_AXIMM_116_BREADY(M_AXIMM_116_BREADY),
        .M_AXIMM_116_ARADDR(M_AXIMM_116_ARADDR),
        .M_AXIMM_116_ARLEN(M_AXIMM_116_ARLEN),
        .M_AXIMM_116_ARSIZE(M_AXIMM_116_ARSIZE),
        .M_AXIMM_116_ARBURST(M_AXIMM_116_ARBURST),
        .M_AXIMM_116_ARLOCK(M_AXIMM_116_ARLOCK),
        .M_AXIMM_116_ARCACHE(M_AXIMM_116_ARCACHE),
        .M_AXIMM_116_ARPROT(M_AXIMM_116_ARPROT),
        .M_AXIMM_116_ARREGION(M_AXIMM_116_ARREGION),
        .M_AXIMM_116_ARQOS(M_AXIMM_116_ARQOS),
        .M_AXIMM_116_ARVALID(M_AXIMM_116_ARVALID),
        .M_AXIMM_116_ARREADY(M_AXIMM_116_ARREADY),
        .M_AXIMM_116_RDATA(M_AXIMM_116_RDATA),
        .M_AXIMM_116_RRESP(M_AXIMM_116_RRESP),
        .M_AXIMM_116_RLAST(M_AXIMM_116_RLAST),
        .M_AXIMM_116_RVALID(M_AXIMM_116_RVALID),
        .M_AXIMM_116_RREADY(M_AXIMM_116_RREADY),
        .AP_AXIMM_117_AWADDR(AP_AXIMM_117_AWADDR),
        .AP_AXIMM_117_AWLEN(AP_AXIMM_117_AWLEN),
        .AP_AXIMM_117_AWSIZE(AP_AXIMM_117_AWSIZE),
        .AP_AXIMM_117_AWBURST(AP_AXIMM_117_AWBURST),
        .AP_AXIMM_117_AWLOCK(AP_AXIMM_117_AWLOCK),
        .AP_AXIMM_117_AWCACHE(AP_AXIMM_117_AWCACHE),
        .AP_AXIMM_117_AWPROT(AP_AXIMM_117_AWPROT),
        .AP_AXIMM_117_AWREGION(AP_AXIMM_117_AWREGION),
        .AP_AXIMM_117_AWQOS(AP_AXIMM_117_AWQOS),
        .AP_AXIMM_117_AWVALID(AP_AXIMM_117_AWVALID),
        .AP_AXIMM_117_AWREADY(AP_AXIMM_117_AWREADY),
        .AP_AXIMM_117_WDATA(AP_AXIMM_117_WDATA),
        .AP_AXIMM_117_WSTRB(AP_AXIMM_117_WSTRB),
        .AP_AXIMM_117_WLAST(AP_AXIMM_117_WLAST),
        .AP_AXIMM_117_WVALID(AP_AXIMM_117_WVALID),
        .AP_AXIMM_117_WREADY(AP_AXIMM_117_WREADY),
        .AP_AXIMM_117_BRESP(AP_AXIMM_117_BRESP),
        .AP_AXIMM_117_BVALID(AP_AXIMM_117_BVALID),
        .AP_AXIMM_117_BREADY(AP_AXIMM_117_BREADY),
        .AP_AXIMM_117_ARADDR(AP_AXIMM_117_ARADDR),
        .AP_AXIMM_117_ARLEN(AP_AXIMM_117_ARLEN),
        .AP_AXIMM_117_ARSIZE(AP_AXIMM_117_ARSIZE),
        .AP_AXIMM_117_ARBURST(AP_AXIMM_117_ARBURST),
        .AP_AXIMM_117_ARLOCK(AP_AXIMM_117_ARLOCK),
        .AP_AXIMM_117_ARCACHE(AP_AXIMM_117_ARCACHE),
        .AP_AXIMM_117_ARPROT(AP_AXIMM_117_ARPROT),
        .AP_AXIMM_117_ARREGION(AP_AXIMM_117_ARREGION),
        .AP_AXIMM_117_ARQOS(AP_AXIMM_117_ARQOS),
        .AP_AXIMM_117_ARVALID(AP_AXIMM_117_ARVALID),
        .AP_AXIMM_117_ARREADY(AP_AXIMM_117_ARREADY),
        .AP_AXIMM_117_RDATA(AP_AXIMM_117_RDATA),
        .AP_AXIMM_117_RRESP(AP_AXIMM_117_RRESP),
        .AP_AXIMM_117_RLAST(AP_AXIMM_117_RLAST),
        .AP_AXIMM_117_RVALID(AP_AXIMM_117_RVALID),
        .AP_AXIMM_117_RREADY(AP_AXIMM_117_RREADY),
        .M_AXIMM_117_AWADDR(M_AXIMM_117_AWADDR),
        .M_AXIMM_117_AWLEN(M_AXIMM_117_AWLEN),
        .M_AXIMM_117_AWSIZE(M_AXIMM_117_AWSIZE),
        .M_AXIMM_117_AWBURST(M_AXIMM_117_AWBURST),
        .M_AXIMM_117_AWLOCK(M_AXIMM_117_AWLOCK),
        .M_AXIMM_117_AWCACHE(M_AXIMM_117_AWCACHE),
        .M_AXIMM_117_AWPROT(M_AXIMM_117_AWPROT),
        .M_AXIMM_117_AWREGION(M_AXIMM_117_AWREGION),
        .M_AXIMM_117_AWQOS(M_AXIMM_117_AWQOS),
        .M_AXIMM_117_AWVALID(M_AXIMM_117_AWVALID),
        .M_AXIMM_117_AWREADY(M_AXIMM_117_AWREADY),
        .M_AXIMM_117_WDATA(M_AXIMM_117_WDATA),
        .M_AXIMM_117_WSTRB(M_AXIMM_117_WSTRB),
        .M_AXIMM_117_WLAST(M_AXIMM_117_WLAST),
        .M_AXIMM_117_WVALID(M_AXIMM_117_WVALID),
        .M_AXIMM_117_WREADY(M_AXIMM_117_WREADY),
        .M_AXIMM_117_BRESP(M_AXIMM_117_BRESP),
        .M_AXIMM_117_BVALID(M_AXIMM_117_BVALID),
        .M_AXIMM_117_BREADY(M_AXIMM_117_BREADY),
        .M_AXIMM_117_ARADDR(M_AXIMM_117_ARADDR),
        .M_AXIMM_117_ARLEN(M_AXIMM_117_ARLEN),
        .M_AXIMM_117_ARSIZE(M_AXIMM_117_ARSIZE),
        .M_AXIMM_117_ARBURST(M_AXIMM_117_ARBURST),
        .M_AXIMM_117_ARLOCK(M_AXIMM_117_ARLOCK),
        .M_AXIMM_117_ARCACHE(M_AXIMM_117_ARCACHE),
        .M_AXIMM_117_ARPROT(M_AXIMM_117_ARPROT),
        .M_AXIMM_117_ARREGION(M_AXIMM_117_ARREGION),
        .M_AXIMM_117_ARQOS(M_AXIMM_117_ARQOS),
        .M_AXIMM_117_ARVALID(M_AXIMM_117_ARVALID),
        .M_AXIMM_117_ARREADY(M_AXIMM_117_ARREADY),
        .M_AXIMM_117_RDATA(M_AXIMM_117_RDATA),
        .M_AXIMM_117_RRESP(M_AXIMM_117_RRESP),
        .M_AXIMM_117_RLAST(M_AXIMM_117_RLAST),
        .M_AXIMM_117_RVALID(M_AXIMM_117_RVALID),
        .M_AXIMM_117_RREADY(M_AXIMM_117_RREADY),
        .AP_AXIMM_118_AWADDR(AP_AXIMM_118_AWADDR),
        .AP_AXIMM_118_AWLEN(AP_AXIMM_118_AWLEN),
        .AP_AXIMM_118_AWSIZE(AP_AXIMM_118_AWSIZE),
        .AP_AXIMM_118_AWBURST(AP_AXIMM_118_AWBURST),
        .AP_AXIMM_118_AWLOCK(AP_AXIMM_118_AWLOCK),
        .AP_AXIMM_118_AWCACHE(AP_AXIMM_118_AWCACHE),
        .AP_AXIMM_118_AWPROT(AP_AXIMM_118_AWPROT),
        .AP_AXIMM_118_AWREGION(AP_AXIMM_118_AWREGION),
        .AP_AXIMM_118_AWQOS(AP_AXIMM_118_AWQOS),
        .AP_AXIMM_118_AWVALID(AP_AXIMM_118_AWVALID),
        .AP_AXIMM_118_AWREADY(AP_AXIMM_118_AWREADY),
        .AP_AXIMM_118_WDATA(AP_AXIMM_118_WDATA),
        .AP_AXIMM_118_WSTRB(AP_AXIMM_118_WSTRB),
        .AP_AXIMM_118_WLAST(AP_AXIMM_118_WLAST),
        .AP_AXIMM_118_WVALID(AP_AXIMM_118_WVALID),
        .AP_AXIMM_118_WREADY(AP_AXIMM_118_WREADY),
        .AP_AXIMM_118_BRESP(AP_AXIMM_118_BRESP),
        .AP_AXIMM_118_BVALID(AP_AXIMM_118_BVALID),
        .AP_AXIMM_118_BREADY(AP_AXIMM_118_BREADY),
        .AP_AXIMM_118_ARADDR(AP_AXIMM_118_ARADDR),
        .AP_AXIMM_118_ARLEN(AP_AXIMM_118_ARLEN),
        .AP_AXIMM_118_ARSIZE(AP_AXIMM_118_ARSIZE),
        .AP_AXIMM_118_ARBURST(AP_AXIMM_118_ARBURST),
        .AP_AXIMM_118_ARLOCK(AP_AXIMM_118_ARLOCK),
        .AP_AXIMM_118_ARCACHE(AP_AXIMM_118_ARCACHE),
        .AP_AXIMM_118_ARPROT(AP_AXIMM_118_ARPROT),
        .AP_AXIMM_118_ARREGION(AP_AXIMM_118_ARREGION),
        .AP_AXIMM_118_ARQOS(AP_AXIMM_118_ARQOS),
        .AP_AXIMM_118_ARVALID(AP_AXIMM_118_ARVALID),
        .AP_AXIMM_118_ARREADY(AP_AXIMM_118_ARREADY),
        .AP_AXIMM_118_RDATA(AP_AXIMM_118_RDATA),
        .AP_AXIMM_118_RRESP(AP_AXIMM_118_RRESP),
        .AP_AXIMM_118_RLAST(AP_AXIMM_118_RLAST),
        .AP_AXIMM_118_RVALID(AP_AXIMM_118_RVALID),
        .AP_AXIMM_118_RREADY(AP_AXIMM_118_RREADY),
        .M_AXIMM_118_AWADDR(M_AXIMM_118_AWADDR),
        .M_AXIMM_118_AWLEN(M_AXIMM_118_AWLEN),
        .M_AXIMM_118_AWSIZE(M_AXIMM_118_AWSIZE),
        .M_AXIMM_118_AWBURST(M_AXIMM_118_AWBURST),
        .M_AXIMM_118_AWLOCK(M_AXIMM_118_AWLOCK),
        .M_AXIMM_118_AWCACHE(M_AXIMM_118_AWCACHE),
        .M_AXIMM_118_AWPROT(M_AXIMM_118_AWPROT),
        .M_AXIMM_118_AWREGION(M_AXIMM_118_AWREGION),
        .M_AXIMM_118_AWQOS(M_AXIMM_118_AWQOS),
        .M_AXIMM_118_AWVALID(M_AXIMM_118_AWVALID),
        .M_AXIMM_118_AWREADY(M_AXIMM_118_AWREADY),
        .M_AXIMM_118_WDATA(M_AXIMM_118_WDATA),
        .M_AXIMM_118_WSTRB(M_AXIMM_118_WSTRB),
        .M_AXIMM_118_WLAST(M_AXIMM_118_WLAST),
        .M_AXIMM_118_WVALID(M_AXIMM_118_WVALID),
        .M_AXIMM_118_WREADY(M_AXIMM_118_WREADY),
        .M_AXIMM_118_BRESP(M_AXIMM_118_BRESP),
        .M_AXIMM_118_BVALID(M_AXIMM_118_BVALID),
        .M_AXIMM_118_BREADY(M_AXIMM_118_BREADY),
        .M_AXIMM_118_ARADDR(M_AXIMM_118_ARADDR),
        .M_AXIMM_118_ARLEN(M_AXIMM_118_ARLEN),
        .M_AXIMM_118_ARSIZE(M_AXIMM_118_ARSIZE),
        .M_AXIMM_118_ARBURST(M_AXIMM_118_ARBURST),
        .M_AXIMM_118_ARLOCK(M_AXIMM_118_ARLOCK),
        .M_AXIMM_118_ARCACHE(M_AXIMM_118_ARCACHE),
        .M_AXIMM_118_ARPROT(M_AXIMM_118_ARPROT),
        .M_AXIMM_118_ARREGION(M_AXIMM_118_ARREGION),
        .M_AXIMM_118_ARQOS(M_AXIMM_118_ARQOS),
        .M_AXIMM_118_ARVALID(M_AXIMM_118_ARVALID),
        .M_AXIMM_118_ARREADY(M_AXIMM_118_ARREADY),
        .M_AXIMM_118_RDATA(M_AXIMM_118_RDATA),
        .M_AXIMM_118_RRESP(M_AXIMM_118_RRESP),
        .M_AXIMM_118_RLAST(M_AXIMM_118_RLAST),
        .M_AXIMM_118_RVALID(M_AXIMM_118_RVALID),
        .M_AXIMM_118_RREADY(M_AXIMM_118_RREADY),
        .AP_AXIMM_119_AWADDR(AP_AXIMM_119_AWADDR),
        .AP_AXIMM_119_AWLEN(AP_AXIMM_119_AWLEN),
        .AP_AXIMM_119_AWSIZE(AP_AXIMM_119_AWSIZE),
        .AP_AXIMM_119_AWBURST(AP_AXIMM_119_AWBURST),
        .AP_AXIMM_119_AWLOCK(AP_AXIMM_119_AWLOCK),
        .AP_AXIMM_119_AWCACHE(AP_AXIMM_119_AWCACHE),
        .AP_AXIMM_119_AWPROT(AP_AXIMM_119_AWPROT),
        .AP_AXIMM_119_AWREGION(AP_AXIMM_119_AWREGION),
        .AP_AXIMM_119_AWQOS(AP_AXIMM_119_AWQOS),
        .AP_AXIMM_119_AWVALID(AP_AXIMM_119_AWVALID),
        .AP_AXIMM_119_AWREADY(AP_AXIMM_119_AWREADY),
        .AP_AXIMM_119_WDATA(AP_AXIMM_119_WDATA),
        .AP_AXIMM_119_WSTRB(AP_AXIMM_119_WSTRB),
        .AP_AXIMM_119_WLAST(AP_AXIMM_119_WLAST),
        .AP_AXIMM_119_WVALID(AP_AXIMM_119_WVALID),
        .AP_AXIMM_119_WREADY(AP_AXIMM_119_WREADY),
        .AP_AXIMM_119_BRESP(AP_AXIMM_119_BRESP),
        .AP_AXIMM_119_BVALID(AP_AXIMM_119_BVALID),
        .AP_AXIMM_119_BREADY(AP_AXIMM_119_BREADY),
        .AP_AXIMM_119_ARADDR(AP_AXIMM_119_ARADDR),
        .AP_AXIMM_119_ARLEN(AP_AXIMM_119_ARLEN),
        .AP_AXIMM_119_ARSIZE(AP_AXIMM_119_ARSIZE),
        .AP_AXIMM_119_ARBURST(AP_AXIMM_119_ARBURST),
        .AP_AXIMM_119_ARLOCK(AP_AXIMM_119_ARLOCK),
        .AP_AXIMM_119_ARCACHE(AP_AXIMM_119_ARCACHE),
        .AP_AXIMM_119_ARPROT(AP_AXIMM_119_ARPROT),
        .AP_AXIMM_119_ARREGION(AP_AXIMM_119_ARREGION),
        .AP_AXIMM_119_ARQOS(AP_AXIMM_119_ARQOS),
        .AP_AXIMM_119_ARVALID(AP_AXIMM_119_ARVALID),
        .AP_AXIMM_119_ARREADY(AP_AXIMM_119_ARREADY),
        .AP_AXIMM_119_RDATA(AP_AXIMM_119_RDATA),
        .AP_AXIMM_119_RRESP(AP_AXIMM_119_RRESP),
        .AP_AXIMM_119_RLAST(AP_AXIMM_119_RLAST),
        .AP_AXIMM_119_RVALID(AP_AXIMM_119_RVALID),
        .AP_AXIMM_119_RREADY(AP_AXIMM_119_RREADY),
        .M_AXIMM_119_AWADDR(M_AXIMM_119_AWADDR),
        .M_AXIMM_119_AWLEN(M_AXIMM_119_AWLEN),
        .M_AXIMM_119_AWSIZE(M_AXIMM_119_AWSIZE),
        .M_AXIMM_119_AWBURST(M_AXIMM_119_AWBURST),
        .M_AXIMM_119_AWLOCK(M_AXIMM_119_AWLOCK),
        .M_AXIMM_119_AWCACHE(M_AXIMM_119_AWCACHE),
        .M_AXIMM_119_AWPROT(M_AXIMM_119_AWPROT),
        .M_AXIMM_119_AWREGION(M_AXIMM_119_AWREGION),
        .M_AXIMM_119_AWQOS(M_AXIMM_119_AWQOS),
        .M_AXIMM_119_AWVALID(M_AXIMM_119_AWVALID),
        .M_AXIMM_119_AWREADY(M_AXIMM_119_AWREADY),
        .M_AXIMM_119_WDATA(M_AXIMM_119_WDATA),
        .M_AXIMM_119_WSTRB(M_AXIMM_119_WSTRB),
        .M_AXIMM_119_WLAST(M_AXIMM_119_WLAST),
        .M_AXIMM_119_WVALID(M_AXIMM_119_WVALID),
        .M_AXIMM_119_WREADY(M_AXIMM_119_WREADY),
        .M_AXIMM_119_BRESP(M_AXIMM_119_BRESP),
        .M_AXIMM_119_BVALID(M_AXIMM_119_BVALID),
        .M_AXIMM_119_BREADY(M_AXIMM_119_BREADY),
        .M_AXIMM_119_ARADDR(M_AXIMM_119_ARADDR),
        .M_AXIMM_119_ARLEN(M_AXIMM_119_ARLEN),
        .M_AXIMM_119_ARSIZE(M_AXIMM_119_ARSIZE),
        .M_AXIMM_119_ARBURST(M_AXIMM_119_ARBURST),
        .M_AXIMM_119_ARLOCK(M_AXIMM_119_ARLOCK),
        .M_AXIMM_119_ARCACHE(M_AXIMM_119_ARCACHE),
        .M_AXIMM_119_ARPROT(M_AXIMM_119_ARPROT),
        .M_AXIMM_119_ARREGION(M_AXIMM_119_ARREGION),
        .M_AXIMM_119_ARQOS(M_AXIMM_119_ARQOS),
        .M_AXIMM_119_ARVALID(M_AXIMM_119_ARVALID),
        .M_AXIMM_119_ARREADY(M_AXIMM_119_ARREADY),
        .M_AXIMM_119_RDATA(M_AXIMM_119_RDATA),
        .M_AXIMM_119_RRESP(M_AXIMM_119_RRESP),
        .M_AXIMM_119_RLAST(M_AXIMM_119_RLAST),
        .M_AXIMM_119_RVALID(M_AXIMM_119_RVALID),
        .M_AXIMM_119_RREADY(M_AXIMM_119_RREADY),
        .AP_AXIMM_120_AWADDR(AP_AXIMM_120_AWADDR),
        .AP_AXIMM_120_AWLEN(AP_AXIMM_120_AWLEN),
        .AP_AXIMM_120_AWSIZE(AP_AXIMM_120_AWSIZE),
        .AP_AXIMM_120_AWBURST(AP_AXIMM_120_AWBURST),
        .AP_AXIMM_120_AWLOCK(AP_AXIMM_120_AWLOCK),
        .AP_AXIMM_120_AWCACHE(AP_AXIMM_120_AWCACHE),
        .AP_AXIMM_120_AWPROT(AP_AXIMM_120_AWPROT),
        .AP_AXIMM_120_AWREGION(AP_AXIMM_120_AWREGION),
        .AP_AXIMM_120_AWQOS(AP_AXIMM_120_AWQOS),
        .AP_AXIMM_120_AWVALID(AP_AXIMM_120_AWVALID),
        .AP_AXIMM_120_AWREADY(AP_AXIMM_120_AWREADY),
        .AP_AXIMM_120_WDATA(AP_AXIMM_120_WDATA),
        .AP_AXIMM_120_WSTRB(AP_AXIMM_120_WSTRB),
        .AP_AXIMM_120_WLAST(AP_AXIMM_120_WLAST),
        .AP_AXIMM_120_WVALID(AP_AXIMM_120_WVALID),
        .AP_AXIMM_120_WREADY(AP_AXIMM_120_WREADY),
        .AP_AXIMM_120_BRESP(AP_AXIMM_120_BRESP),
        .AP_AXIMM_120_BVALID(AP_AXIMM_120_BVALID),
        .AP_AXIMM_120_BREADY(AP_AXIMM_120_BREADY),
        .AP_AXIMM_120_ARADDR(AP_AXIMM_120_ARADDR),
        .AP_AXIMM_120_ARLEN(AP_AXIMM_120_ARLEN),
        .AP_AXIMM_120_ARSIZE(AP_AXIMM_120_ARSIZE),
        .AP_AXIMM_120_ARBURST(AP_AXIMM_120_ARBURST),
        .AP_AXIMM_120_ARLOCK(AP_AXIMM_120_ARLOCK),
        .AP_AXIMM_120_ARCACHE(AP_AXIMM_120_ARCACHE),
        .AP_AXIMM_120_ARPROT(AP_AXIMM_120_ARPROT),
        .AP_AXIMM_120_ARREGION(AP_AXIMM_120_ARREGION),
        .AP_AXIMM_120_ARQOS(AP_AXIMM_120_ARQOS),
        .AP_AXIMM_120_ARVALID(AP_AXIMM_120_ARVALID),
        .AP_AXIMM_120_ARREADY(AP_AXIMM_120_ARREADY),
        .AP_AXIMM_120_RDATA(AP_AXIMM_120_RDATA),
        .AP_AXIMM_120_RRESP(AP_AXIMM_120_RRESP),
        .AP_AXIMM_120_RLAST(AP_AXIMM_120_RLAST),
        .AP_AXIMM_120_RVALID(AP_AXIMM_120_RVALID),
        .AP_AXIMM_120_RREADY(AP_AXIMM_120_RREADY),
        .M_AXIMM_120_AWADDR(M_AXIMM_120_AWADDR),
        .M_AXIMM_120_AWLEN(M_AXIMM_120_AWLEN),
        .M_AXIMM_120_AWSIZE(M_AXIMM_120_AWSIZE),
        .M_AXIMM_120_AWBURST(M_AXIMM_120_AWBURST),
        .M_AXIMM_120_AWLOCK(M_AXIMM_120_AWLOCK),
        .M_AXIMM_120_AWCACHE(M_AXIMM_120_AWCACHE),
        .M_AXIMM_120_AWPROT(M_AXIMM_120_AWPROT),
        .M_AXIMM_120_AWREGION(M_AXIMM_120_AWREGION),
        .M_AXIMM_120_AWQOS(M_AXIMM_120_AWQOS),
        .M_AXIMM_120_AWVALID(M_AXIMM_120_AWVALID),
        .M_AXIMM_120_AWREADY(M_AXIMM_120_AWREADY),
        .M_AXIMM_120_WDATA(M_AXIMM_120_WDATA),
        .M_AXIMM_120_WSTRB(M_AXIMM_120_WSTRB),
        .M_AXIMM_120_WLAST(M_AXIMM_120_WLAST),
        .M_AXIMM_120_WVALID(M_AXIMM_120_WVALID),
        .M_AXIMM_120_WREADY(M_AXIMM_120_WREADY),
        .M_AXIMM_120_BRESP(M_AXIMM_120_BRESP),
        .M_AXIMM_120_BVALID(M_AXIMM_120_BVALID),
        .M_AXIMM_120_BREADY(M_AXIMM_120_BREADY),
        .M_AXIMM_120_ARADDR(M_AXIMM_120_ARADDR),
        .M_AXIMM_120_ARLEN(M_AXIMM_120_ARLEN),
        .M_AXIMM_120_ARSIZE(M_AXIMM_120_ARSIZE),
        .M_AXIMM_120_ARBURST(M_AXIMM_120_ARBURST),
        .M_AXIMM_120_ARLOCK(M_AXIMM_120_ARLOCK),
        .M_AXIMM_120_ARCACHE(M_AXIMM_120_ARCACHE),
        .M_AXIMM_120_ARPROT(M_AXIMM_120_ARPROT),
        .M_AXIMM_120_ARREGION(M_AXIMM_120_ARREGION),
        .M_AXIMM_120_ARQOS(M_AXIMM_120_ARQOS),
        .M_AXIMM_120_ARVALID(M_AXIMM_120_ARVALID),
        .M_AXIMM_120_ARREADY(M_AXIMM_120_ARREADY),
        .M_AXIMM_120_RDATA(M_AXIMM_120_RDATA),
        .M_AXIMM_120_RRESP(M_AXIMM_120_RRESP),
        .M_AXIMM_120_RLAST(M_AXIMM_120_RLAST),
        .M_AXIMM_120_RVALID(M_AXIMM_120_RVALID),
        .M_AXIMM_120_RREADY(M_AXIMM_120_RREADY),
        .AP_AXIMM_121_AWADDR(AP_AXIMM_121_AWADDR),
        .AP_AXIMM_121_AWLEN(AP_AXIMM_121_AWLEN),
        .AP_AXIMM_121_AWSIZE(AP_AXIMM_121_AWSIZE),
        .AP_AXIMM_121_AWBURST(AP_AXIMM_121_AWBURST),
        .AP_AXIMM_121_AWLOCK(AP_AXIMM_121_AWLOCK),
        .AP_AXIMM_121_AWCACHE(AP_AXIMM_121_AWCACHE),
        .AP_AXIMM_121_AWPROT(AP_AXIMM_121_AWPROT),
        .AP_AXIMM_121_AWREGION(AP_AXIMM_121_AWREGION),
        .AP_AXIMM_121_AWQOS(AP_AXIMM_121_AWQOS),
        .AP_AXIMM_121_AWVALID(AP_AXIMM_121_AWVALID),
        .AP_AXIMM_121_AWREADY(AP_AXIMM_121_AWREADY),
        .AP_AXIMM_121_WDATA(AP_AXIMM_121_WDATA),
        .AP_AXIMM_121_WSTRB(AP_AXIMM_121_WSTRB),
        .AP_AXIMM_121_WLAST(AP_AXIMM_121_WLAST),
        .AP_AXIMM_121_WVALID(AP_AXIMM_121_WVALID),
        .AP_AXIMM_121_WREADY(AP_AXIMM_121_WREADY),
        .AP_AXIMM_121_BRESP(AP_AXIMM_121_BRESP),
        .AP_AXIMM_121_BVALID(AP_AXIMM_121_BVALID),
        .AP_AXIMM_121_BREADY(AP_AXIMM_121_BREADY),
        .AP_AXIMM_121_ARADDR(AP_AXIMM_121_ARADDR),
        .AP_AXIMM_121_ARLEN(AP_AXIMM_121_ARLEN),
        .AP_AXIMM_121_ARSIZE(AP_AXIMM_121_ARSIZE),
        .AP_AXIMM_121_ARBURST(AP_AXIMM_121_ARBURST),
        .AP_AXIMM_121_ARLOCK(AP_AXIMM_121_ARLOCK),
        .AP_AXIMM_121_ARCACHE(AP_AXIMM_121_ARCACHE),
        .AP_AXIMM_121_ARPROT(AP_AXIMM_121_ARPROT),
        .AP_AXIMM_121_ARREGION(AP_AXIMM_121_ARREGION),
        .AP_AXIMM_121_ARQOS(AP_AXIMM_121_ARQOS),
        .AP_AXIMM_121_ARVALID(AP_AXIMM_121_ARVALID),
        .AP_AXIMM_121_ARREADY(AP_AXIMM_121_ARREADY),
        .AP_AXIMM_121_RDATA(AP_AXIMM_121_RDATA),
        .AP_AXIMM_121_RRESP(AP_AXIMM_121_RRESP),
        .AP_AXIMM_121_RLAST(AP_AXIMM_121_RLAST),
        .AP_AXIMM_121_RVALID(AP_AXIMM_121_RVALID),
        .AP_AXIMM_121_RREADY(AP_AXIMM_121_RREADY),
        .M_AXIMM_121_AWADDR(M_AXIMM_121_AWADDR),
        .M_AXIMM_121_AWLEN(M_AXIMM_121_AWLEN),
        .M_AXIMM_121_AWSIZE(M_AXIMM_121_AWSIZE),
        .M_AXIMM_121_AWBURST(M_AXIMM_121_AWBURST),
        .M_AXIMM_121_AWLOCK(M_AXIMM_121_AWLOCK),
        .M_AXIMM_121_AWCACHE(M_AXIMM_121_AWCACHE),
        .M_AXIMM_121_AWPROT(M_AXIMM_121_AWPROT),
        .M_AXIMM_121_AWREGION(M_AXIMM_121_AWREGION),
        .M_AXIMM_121_AWQOS(M_AXIMM_121_AWQOS),
        .M_AXIMM_121_AWVALID(M_AXIMM_121_AWVALID),
        .M_AXIMM_121_AWREADY(M_AXIMM_121_AWREADY),
        .M_AXIMM_121_WDATA(M_AXIMM_121_WDATA),
        .M_AXIMM_121_WSTRB(M_AXIMM_121_WSTRB),
        .M_AXIMM_121_WLAST(M_AXIMM_121_WLAST),
        .M_AXIMM_121_WVALID(M_AXIMM_121_WVALID),
        .M_AXIMM_121_WREADY(M_AXIMM_121_WREADY),
        .M_AXIMM_121_BRESP(M_AXIMM_121_BRESP),
        .M_AXIMM_121_BVALID(M_AXIMM_121_BVALID),
        .M_AXIMM_121_BREADY(M_AXIMM_121_BREADY),
        .M_AXIMM_121_ARADDR(M_AXIMM_121_ARADDR),
        .M_AXIMM_121_ARLEN(M_AXIMM_121_ARLEN),
        .M_AXIMM_121_ARSIZE(M_AXIMM_121_ARSIZE),
        .M_AXIMM_121_ARBURST(M_AXIMM_121_ARBURST),
        .M_AXIMM_121_ARLOCK(M_AXIMM_121_ARLOCK),
        .M_AXIMM_121_ARCACHE(M_AXIMM_121_ARCACHE),
        .M_AXIMM_121_ARPROT(M_AXIMM_121_ARPROT),
        .M_AXIMM_121_ARREGION(M_AXIMM_121_ARREGION),
        .M_AXIMM_121_ARQOS(M_AXIMM_121_ARQOS),
        .M_AXIMM_121_ARVALID(M_AXIMM_121_ARVALID),
        .M_AXIMM_121_ARREADY(M_AXIMM_121_ARREADY),
        .M_AXIMM_121_RDATA(M_AXIMM_121_RDATA),
        .M_AXIMM_121_RRESP(M_AXIMM_121_RRESP),
        .M_AXIMM_121_RLAST(M_AXIMM_121_RLAST),
        .M_AXIMM_121_RVALID(M_AXIMM_121_RVALID),
        .M_AXIMM_121_RREADY(M_AXIMM_121_RREADY),
        .AP_AXIMM_122_AWADDR(AP_AXIMM_122_AWADDR),
        .AP_AXIMM_122_AWLEN(AP_AXIMM_122_AWLEN),
        .AP_AXIMM_122_AWSIZE(AP_AXIMM_122_AWSIZE),
        .AP_AXIMM_122_AWBURST(AP_AXIMM_122_AWBURST),
        .AP_AXIMM_122_AWLOCK(AP_AXIMM_122_AWLOCK),
        .AP_AXIMM_122_AWCACHE(AP_AXIMM_122_AWCACHE),
        .AP_AXIMM_122_AWPROT(AP_AXIMM_122_AWPROT),
        .AP_AXIMM_122_AWREGION(AP_AXIMM_122_AWREGION),
        .AP_AXIMM_122_AWQOS(AP_AXIMM_122_AWQOS),
        .AP_AXIMM_122_AWVALID(AP_AXIMM_122_AWVALID),
        .AP_AXIMM_122_AWREADY(AP_AXIMM_122_AWREADY),
        .AP_AXIMM_122_WDATA(AP_AXIMM_122_WDATA),
        .AP_AXIMM_122_WSTRB(AP_AXIMM_122_WSTRB),
        .AP_AXIMM_122_WLAST(AP_AXIMM_122_WLAST),
        .AP_AXIMM_122_WVALID(AP_AXIMM_122_WVALID),
        .AP_AXIMM_122_WREADY(AP_AXIMM_122_WREADY),
        .AP_AXIMM_122_BRESP(AP_AXIMM_122_BRESP),
        .AP_AXIMM_122_BVALID(AP_AXIMM_122_BVALID),
        .AP_AXIMM_122_BREADY(AP_AXIMM_122_BREADY),
        .AP_AXIMM_122_ARADDR(AP_AXIMM_122_ARADDR),
        .AP_AXIMM_122_ARLEN(AP_AXIMM_122_ARLEN),
        .AP_AXIMM_122_ARSIZE(AP_AXIMM_122_ARSIZE),
        .AP_AXIMM_122_ARBURST(AP_AXIMM_122_ARBURST),
        .AP_AXIMM_122_ARLOCK(AP_AXIMM_122_ARLOCK),
        .AP_AXIMM_122_ARCACHE(AP_AXIMM_122_ARCACHE),
        .AP_AXIMM_122_ARPROT(AP_AXIMM_122_ARPROT),
        .AP_AXIMM_122_ARREGION(AP_AXIMM_122_ARREGION),
        .AP_AXIMM_122_ARQOS(AP_AXIMM_122_ARQOS),
        .AP_AXIMM_122_ARVALID(AP_AXIMM_122_ARVALID),
        .AP_AXIMM_122_ARREADY(AP_AXIMM_122_ARREADY),
        .AP_AXIMM_122_RDATA(AP_AXIMM_122_RDATA),
        .AP_AXIMM_122_RRESP(AP_AXIMM_122_RRESP),
        .AP_AXIMM_122_RLAST(AP_AXIMM_122_RLAST),
        .AP_AXIMM_122_RVALID(AP_AXIMM_122_RVALID),
        .AP_AXIMM_122_RREADY(AP_AXIMM_122_RREADY),
        .M_AXIMM_122_AWADDR(M_AXIMM_122_AWADDR),
        .M_AXIMM_122_AWLEN(M_AXIMM_122_AWLEN),
        .M_AXIMM_122_AWSIZE(M_AXIMM_122_AWSIZE),
        .M_AXIMM_122_AWBURST(M_AXIMM_122_AWBURST),
        .M_AXIMM_122_AWLOCK(M_AXIMM_122_AWLOCK),
        .M_AXIMM_122_AWCACHE(M_AXIMM_122_AWCACHE),
        .M_AXIMM_122_AWPROT(M_AXIMM_122_AWPROT),
        .M_AXIMM_122_AWREGION(M_AXIMM_122_AWREGION),
        .M_AXIMM_122_AWQOS(M_AXIMM_122_AWQOS),
        .M_AXIMM_122_AWVALID(M_AXIMM_122_AWVALID),
        .M_AXIMM_122_AWREADY(M_AXIMM_122_AWREADY),
        .M_AXIMM_122_WDATA(M_AXIMM_122_WDATA),
        .M_AXIMM_122_WSTRB(M_AXIMM_122_WSTRB),
        .M_AXIMM_122_WLAST(M_AXIMM_122_WLAST),
        .M_AXIMM_122_WVALID(M_AXIMM_122_WVALID),
        .M_AXIMM_122_WREADY(M_AXIMM_122_WREADY),
        .M_AXIMM_122_BRESP(M_AXIMM_122_BRESP),
        .M_AXIMM_122_BVALID(M_AXIMM_122_BVALID),
        .M_AXIMM_122_BREADY(M_AXIMM_122_BREADY),
        .M_AXIMM_122_ARADDR(M_AXIMM_122_ARADDR),
        .M_AXIMM_122_ARLEN(M_AXIMM_122_ARLEN),
        .M_AXIMM_122_ARSIZE(M_AXIMM_122_ARSIZE),
        .M_AXIMM_122_ARBURST(M_AXIMM_122_ARBURST),
        .M_AXIMM_122_ARLOCK(M_AXIMM_122_ARLOCK),
        .M_AXIMM_122_ARCACHE(M_AXIMM_122_ARCACHE),
        .M_AXIMM_122_ARPROT(M_AXIMM_122_ARPROT),
        .M_AXIMM_122_ARREGION(M_AXIMM_122_ARREGION),
        .M_AXIMM_122_ARQOS(M_AXIMM_122_ARQOS),
        .M_AXIMM_122_ARVALID(M_AXIMM_122_ARVALID),
        .M_AXIMM_122_ARREADY(M_AXIMM_122_ARREADY),
        .M_AXIMM_122_RDATA(M_AXIMM_122_RDATA),
        .M_AXIMM_122_RRESP(M_AXIMM_122_RRESP),
        .M_AXIMM_122_RLAST(M_AXIMM_122_RLAST),
        .M_AXIMM_122_RVALID(M_AXIMM_122_RVALID),
        .M_AXIMM_122_RREADY(M_AXIMM_122_RREADY),
        .AP_AXIMM_123_AWADDR(AP_AXIMM_123_AWADDR),
        .AP_AXIMM_123_AWLEN(AP_AXIMM_123_AWLEN),
        .AP_AXIMM_123_AWSIZE(AP_AXIMM_123_AWSIZE),
        .AP_AXIMM_123_AWBURST(AP_AXIMM_123_AWBURST),
        .AP_AXIMM_123_AWLOCK(AP_AXIMM_123_AWLOCK),
        .AP_AXIMM_123_AWCACHE(AP_AXIMM_123_AWCACHE),
        .AP_AXIMM_123_AWPROT(AP_AXIMM_123_AWPROT),
        .AP_AXIMM_123_AWREGION(AP_AXIMM_123_AWREGION),
        .AP_AXIMM_123_AWQOS(AP_AXIMM_123_AWQOS),
        .AP_AXIMM_123_AWVALID(AP_AXIMM_123_AWVALID),
        .AP_AXIMM_123_AWREADY(AP_AXIMM_123_AWREADY),
        .AP_AXIMM_123_WDATA(AP_AXIMM_123_WDATA),
        .AP_AXIMM_123_WSTRB(AP_AXIMM_123_WSTRB),
        .AP_AXIMM_123_WLAST(AP_AXIMM_123_WLAST),
        .AP_AXIMM_123_WVALID(AP_AXIMM_123_WVALID),
        .AP_AXIMM_123_WREADY(AP_AXIMM_123_WREADY),
        .AP_AXIMM_123_BRESP(AP_AXIMM_123_BRESP),
        .AP_AXIMM_123_BVALID(AP_AXIMM_123_BVALID),
        .AP_AXIMM_123_BREADY(AP_AXIMM_123_BREADY),
        .AP_AXIMM_123_ARADDR(AP_AXIMM_123_ARADDR),
        .AP_AXIMM_123_ARLEN(AP_AXIMM_123_ARLEN),
        .AP_AXIMM_123_ARSIZE(AP_AXIMM_123_ARSIZE),
        .AP_AXIMM_123_ARBURST(AP_AXIMM_123_ARBURST),
        .AP_AXIMM_123_ARLOCK(AP_AXIMM_123_ARLOCK),
        .AP_AXIMM_123_ARCACHE(AP_AXIMM_123_ARCACHE),
        .AP_AXIMM_123_ARPROT(AP_AXIMM_123_ARPROT),
        .AP_AXIMM_123_ARREGION(AP_AXIMM_123_ARREGION),
        .AP_AXIMM_123_ARQOS(AP_AXIMM_123_ARQOS),
        .AP_AXIMM_123_ARVALID(AP_AXIMM_123_ARVALID),
        .AP_AXIMM_123_ARREADY(AP_AXIMM_123_ARREADY),
        .AP_AXIMM_123_RDATA(AP_AXIMM_123_RDATA),
        .AP_AXIMM_123_RRESP(AP_AXIMM_123_RRESP),
        .AP_AXIMM_123_RLAST(AP_AXIMM_123_RLAST),
        .AP_AXIMM_123_RVALID(AP_AXIMM_123_RVALID),
        .AP_AXIMM_123_RREADY(AP_AXIMM_123_RREADY),
        .M_AXIMM_123_AWADDR(M_AXIMM_123_AWADDR),
        .M_AXIMM_123_AWLEN(M_AXIMM_123_AWLEN),
        .M_AXIMM_123_AWSIZE(M_AXIMM_123_AWSIZE),
        .M_AXIMM_123_AWBURST(M_AXIMM_123_AWBURST),
        .M_AXIMM_123_AWLOCK(M_AXIMM_123_AWLOCK),
        .M_AXIMM_123_AWCACHE(M_AXIMM_123_AWCACHE),
        .M_AXIMM_123_AWPROT(M_AXIMM_123_AWPROT),
        .M_AXIMM_123_AWREGION(M_AXIMM_123_AWREGION),
        .M_AXIMM_123_AWQOS(M_AXIMM_123_AWQOS),
        .M_AXIMM_123_AWVALID(M_AXIMM_123_AWVALID),
        .M_AXIMM_123_AWREADY(M_AXIMM_123_AWREADY),
        .M_AXIMM_123_WDATA(M_AXIMM_123_WDATA),
        .M_AXIMM_123_WSTRB(M_AXIMM_123_WSTRB),
        .M_AXIMM_123_WLAST(M_AXIMM_123_WLAST),
        .M_AXIMM_123_WVALID(M_AXIMM_123_WVALID),
        .M_AXIMM_123_WREADY(M_AXIMM_123_WREADY),
        .M_AXIMM_123_BRESP(M_AXIMM_123_BRESP),
        .M_AXIMM_123_BVALID(M_AXIMM_123_BVALID),
        .M_AXIMM_123_BREADY(M_AXIMM_123_BREADY),
        .M_AXIMM_123_ARADDR(M_AXIMM_123_ARADDR),
        .M_AXIMM_123_ARLEN(M_AXIMM_123_ARLEN),
        .M_AXIMM_123_ARSIZE(M_AXIMM_123_ARSIZE),
        .M_AXIMM_123_ARBURST(M_AXIMM_123_ARBURST),
        .M_AXIMM_123_ARLOCK(M_AXIMM_123_ARLOCK),
        .M_AXIMM_123_ARCACHE(M_AXIMM_123_ARCACHE),
        .M_AXIMM_123_ARPROT(M_AXIMM_123_ARPROT),
        .M_AXIMM_123_ARREGION(M_AXIMM_123_ARREGION),
        .M_AXIMM_123_ARQOS(M_AXIMM_123_ARQOS),
        .M_AXIMM_123_ARVALID(M_AXIMM_123_ARVALID),
        .M_AXIMM_123_ARREADY(M_AXIMM_123_ARREADY),
        .M_AXIMM_123_RDATA(M_AXIMM_123_RDATA),
        .M_AXIMM_123_RRESP(M_AXIMM_123_RRESP),
        .M_AXIMM_123_RLAST(M_AXIMM_123_RLAST),
        .M_AXIMM_123_RVALID(M_AXIMM_123_RVALID),
        .M_AXIMM_123_RREADY(M_AXIMM_123_RREADY),
        .AP_AXIMM_124_AWADDR(AP_AXIMM_124_AWADDR),
        .AP_AXIMM_124_AWLEN(AP_AXIMM_124_AWLEN),
        .AP_AXIMM_124_AWSIZE(AP_AXIMM_124_AWSIZE),
        .AP_AXIMM_124_AWBURST(AP_AXIMM_124_AWBURST),
        .AP_AXIMM_124_AWLOCK(AP_AXIMM_124_AWLOCK),
        .AP_AXIMM_124_AWCACHE(AP_AXIMM_124_AWCACHE),
        .AP_AXIMM_124_AWPROT(AP_AXIMM_124_AWPROT),
        .AP_AXIMM_124_AWREGION(AP_AXIMM_124_AWREGION),
        .AP_AXIMM_124_AWQOS(AP_AXIMM_124_AWQOS),
        .AP_AXIMM_124_AWVALID(AP_AXIMM_124_AWVALID),
        .AP_AXIMM_124_AWREADY(AP_AXIMM_124_AWREADY),
        .AP_AXIMM_124_WDATA(AP_AXIMM_124_WDATA),
        .AP_AXIMM_124_WSTRB(AP_AXIMM_124_WSTRB),
        .AP_AXIMM_124_WLAST(AP_AXIMM_124_WLAST),
        .AP_AXIMM_124_WVALID(AP_AXIMM_124_WVALID),
        .AP_AXIMM_124_WREADY(AP_AXIMM_124_WREADY),
        .AP_AXIMM_124_BRESP(AP_AXIMM_124_BRESP),
        .AP_AXIMM_124_BVALID(AP_AXIMM_124_BVALID),
        .AP_AXIMM_124_BREADY(AP_AXIMM_124_BREADY),
        .AP_AXIMM_124_ARADDR(AP_AXIMM_124_ARADDR),
        .AP_AXIMM_124_ARLEN(AP_AXIMM_124_ARLEN),
        .AP_AXIMM_124_ARSIZE(AP_AXIMM_124_ARSIZE),
        .AP_AXIMM_124_ARBURST(AP_AXIMM_124_ARBURST),
        .AP_AXIMM_124_ARLOCK(AP_AXIMM_124_ARLOCK),
        .AP_AXIMM_124_ARCACHE(AP_AXIMM_124_ARCACHE),
        .AP_AXIMM_124_ARPROT(AP_AXIMM_124_ARPROT),
        .AP_AXIMM_124_ARREGION(AP_AXIMM_124_ARREGION),
        .AP_AXIMM_124_ARQOS(AP_AXIMM_124_ARQOS),
        .AP_AXIMM_124_ARVALID(AP_AXIMM_124_ARVALID),
        .AP_AXIMM_124_ARREADY(AP_AXIMM_124_ARREADY),
        .AP_AXIMM_124_RDATA(AP_AXIMM_124_RDATA),
        .AP_AXIMM_124_RRESP(AP_AXIMM_124_RRESP),
        .AP_AXIMM_124_RLAST(AP_AXIMM_124_RLAST),
        .AP_AXIMM_124_RVALID(AP_AXIMM_124_RVALID),
        .AP_AXIMM_124_RREADY(AP_AXIMM_124_RREADY),
        .M_AXIMM_124_AWADDR(M_AXIMM_124_AWADDR),
        .M_AXIMM_124_AWLEN(M_AXIMM_124_AWLEN),
        .M_AXIMM_124_AWSIZE(M_AXIMM_124_AWSIZE),
        .M_AXIMM_124_AWBURST(M_AXIMM_124_AWBURST),
        .M_AXIMM_124_AWLOCK(M_AXIMM_124_AWLOCK),
        .M_AXIMM_124_AWCACHE(M_AXIMM_124_AWCACHE),
        .M_AXIMM_124_AWPROT(M_AXIMM_124_AWPROT),
        .M_AXIMM_124_AWREGION(M_AXIMM_124_AWREGION),
        .M_AXIMM_124_AWQOS(M_AXIMM_124_AWQOS),
        .M_AXIMM_124_AWVALID(M_AXIMM_124_AWVALID),
        .M_AXIMM_124_AWREADY(M_AXIMM_124_AWREADY),
        .M_AXIMM_124_WDATA(M_AXIMM_124_WDATA),
        .M_AXIMM_124_WSTRB(M_AXIMM_124_WSTRB),
        .M_AXIMM_124_WLAST(M_AXIMM_124_WLAST),
        .M_AXIMM_124_WVALID(M_AXIMM_124_WVALID),
        .M_AXIMM_124_WREADY(M_AXIMM_124_WREADY),
        .M_AXIMM_124_BRESP(M_AXIMM_124_BRESP),
        .M_AXIMM_124_BVALID(M_AXIMM_124_BVALID),
        .M_AXIMM_124_BREADY(M_AXIMM_124_BREADY),
        .M_AXIMM_124_ARADDR(M_AXIMM_124_ARADDR),
        .M_AXIMM_124_ARLEN(M_AXIMM_124_ARLEN),
        .M_AXIMM_124_ARSIZE(M_AXIMM_124_ARSIZE),
        .M_AXIMM_124_ARBURST(M_AXIMM_124_ARBURST),
        .M_AXIMM_124_ARLOCK(M_AXIMM_124_ARLOCK),
        .M_AXIMM_124_ARCACHE(M_AXIMM_124_ARCACHE),
        .M_AXIMM_124_ARPROT(M_AXIMM_124_ARPROT),
        .M_AXIMM_124_ARREGION(M_AXIMM_124_ARREGION),
        .M_AXIMM_124_ARQOS(M_AXIMM_124_ARQOS),
        .M_AXIMM_124_ARVALID(M_AXIMM_124_ARVALID),
        .M_AXIMM_124_ARREADY(M_AXIMM_124_ARREADY),
        .M_AXIMM_124_RDATA(M_AXIMM_124_RDATA),
        .M_AXIMM_124_RRESP(M_AXIMM_124_RRESP),
        .M_AXIMM_124_RLAST(M_AXIMM_124_RLAST),
        .M_AXIMM_124_RVALID(M_AXIMM_124_RVALID),
        .M_AXIMM_124_RREADY(M_AXIMM_124_RREADY),
        .AP_AXIMM_125_AWADDR(AP_AXIMM_125_AWADDR),
        .AP_AXIMM_125_AWLEN(AP_AXIMM_125_AWLEN),
        .AP_AXIMM_125_AWSIZE(AP_AXIMM_125_AWSIZE),
        .AP_AXIMM_125_AWBURST(AP_AXIMM_125_AWBURST),
        .AP_AXIMM_125_AWLOCK(AP_AXIMM_125_AWLOCK),
        .AP_AXIMM_125_AWCACHE(AP_AXIMM_125_AWCACHE),
        .AP_AXIMM_125_AWPROT(AP_AXIMM_125_AWPROT),
        .AP_AXIMM_125_AWREGION(AP_AXIMM_125_AWREGION),
        .AP_AXIMM_125_AWQOS(AP_AXIMM_125_AWQOS),
        .AP_AXIMM_125_AWVALID(AP_AXIMM_125_AWVALID),
        .AP_AXIMM_125_AWREADY(AP_AXIMM_125_AWREADY),
        .AP_AXIMM_125_WDATA(AP_AXIMM_125_WDATA),
        .AP_AXIMM_125_WSTRB(AP_AXIMM_125_WSTRB),
        .AP_AXIMM_125_WLAST(AP_AXIMM_125_WLAST),
        .AP_AXIMM_125_WVALID(AP_AXIMM_125_WVALID),
        .AP_AXIMM_125_WREADY(AP_AXIMM_125_WREADY),
        .AP_AXIMM_125_BRESP(AP_AXIMM_125_BRESP),
        .AP_AXIMM_125_BVALID(AP_AXIMM_125_BVALID),
        .AP_AXIMM_125_BREADY(AP_AXIMM_125_BREADY),
        .AP_AXIMM_125_ARADDR(AP_AXIMM_125_ARADDR),
        .AP_AXIMM_125_ARLEN(AP_AXIMM_125_ARLEN),
        .AP_AXIMM_125_ARSIZE(AP_AXIMM_125_ARSIZE),
        .AP_AXIMM_125_ARBURST(AP_AXIMM_125_ARBURST),
        .AP_AXIMM_125_ARLOCK(AP_AXIMM_125_ARLOCK),
        .AP_AXIMM_125_ARCACHE(AP_AXIMM_125_ARCACHE),
        .AP_AXIMM_125_ARPROT(AP_AXIMM_125_ARPROT),
        .AP_AXIMM_125_ARREGION(AP_AXIMM_125_ARREGION),
        .AP_AXIMM_125_ARQOS(AP_AXIMM_125_ARQOS),
        .AP_AXIMM_125_ARVALID(AP_AXIMM_125_ARVALID),
        .AP_AXIMM_125_ARREADY(AP_AXIMM_125_ARREADY),
        .AP_AXIMM_125_RDATA(AP_AXIMM_125_RDATA),
        .AP_AXIMM_125_RRESP(AP_AXIMM_125_RRESP),
        .AP_AXIMM_125_RLAST(AP_AXIMM_125_RLAST),
        .AP_AXIMM_125_RVALID(AP_AXIMM_125_RVALID),
        .AP_AXIMM_125_RREADY(AP_AXIMM_125_RREADY),
        .M_AXIMM_125_AWADDR(M_AXIMM_125_AWADDR),
        .M_AXIMM_125_AWLEN(M_AXIMM_125_AWLEN),
        .M_AXIMM_125_AWSIZE(M_AXIMM_125_AWSIZE),
        .M_AXIMM_125_AWBURST(M_AXIMM_125_AWBURST),
        .M_AXIMM_125_AWLOCK(M_AXIMM_125_AWLOCK),
        .M_AXIMM_125_AWCACHE(M_AXIMM_125_AWCACHE),
        .M_AXIMM_125_AWPROT(M_AXIMM_125_AWPROT),
        .M_AXIMM_125_AWREGION(M_AXIMM_125_AWREGION),
        .M_AXIMM_125_AWQOS(M_AXIMM_125_AWQOS),
        .M_AXIMM_125_AWVALID(M_AXIMM_125_AWVALID),
        .M_AXIMM_125_AWREADY(M_AXIMM_125_AWREADY),
        .M_AXIMM_125_WDATA(M_AXIMM_125_WDATA),
        .M_AXIMM_125_WSTRB(M_AXIMM_125_WSTRB),
        .M_AXIMM_125_WLAST(M_AXIMM_125_WLAST),
        .M_AXIMM_125_WVALID(M_AXIMM_125_WVALID),
        .M_AXIMM_125_WREADY(M_AXIMM_125_WREADY),
        .M_AXIMM_125_BRESP(M_AXIMM_125_BRESP),
        .M_AXIMM_125_BVALID(M_AXIMM_125_BVALID),
        .M_AXIMM_125_BREADY(M_AXIMM_125_BREADY),
        .M_AXIMM_125_ARADDR(M_AXIMM_125_ARADDR),
        .M_AXIMM_125_ARLEN(M_AXIMM_125_ARLEN),
        .M_AXIMM_125_ARSIZE(M_AXIMM_125_ARSIZE),
        .M_AXIMM_125_ARBURST(M_AXIMM_125_ARBURST),
        .M_AXIMM_125_ARLOCK(M_AXIMM_125_ARLOCK),
        .M_AXIMM_125_ARCACHE(M_AXIMM_125_ARCACHE),
        .M_AXIMM_125_ARPROT(M_AXIMM_125_ARPROT),
        .M_AXIMM_125_ARREGION(M_AXIMM_125_ARREGION),
        .M_AXIMM_125_ARQOS(M_AXIMM_125_ARQOS),
        .M_AXIMM_125_ARVALID(M_AXIMM_125_ARVALID),
        .M_AXIMM_125_ARREADY(M_AXIMM_125_ARREADY),
        .M_AXIMM_125_RDATA(M_AXIMM_125_RDATA),
        .M_AXIMM_125_RRESP(M_AXIMM_125_RRESP),
        .M_AXIMM_125_RLAST(M_AXIMM_125_RLAST),
        .M_AXIMM_125_RVALID(M_AXIMM_125_RVALID),
        .M_AXIMM_125_RREADY(M_AXIMM_125_RREADY),
        .AP_AXIMM_126_AWADDR(AP_AXIMM_126_AWADDR),
        .AP_AXIMM_126_AWLEN(AP_AXIMM_126_AWLEN),
        .AP_AXIMM_126_AWSIZE(AP_AXIMM_126_AWSIZE),
        .AP_AXIMM_126_AWBURST(AP_AXIMM_126_AWBURST),
        .AP_AXIMM_126_AWLOCK(AP_AXIMM_126_AWLOCK),
        .AP_AXIMM_126_AWCACHE(AP_AXIMM_126_AWCACHE),
        .AP_AXIMM_126_AWPROT(AP_AXIMM_126_AWPROT),
        .AP_AXIMM_126_AWREGION(AP_AXIMM_126_AWREGION),
        .AP_AXIMM_126_AWQOS(AP_AXIMM_126_AWQOS),
        .AP_AXIMM_126_AWVALID(AP_AXIMM_126_AWVALID),
        .AP_AXIMM_126_AWREADY(AP_AXIMM_126_AWREADY),
        .AP_AXIMM_126_WDATA(AP_AXIMM_126_WDATA),
        .AP_AXIMM_126_WSTRB(AP_AXIMM_126_WSTRB),
        .AP_AXIMM_126_WLAST(AP_AXIMM_126_WLAST),
        .AP_AXIMM_126_WVALID(AP_AXIMM_126_WVALID),
        .AP_AXIMM_126_WREADY(AP_AXIMM_126_WREADY),
        .AP_AXIMM_126_BRESP(AP_AXIMM_126_BRESP),
        .AP_AXIMM_126_BVALID(AP_AXIMM_126_BVALID),
        .AP_AXIMM_126_BREADY(AP_AXIMM_126_BREADY),
        .AP_AXIMM_126_ARADDR(AP_AXIMM_126_ARADDR),
        .AP_AXIMM_126_ARLEN(AP_AXIMM_126_ARLEN),
        .AP_AXIMM_126_ARSIZE(AP_AXIMM_126_ARSIZE),
        .AP_AXIMM_126_ARBURST(AP_AXIMM_126_ARBURST),
        .AP_AXIMM_126_ARLOCK(AP_AXIMM_126_ARLOCK),
        .AP_AXIMM_126_ARCACHE(AP_AXIMM_126_ARCACHE),
        .AP_AXIMM_126_ARPROT(AP_AXIMM_126_ARPROT),
        .AP_AXIMM_126_ARREGION(AP_AXIMM_126_ARREGION),
        .AP_AXIMM_126_ARQOS(AP_AXIMM_126_ARQOS),
        .AP_AXIMM_126_ARVALID(AP_AXIMM_126_ARVALID),
        .AP_AXIMM_126_ARREADY(AP_AXIMM_126_ARREADY),
        .AP_AXIMM_126_RDATA(AP_AXIMM_126_RDATA),
        .AP_AXIMM_126_RRESP(AP_AXIMM_126_RRESP),
        .AP_AXIMM_126_RLAST(AP_AXIMM_126_RLAST),
        .AP_AXIMM_126_RVALID(AP_AXIMM_126_RVALID),
        .AP_AXIMM_126_RREADY(AP_AXIMM_126_RREADY),
        .M_AXIMM_126_AWADDR(M_AXIMM_126_AWADDR),
        .M_AXIMM_126_AWLEN(M_AXIMM_126_AWLEN),
        .M_AXIMM_126_AWSIZE(M_AXIMM_126_AWSIZE),
        .M_AXIMM_126_AWBURST(M_AXIMM_126_AWBURST),
        .M_AXIMM_126_AWLOCK(M_AXIMM_126_AWLOCK),
        .M_AXIMM_126_AWCACHE(M_AXIMM_126_AWCACHE),
        .M_AXIMM_126_AWPROT(M_AXIMM_126_AWPROT),
        .M_AXIMM_126_AWREGION(M_AXIMM_126_AWREGION),
        .M_AXIMM_126_AWQOS(M_AXIMM_126_AWQOS),
        .M_AXIMM_126_AWVALID(M_AXIMM_126_AWVALID),
        .M_AXIMM_126_AWREADY(M_AXIMM_126_AWREADY),
        .M_AXIMM_126_WDATA(M_AXIMM_126_WDATA),
        .M_AXIMM_126_WSTRB(M_AXIMM_126_WSTRB),
        .M_AXIMM_126_WLAST(M_AXIMM_126_WLAST),
        .M_AXIMM_126_WVALID(M_AXIMM_126_WVALID),
        .M_AXIMM_126_WREADY(M_AXIMM_126_WREADY),
        .M_AXIMM_126_BRESP(M_AXIMM_126_BRESP),
        .M_AXIMM_126_BVALID(M_AXIMM_126_BVALID),
        .M_AXIMM_126_BREADY(M_AXIMM_126_BREADY),
        .M_AXIMM_126_ARADDR(M_AXIMM_126_ARADDR),
        .M_AXIMM_126_ARLEN(M_AXIMM_126_ARLEN),
        .M_AXIMM_126_ARSIZE(M_AXIMM_126_ARSIZE),
        .M_AXIMM_126_ARBURST(M_AXIMM_126_ARBURST),
        .M_AXIMM_126_ARLOCK(M_AXIMM_126_ARLOCK),
        .M_AXIMM_126_ARCACHE(M_AXIMM_126_ARCACHE),
        .M_AXIMM_126_ARPROT(M_AXIMM_126_ARPROT),
        .M_AXIMM_126_ARREGION(M_AXIMM_126_ARREGION),
        .M_AXIMM_126_ARQOS(M_AXIMM_126_ARQOS),
        .M_AXIMM_126_ARVALID(M_AXIMM_126_ARVALID),
        .M_AXIMM_126_ARREADY(M_AXIMM_126_ARREADY),
        .M_AXIMM_126_RDATA(M_AXIMM_126_RDATA),
        .M_AXIMM_126_RRESP(M_AXIMM_126_RRESP),
        .M_AXIMM_126_RLAST(M_AXIMM_126_RLAST),
        .M_AXIMM_126_RVALID(M_AXIMM_126_RVALID),
        .M_AXIMM_126_RREADY(M_AXIMM_126_RREADY),
        .AP_AXIMM_127_AWADDR(AP_AXIMM_127_AWADDR),
        .AP_AXIMM_127_AWLEN(AP_AXIMM_127_AWLEN),
        .AP_AXIMM_127_AWSIZE(AP_AXIMM_127_AWSIZE),
        .AP_AXIMM_127_AWBURST(AP_AXIMM_127_AWBURST),
        .AP_AXIMM_127_AWLOCK(AP_AXIMM_127_AWLOCK),
        .AP_AXIMM_127_AWCACHE(AP_AXIMM_127_AWCACHE),
        .AP_AXIMM_127_AWPROT(AP_AXIMM_127_AWPROT),
        .AP_AXIMM_127_AWREGION(AP_AXIMM_127_AWREGION),
        .AP_AXIMM_127_AWQOS(AP_AXIMM_127_AWQOS),
        .AP_AXIMM_127_AWVALID(AP_AXIMM_127_AWVALID),
        .AP_AXIMM_127_AWREADY(AP_AXIMM_127_AWREADY),
        .AP_AXIMM_127_WDATA(AP_AXIMM_127_WDATA),
        .AP_AXIMM_127_WSTRB(AP_AXIMM_127_WSTRB),
        .AP_AXIMM_127_WLAST(AP_AXIMM_127_WLAST),
        .AP_AXIMM_127_WVALID(AP_AXIMM_127_WVALID),
        .AP_AXIMM_127_WREADY(AP_AXIMM_127_WREADY),
        .AP_AXIMM_127_BRESP(AP_AXIMM_127_BRESP),
        .AP_AXIMM_127_BVALID(AP_AXIMM_127_BVALID),
        .AP_AXIMM_127_BREADY(AP_AXIMM_127_BREADY),
        .AP_AXIMM_127_ARADDR(AP_AXIMM_127_ARADDR),
        .AP_AXIMM_127_ARLEN(AP_AXIMM_127_ARLEN),
        .AP_AXIMM_127_ARSIZE(AP_AXIMM_127_ARSIZE),
        .AP_AXIMM_127_ARBURST(AP_AXIMM_127_ARBURST),
        .AP_AXIMM_127_ARLOCK(AP_AXIMM_127_ARLOCK),
        .AP_AXIMM_127_ARCACHE(AP_AXIMM_127_ARCACHE),
        .AP_AXIMM_127_ARPROT(AP_AXIMM_127_ARPROT),
        .AP_AXIMM_127_ARREGION(AP_AXIMM_127_ARREGION),
        .AP_AXIMM_127_ARQOS(AP_AXIMM_127_ARQOS),
        .AP_AXIMM_127_ARVALID(AP_AXIMM_127_ARVALID),
        .AP_AXIMM_127_ARREADY(AP_AXIMM_127_ARREADY),
        .AP_AXIMM_127_RDATA(AP_AXIMM_127_RDATA),
        .AP_AXIMM_127_RRESP(AP_AXIMM_127_RRESP),
        .AP_AXIMM_127_RLAST(AP_AXIMM_127_RLAST),
        .AP_AXIMM_127_RVALID(AP_AXIMM_127_RVALID),
        .AP_AXIMM_127_RREADY(AP_AXIMM_127_RREADY),
        .M_AXIMM_127_AWADDR(M_AXIMM_127_AWADDR),
        .M_AXIMM_127_AWLEN(M_AXIMM_127_AWLEN),
        .M_AXIMM_127_AWSIZE(M_AXIMM_127_AWSIZE),
        .M_AXIMM_127_AWBURST(M_AXIMM_127_AWBURST),
        .M_AXIMM_127_AWLOCK(M_AXIMM_127_AWLOCK),
        .M_AXIMM_127_AWCACHE(M_AXIMM_127_AWCACHE),
        .M_AXIMM_127_AWPROT(M_AXIMM_127_AWPROT),
        .M_AXIMM_127_AWREGION(M_AXIMM_127_AWREGION),
        .M_AXIMM_127_AWQOS(M_AXIMM_127_AWQOS),
        .M_AXIMM_127_AWVALID(M_AXIMM_127_AWVALID),
        .M_AXIMM_127_AWREADY(M_AXIMM_127_AWREADY),
        .M_AXIMM_127_WDATA(M_AXIMM_127_WDATA),
        .M_AXIMM_127_WSTRB(M_AXIMM_127_WSTRB),
        .M_AXIMM_127_WLAST(M_AXIMM_127_WLAST),
        .M_AXIMM_127_WVALID(M_AXIMM_127_WVALID),
        .M_AXIMM_127_WREADY(M_AXIMM_127_WREADY),
        .M_AXIMM_127_BRESP(M_AXIMM_127_BRESP),
        .M_AXIMM_127_BVALID(M_AXIMM_127_BVALID),
        .M_AXIMM_127_BREADY(M_AXIMM_127_BREADY),
        .M_AXIMM_127_ARADDR(M_AXIMM_127_ARADDR),
        .M_AXIMM_127_ARLEN(M_AXIMM_127_ARLEN),
        .M_AXIMM_127_ARSIZE(M_AXIMM_127_ARSIZE),
        .M_AXIMM_127_ARBURST(M_AXIMM_127_ARBURST),
        .M_AXIMM_127_ARLOCK(M_AXIMM_127_ARLOCK),
        .M_AXIMM_127_ARCACHE(M_AXIMM_127_ARCACHE),
        .M_AXIMM_127_ARPROT(M_AXIMM_127_ARPROT),
        .M_AXIMM_127_ARREGION(M_AXIMM_127_ARREGION),
        .M_AXIMM_127_ARQOS(M_AXIMM_127_ARQOS),
        .M_AXIMM_127_ARVALID(M_AXIMM_127_ARVALID),
        .M_AXIMM_127_ARREADY(M_AXIMM_127_ARREADY),
        .M_AXIMM_127_RDATA(M_AXIMM_127_RDATA),
        .M_AXIMM_127_RRESP(M_AXIMM_127_RRESP),
        .M_AXIMM_127_RLAST(M_AXIMM_127_RLAST),
        .M_AXIMM_127_RVALID(M_AXIMM_127_RVALID),
        .M_AXIMM_127_RREADY(M_AXIMM_127_RREADY)
    );
    
    in_bram_args #(
        .C_NUM_INPUT_BRAMs(C_NUM_INPUT_BRAMs),
        .S_AXIS_BRAM_0_PORTS(S_AXIS_BRAM_0_PORTS),
        .S_AXIS_BRAM_1_PORTS(S_AXIS_BRAM_1_PORTS),
        .S_AXIS_BRAM_2_PORTS(S_AXIS_BRAM_2_PORTS),
        .S_AXIS_BRAM_3_PORTS(S_AXIS_BRAM_3_PORTS),
        .S_AXIS_BRAM_4_PORTS(S_AXIS_BRAM_4_PORTS),
        .S_AXIS_BRAM_5_PORTS(S_AXIS_BRAM_5_PORTS),
        .S_AXIS_BRAM_6_PORTS(S_AXIS_BRAM_6_PORTS),
        .S_AXIS_BRAM_7_PORTS(S_AXIS_BRAM_7_PORTS),
        .S_AXIS_BRAM_8_PORTS(S_AXIS_BRAM_8_PORTS),
        .S_AXIS_BRAM_9_PORTS(S_AXIS_BRAM_9_PORTS),
        .S_AXIS_BRAM_10_PORTS(S_AXIS_BRAM_10_PORTS),
        .S_AXIS_BRAM_11_PORTS(S_AXIS_BRAM_11_PORTS),
        .S_AXIS_BRAM_12_PORTS(S_AXIS_BRAM_12_PORTS),
        .S_AXIS_BRAM_13_PORTS(S_AXIS_BRAM_13_PORTS),
        .S_AXIS_BRAM_14_PORTS(S_AXIS_BRAM_14_PORTS),
        .S_AXIS_BRAM_15_PORTS(S_AXIS_BRAM_15_PORTS),
        .S_AXIS_BRAM_16_PORTS(S_AXIS_BRAM_16_PORTS),
        .S_AXIS_BRAM_17_PORTS(S_AXIS_BRAM_17_PORTS),
        .S_AXIS_BRAM_18_PORTS(S_AXIS_BRAM_18_PORTS),
        .S_AXIS_BRAM_19_PORTS(S_AXIS_BRAM_19_PORTS),
        .S_AXIS_BRAM_20_PORTS(S_AXIS_BRAM_20_PORTS),
        .S_AXIS_BRAM_21_PORTS(S_AXIS_BRAM_21_PORTS),
        .S_AXIS_BRAM_22_PORTS(S_AXIS_BRAM_22_PORTS),
        .S_AXIS_BRAM_23_PORTS(S_AXIS_BRAM_23_PORTS),
        .S_AXIS_BRAM_24_PORTS(S_AXIS_BRAM_24_PORTS),
        .S_AXIS_BRAM_25_PORTS(S_AXIS_BRAM_25_PORTS),
        .S_AXIS_BRAM_26_PORTS(S_AXIS_BRAM_26_PORTS),
        .S_AXIS_BRAM_27_PORTS(S_AXIS_BRAM_27_PORTS),
        .S_AXIS_BRAM_28_PORTS(S_AXIS_BRAM_28_PORTS),
        .S_AXIS_BRAM_29_PORTS(S_AXIS_BRAM_29_PORTS),
        .S_AXIS_BRAM_30_PORTS(S_AXIS_BRAM_30_PORTS),
        .S_AXIS_BRAM_31_PORTS(S_AXIS_BRAM_31_PORTS),
        .S_AXIS_BRAM_32_PORTS(S_AXIS_BRAM_32_PORTS),
        .S_AXIS_BRAM_33_PORTS(S_AXIS_BRAM_33_PORTS),
        .S_AXIS_BRAM_34_PORTS(S_AXIS_BRAM_34_PORTS),
        .S_AXIS_BRAM_35_PORTS(S_AXIS_BRAM_35_PORTS),
        .S_AXIS_BRAM_36_PORTS(S_AXIS_BRAM_36_PORTS),
        .S_AXIS_BRAM_37_PORTS(S_AXIS_BRAM_37_PORTS),
        .S_AXIS_BRAM_38_PORTS(S_AXIS_BRAM_38_PORTS),
        .S_AXIS_BRAM_39_PORTS(S_AXIS_BRAM_39_PORTS),
        .S_AXIS_BRAM_40_PORTS(S_AXIS_BRAM_40_PORTS),
        .S_AXIS_BRAM_41_PORTS(S_AXIS_BRAM_41_PORTS),
        .S_AXIS_BRAM_42_PORTS(S_AXIS_BRAM_42_PORTS),
        .S_AXIS_BRAM_43_PORTS(S_AXIS_BRAM_43_PORTS),
        .S_AXIS_BRAM_44_PORTS(S_AXIS_BRAM_44_PORTS),
        .S_AXIS_BRAM_45_PORTS(S_AXIS_BRAM_45_PORTS),
        .S_AXIS_BRAM_46_PORTS(S_AXIS_BRAM_46_PORTS),
        .S_AXIS_BRAM_47_PORTS(S_AXIS_BRAM_47_PORTS),
        .S_AXIS_BRAM_48_PORTS(S_AXIS_BRAM_48_PORTS),
        .S_AXIS_BRAM_49_PORTS(S_AXIS_BRAM_49_PORTS),
        .S_AXIS_BRAM_50_PORTS(S_AXIS_BRAM_50_PORTS),
        .S_AXIS_BRAM_51_PORTS(S_AXIS_BRAM_51_PORTS),
        .S_AXIS_BRAM_52_PORTS(S_AXIS_BRAM_52_PORTS),
        .S_AXIS_BRAM_53_PORTS(S_AXIS_BRAM_53_PORTS),
        .S_AXIS_BRAM_54_PORTS(S_AXIS_BRAM_54_PORTS),
        .S_AXIS_BRAM_55_PORTS(S_AXIS_BRAM_55_PORTS),
        .S_AXIS_BRAM_56_PORTS(S_AXIS_BRAM_56_PORTS),
        .S_AXIS_BRAM_57_PORTS(S_AXIS_BRAM_57_PORTS),
        .S_AXIS_BRAM_58_PORTS(S_AXIS_BRAM_58_PORTS),
        .S_AXIS_BRAM_59_PORTS(S_AXIS_BRAM_59_PORTS),
        .S_AXIS_BRAM_60_PORTS(S_AXIS_BRAM_60_PORTS),
        .S_AXIS_BRAM_61_PORTS(S_AXIS_BRAM_61_PORTS),
        .S_AXIS_BRAM_62_PORTS(S_AXIS_BRAM_62_PORTS),
        .S_AXIS_BRAM_63_PORTS(S_AXIS_BRAM_63_PORTS),
        .S_AXIS_BRAM_64_PORTS(S_AXIS_BRAM_64_PORTS),
        .S_AXIS_BRAM_65_PORTS(S_AXIS_BRAM_65_PORTS),
        .S_AXIS_BRAM_66_PORTS(S_AXIS_BRAM_66_PORTS),
        .S_AXIS_BRAM_67_PORTS(S_AXIS_BRAM_67_PORTS),
        .S_AXIS_BRAM_68_PORTS(S_AXIS_BRAM_68_PORTS),
        .S_AXIS_BRAM_69_PORTS(S_AXIS_BRAM_69_PORTS),
        .S_AXIS_BRAM_70_PORTS(S_AXIS_BRAM_70_PORTS),
        .S_AXIS_BRAM_71_PORTS(S_AXIS_BRAM_71_PORTS),
        .S_AXIS_BRAM_72_PORTS(S_AXIS_BRAM_72_PORTS),
        .S_AXIS_BRAM_73_PORTS(S_AXIS_BRAM_73_PORTS),
        .S_AXIS_BRAM_74_PORTS(S_AXIS_BRAM_74_PORTS),
        .S_AXIS_BRAM_75_PORTS(S_AXIS_BRAM_75_PORTS),
        .S_AXIS_BRAM_76_PORTS(S_AXIS_BRAM_76_PORTS),
        .S_AXIS_BRAM_77_PORTS(S_AXIS_BRAM_77_PORTS),
        .S_AXIS_BRAM_78_PORTS(S_AXIS_BRAM_78_PORTS),
        .S_AXIS_BRAM_79_PORTS(S_AXIS_BRAM_79_PORTS),
        .S_AXIS_BRAM_80_PORTS(S_AXIS_BRAM_80_PORTS),
        .S_AXIS_BRAM_81_PORTS(S_AXIS_BRAM_81_PORTS),
        .S_AXIS_BRAM_82_PORTS(S_AXIS_BRAM_82_PORTS),
        .S_AXIS_BRAM_83_PORTS(S_AXIS_BRAM_83_PORTS),
        .S_AXIS_BRAM_84_PORTS(S_AXIS_BRAM_84_PORTS),
        .S_AXIS_BRAM_85_PORTS(S_AXIS_BRAM_85_PORTS),
        .S_AXIS_BRAM_86_PORTS(S_AXIS_BRAM_86_PORTS),
        .S_AXIS_BRAM_87_PORTS(S_AXIS_BRAM_87_PORTS),
        .S_AXIS_BRAM_88_PORTS(S_AXIS_BRAM_88_PORTS),
        .S_AXIS_BRAM_89_PORTS(S_AXIS_BRAM_89_PORTS),
        .S_AXIS_BRAM_90_PORTS(S_AXIS_BRAM_90_PORTS),
        .S_AXIS_BRAM_91_PORTS(S_AXIS_BRAM_91_PORTS),
        .S_AXIS_BRAM_92_PORTS(S_AXIS_BRAM_92_PORTS),
        .S_AXIS_BRAM_93_PORTS(S_AXIS_BRAM_93_PORTS),
        .S_AXIS_BRAM_94_PORTS(S_AXIS_BRAM_94_PORTS),
        .S_AXIS_BRAM_95_PORTS(S_AXIS_BRAM_95_PORTS),
        .S_AXIS_BRAM_96_PORTS(S_AXIS_BRAM_96_PORTS),
        .S_AXIS_BRAM_97_PORTS(S_AXIS_BRAM_97_PORTS),
        .S_AXIS_BRAM_98_PORTS(S_AXIS_BRAM_98_PORTS),
        .S_AXIS_BRAM_99_PORTS(S_AXIS_BRAM_99_PORTS),
        .S_AXIS_BRAM_100_PORTS(S_AXIS_BRAM_100_PORTS),
        .S_AXIS_BRAM_101_PORTS(S_AXIS_BRAM_101_PORTS),
        .S_AXIS_BRAM_102_PORTS(S_AXIS_BRAM_102_PORTS),
        .S_AXIS_BRAM_103_PORTS(S_AXIS_BRAM_103_PORTS),
        .S_AXIS_BRAM_104_PORTS(S_AXIS_BRAM_104_PORTS),
        .S_AXIS_BRAM_105_PORTS(S_AXIS_BRAM_105_PORTS),
        .S_AXIS_BRAM_106_PORTS(S_AXIS_BRAM_106_PORTS),
        .S_AXIS_BRAM_107_PORTS(S_AXIS_BRAM_107_PORTS),
        .S_AXIS_BRAM_108_PORTS(S_AXIS_BRAM_108_PORTS),
        .S_AXIS_BRAM_109_PORTS(S_AXIS_BRAM_109_PORTS),
        .S_AXIS_BRAM_110_PORTS(S_AXIS_BRAM_110_PORTS),
        .S_AXIS_BRAM_111_PORTS(S_AXIS_BRAM_111_PORTS),
        .S_AXIS_BRAM_112_PORTS(S_AXIS_BRAM_112_PORTS),
        .S_AXIS_BRAM_113_PORTS(S_AXIS_BRAM_113_PORTS),
        .S_AXIS_BRAM_114_PORTS(S_AXIS_BRAM_114_PORTS),
        .S_AXIS_BRAM_115_PORTS(S_AXIS_BRAM_115_PORTS),
        .S_AXIS_BRAM_116_PORTS(S_AXIS_BRAM_116_PORTS),
        .S_AXIS_BRAM_117_PORTS(S_AXIS_BRAM_117_PORTS),
        .S_AXIS_BRAM_118_PORTS(S_AXIS_BRAM_118_PORTS),
        .S_AXIS_BRAM_119_PORTS(S_AXIS_BRAM_119_PORTS),
        .S_AXIS_BRAM_120_PORTS(S_AXIS_BRAM_120_PORTS),
        .S_AXIS_BRAM_121_PORTS(S_AXIS_BRAM_121_PORTS),
        .S_AXIS_BRAM_122_PORTS(S_AXIS_BRAM_122_PORTS),
        .S_AXIS_BRAM_123_PORTS(S_AXIS_BRAM_123_PORTS),
        .S_AXIS_BRAM_124_PORTS(S_AXIS_BRAM_124_PORTS),
        .S_AXIS_BRAM_125_PORTS(S_AXIS_BRAM_125_PORTS),
        .S_AXIS_BRAM_126_PORTS(S_AXIS_BRAM_126_PORTS),
        .S_AXIS_BRAM_127_PORTS(S_AXIS_BRAM_127_PORTS),
        .S_AXIS_BRAM_0_WIDTH(S_AXIS_BRAM_0_WIDTH),
        .S_AXIS_BRAM_1_WIDTH(S_AXIS_BRAM_1_WIDTH),
        .S_AXIS_BRAM_2_WIDTH(S_AXIS_BRAM_2_WIDTH),
        .S_AXIS_BRAM_3_WIDTH(S_AXIS_BRAM_3_WIDTH),
        .S_AXIS_BRAM_4_WIDTH(S_AXIS_BRAM_4_WIDTH),
        .S_AXIS_BRAM_5_WIDTH(S_AXIS_BRAM_5_WIDTH),
        .S_AXIS_BRAM_6_WIDTH(S_AXIS_BRAM_6_WIDTH),
        .S_AXIS_BRAM_7_WIDTH(S_AXIS_BRAM_7_WIDTH),
        .S_AXIS_BRAM_8_WIDTH(S_AXIS_BRAM_8_WIDTH),
        .S_AXIS_BRAM_9_WIDTH(S_AXIS_BRAM_9_WIDTH),
        .S_AXIS_BRAM_10_WIDTH(S_AXIS_BRAM_10_WIDTH),
        .S_AXIS_BRAM_11_WIDTH(S_AXIS_BRAM_11_WIDTH),
        .S_AXIS_BRAM_12_WIDTH(S_AXIS_BRAM_12_WIDTH),
        .S_AXIS_BRAM_13_WIDTH(S_AXIS_BRAM_13_WIDTH),
        .S_AXIS_BRAM_14_WIDTH(S_AXIS_BRAM_14_WIDTH),
        .S_AXIS_BRAM_15_WIDTH(S_AXIS_BRAM_15_WIDTH),
        .S_AXIS_BRAM_16_WIDTH(S_AXIS_BRAM_16_WIDTH),
        .S_AXIS_BRAM_17_WIDTH(S_AXIS_BRAM_17_WIDTH),
        .S_AXIS_BRAM_18_WIDTH(S_AXIS_BRAM_18_WIDTH),
        .S_AXIS_BRAM_19_WIDTH(S_AXIS_BRAM_19_WIDTH),
        .S_AXIS_BRAM_20_WIDTH(S_AXIS_BRAM_20_WIDTH),
        .S_AXIS_BRAM_21_WIDTH(S_AXIS_BRAM_21_WIDTH),
        .S_AXIS_BRAM_22_WIDTH(S_AXIS_BRAM_22_WIDTH),
        .S_AXIS_BRAM_23_WIDTH(S_AXIS_BRAM_23_WIDTH),
        .S_AXIS_BRAM_24_WIDTH(S_AXIS_BRAM_24_WIDTH),
        .S_AXIS_BRAM_25_WIDTH(S_AXIS_BRAM_25_WIDTH),
        .S_AXIS_BRAM_26_WIDTH(S_AXIS_BRAM_26_WIDTH),
        .S_AXIS_BRAM_27_WIDTH(S_AXIS_BRAM_27_WIDTH),
        .S_AXIS_BRAM_28_WIDTH(S_AXIS_BRAM_28_WIDTH),
        .S_AXIS_BRAM_29_WIDTH(S_AXIS_BRAM_29_WIDTH),
        .S_AXIS_BRAM_30_WIDTH(S_AXIS_BRAM_30_WIDTH),
        .S_AXIS_BRAM_31_WIDTH(S_AXIS_BRAM_31_WIDTH),
        .S_AXIS_BRAM_32_WIDTH(S_AXIS_BRAM_32_WIDTH),
        .S_AXIS_BRAM_33_WIDTH(S_AXIS_BRAM_33_WIDTH),
        .S_AXIS_BRAM_34_WIDTH(S_AXIS_BRAM_34_WIDTH),
        .S_AXIS_BRAM_35_WIDTH(S_AXIS_BRAM_35_WIDTH),
        .S_AXIS_BRAM_36_WIDTH(S_AXIS_BRAM_36_WIDTH),
        .S_AXIS_BRAM_37_WIDTH(S_AXIS_BRAM_37_WIDTH),
        .S_AXIS_BRAM_38_WIDTH(S_AXIS_BRAM_38_WIDTH),
        .S_AXIS_BRAM_39_WIDTH(S_AXIS_BRAM_39_WIDTH),
        .S_AXIS_BRAM_40_WIDTH(S_AXIS_BRAM_40_WIDTH),
        .S_AXIS_BRAM_41_WIDTH(S_AXIS_BRAM_41_WIDTH),
        .S_AXIS_BRAM_42_WIDTH(S_AXIS_BRAM_42_WIDTH),
        .S_AXIS_BRAM_43_WIDTH(S_AXIS_BRAM_43_WIDTH),
        .S_AXIS_BRAM_44_WIDTH(S_AXIS_BRAM_44_WIDTH),
        .S_AXIS_BRAM_45_WIDTH(S_AXIS_BRAM_45_WIDTH),
        .S_AXIS_BRAM_46_WIDTH(S_AXIS_BRAM_46_WIDTH),
        .S_AXIS_BRAM_47_WIDTH(S_AXIS_BRAM_47_WIDTH),
        .S_AXIS_BRAM_48_WIDTH(S_AXIS_BRAM_48_WIDTH),
        .S_AXIS_BRAM_49_WIDTH(S_AXIS_BRAM_49_WIDTH),
        .S_AXIS_BRAM_50_WIDTH(S_AXIS_BRAM_50_WIDTH),
        .S_AXIS_BRAM_51_WIDTH(S_AXIS_BRAM_51_WIDTH),
        .S_AXIS_BRAM_52_WIDTH(S_AXIS_BRAM_52_WIDTH),
        .S_AXIS_BRAM_53_WIDTH(S_AXIS_BRAM_53_WIDTH),
        .S_AXIS_BRAM_54_WIDTH(S_AXIS_BRAM_54_WIDTH),
        .S_AXIS_BRAM_55_WIDTH(S_AXIS_BRAM_55_WIDTH),
        .S_AXIS_BRAM_56_WIDTH(S_AXIS_BRAM_56_WIDTH),
        .S_AXIS_BRAM_57_WIDTH(S_AXIS_BRAM_57_WIDTH),
        .S_AXIS_BRAM_58_WIDTH(S_AXIS_BRAM_58_WIDTH),
        .S_AXIS_BRAM_59_WIDTH(S_AXIS_BRAM_59_WIDTH),
        .S_AXIS_BRAM_60_WIDTH(S_AXIS_BRAM_60_WIDTH),
        .S_AXIS_BRAM_61_WIDTH(S_AXIS_BRAM_61_WIDTH),
        .S_AXIS_BRAM_62_WIDTH(S_AXIS_BRAM_62_WIDTH),
        .S_AXIS_BRAM_63_WIDTH(S_AXIS_BRAM_63_WIDTH),
        .S_AXIS_BRAM_64_WIDTH(S_AXIS_BRAM_64_WIDTH),
        .S_AXIS_BRAM_65_WIDTH(S_AXIS_BRAM_65_WIDTH),
        .S_AXIS_BRAM_66_WIDTH(S_AXIS_BRAM_66_WIDTH),
        .S_AXIS_BRAM_67_WIDTH(S_AXIS_BRAM_67_WIDTH),
        .S_AXIS_BRAM_68_WIDTH(S_AXIS_BRAM_68_WIDTH),
        .S_AXIS_BRAM_69_WIDTH(S_AXIS_BRAM_69_WIDTH),
        .S_AXIS_BRAM_70_WIDTH(S_AXIS_BRAM_70_WIDTH),
        .S_AXIS_BRAM_71_WIDTH(S_AXIS_BRAM_71_WIDTH),
        .S_AXIS_BRAM_72_WIDTH(S_AXIS_BRAM_72_WIDTH),
        .S_AXIS_BRAM_73_WIDTH(S_AXIS_BRAM_73_WIDTH),
        .S_AXIS_BRAM_74_WIDTH(S_AXIS_BRAM_74_WIDTH),
        .S_AXIS_BRAM_75_WIDTH(S_AXIS_BRAM_75_WIDTH),
        .S_AXIS_BRAM_76_WIDTH(S_AXIS_BRAM_76_WIDTH),
        .S_AXIS_BRAM_77_WIDTH(S_AXIS_BRAM_77_WIDTH),
        .S_AXIS_BRAM_78_WIDTH(S_AXIS_BRAM_78_WIDTH),
        .S_AXIS_BRAM_79_WIDTH(S_AXIS_BRAM_79_WIDTH),
        .S_AXIS_BRAM_80_WIDTH(S_AXIS_BRAM_80_WIDTH),
        .S_AXIS_BRAM_81_WIDTH(S_AXIS_BRAM_81_WIDTH),
        .S_AXIS_BRAM_82_WIDTH(S_AXIS_BRAM_82_WIDTH),
        .S_AXIS_BRAM_83_WIDTH(S_AXIS_BRAM_83_WIDTH),
        .S_AXIS_BRAM_84_WIDTH(S_AXIS_BRAM_84_WIDTH),
        .S_AXIS_BRAM_85_WIDTH(S_AXIS_BRAM_85_WIDTH),
        .S_AXIS_BRAM_86_WIDTH(S_AXIS_BRAM_86_WIDTH),
        .S_AXIS_BRAM_87_WIDTH(S_AXIS_BRAM_87_WIDTH),
        .S_AXIS_BRAM_88_WIDTH(S_AXIS_BRAM_88_WIDTH),
        .S_AXIS_BRAM_89_WIDTH(S_AXIS_BRAM_89_WIDTH),
        .S_AXIS_BRAM_90_WIDTH(S_AXIS_BRAM_90_WIDTH),
        .S_AXIS_BRAM_91_WIDTH(S_AXIS_BRAM_91_WIDTH),
        .S_AXIS_BRAM_92_WIDTH(S_AXIS_BRAM_92_WIDTH),
        .S_AXIS_BRAM_93_WIDTH(S_AXIS_BRAM_93_WIDTH),
        .S_AXIS_BRAM_94_WIDTH(S_AXIS_BRAM_94_WIDTH),
        .S_AXIS_BRAM_95_WIDTH(S_AXIS_BRAM_95_WIDTH),
        .S_AXIS_BRAM_96_WIDTH(S_AXIS_BRAM_96_WIDTH),
        .S_AXIS_BRAM_97_WIDTH(S_AXIS_BRAM_97_WIDTH),
        .S_AXIS_BRAM_98_WIDTH(S_AXIS_BRAM_98_WIDTH),
        .S_AXIS_BRAM_99_WIDTH(S_AXIS_BRAM_99_WIDTH),
        .S_AXIS_BRAM_100_WIDTH(S_AXIS_BRAM_100_WIDTH),
        .S_AXIS_BRAM_101_WIDTH(S_AXIS_BRAM_101_WIDTH),
        .S_AXIS_BRAM_102_WIDTH(S_AXIS_BRAM_102_WIDTH),
        .S_AXIS_BRAM_103_WIDTH(S_AXIS_BRAM_103_WIDTH),
        .S_AXIS_BRAM_104_WIDTH(S_AXIS_BRAM_104_WIDTH),
        .S_AXIS_BRAM_105_WIDTH(S_AXIS_BRAM_105_WIDTH),
        .S_AXIS_BRAM_106_WIDTH(S_AXIS_BRAM_106_WIDTH),
        .S_AXIS_BRAM_107_WIDTH(S_AXIS_BRAM_107_WIDTH),
        .S_AXIS_BRAM_108_WIDTH(S_AXIS_BRAM_108_WIDTH),
        .S_AXIS_BRAM_109_WIDTH(S_AXIS_BRAM_109_WIDTH),
        .S_AXIS_BRAM_110_WIDTH(S_AXIS_BRAM_110_WIDTH),
        .S_AXIS_BRAM_111_WIDTH(S_AXIS_BRAM_111_WIDTH),
        .S_AXIS_BRAM_112_WIDTH(S_AXIS_BRAM_112_WIDTH),
        .S_AXIS_BRAM_113_WIDTH(S_AXIS_BRAM_113_WIDTH),
        .S_AXIS_BRAM_114_WIDTH(S_AXIS_BRAM_114_WIDTH),
        .S_AXIS_BRAM_115_WIDTH(S_AXIS_BRAM_115_WIDTH),
        .S_AXIS_BRAM_116_WIDTH(S_AXIS_BRAM_116_WIDTH),
        .S_AXIS_BRAM_117_WIDTH(S_AXIS_BRAM_117_WIDTH),
        .S_AXIS_BRAM_118_WIDTH(S_AXIS_BRAM_118_WIDTH),
        .S_AXIS_BRAM_119_WIDTH(S_AXIS_BRAM_119_WIDTH),
        .S_AXIS_BRAM_120_WIDTH(S_AXIS_BRAM_120_WIDTH),
        .S_AXIS_BRAM_121_WIDTH(S_AXIS_BRAM_121_WIDTH),
        .S_AXIS_BRAM_122_WIDTH(S_AXIS_BRAM_122_WIDTH),
        .S_AXIS_BRAM_123_WIDTH(S_AXIS_BRAM_123_WIDTH),
        .S_AXIS_BRAM_124_WIDTH(S_AXIS_BRAM_124_WIDTH),
        .S_AXIS_BRAM_125_WIDTH(S_AXIS_BRAM_125_WIDTH),
        .S_AXIS_BRAM_126_WIDTH(S_AXIS_BRAM_126_WIDTH),
        .S_AXIS_BRAM_127_WIDTH(S_AXIS_BRAM_127_WIDTH),
        .S_AXIS_BRAM_0_DEPTH(S_AXIS_BRAM_0_DEPTH),
        .S_AXIS_BRAM_1_DEPTH(S_AXIS_BRAM_1_DEPTH),
        .S_AXIS_BRAM_2_DEPTH(S_AXIS_BRAM_2_DEPTH),
        .S_AXIS_BRAM_3_DEPTH(S_AXIS_BRAM_3_DEPTH),
        .S_AXIS_BRAM_4_DEPTH(S_AXIS_BRAM_4_DEPTH),
        .S_AXIS_BRAM_5_DEPTH(S_AXIS_BRAM_5_DEPTH),
        .S_AXIS_BRAM_6_DEPTH(S_AXIS_BRAM_6_DEPTH),
        .S_AXIS_BRAM_7_DEPTH(S_AXIS_BRAM_7_DEPTH),
        .S_AXIS_BRAM_8_DEPTH(S_AXIS_BRAM_8_DEPTH),
        .S_AXIS_BRAM_9_DEPTH(S_AXIS_BRAM_9_DEPTH),
        .S_AXIS_BRAM_10_DEPTH(S_AXIS_BRAM_10_DEPTH),
        .S_AXIS_BRAM_11_DEPTH(S_AXIS_BRAM_11_DEPTH),
        .S_AXIS_BRAM_12_DEPTH(S_AXIS_BRAM_12_DEPTH),
        .S_AXIS_BRAM_13_DEPTH(S_AXIS_BRAM_13_DEPTH),
        .S_AXIS_BRAM_14_DEPTH(S_AXIS_BRAM_14_DEPTH),
        .S_AXIS_BRAM_15_DEPTH(S_AXIS_BRAM_15_DEPTH),
        .S_AXIS_BRAM_16_DEPTH(S_AXIS_BRAM_16_DEPTH),
        .S_AXIS_BRAM_17_DEPTH(S_AXIS_BRAM_17_DEPTH),
        .S_AXIS_BRAM_18_DEPTH(S_AXIS_BRAM_18_DEPTH),
        .S_AXIS_BRAM_19_DEPTH(S_AXIS_BRAM_19_DEPTH),
        .S_AXIS_BRAM_20_DEPTH(S_AXIS_BRAM_20_DEPTH),
        .S_AXIS_BRAM_21_DEPTH(S_AXIS_BRAM_21_DEPTH),
        .S_AXIS_BRAM_22_DEPTH(S_AXIS_BRAM_22_DEPTH),
        .S_AXIS_BRAM_23_DEPTH(S_AXIS_BRAM_23_DEPTH),
        .S_AXIS_BRAM_24_DEPTH(S_AXIS_BRAM_24_DEPTH),
        .S_AXIS_BRAM_25_DEPTH(S_AXIS_BRAM_25_DEPTH),
        .S_AXIS_BRAM_26_DEPTH(S_AXIS_BRAM_26_DEPTH),
        .S_AXIS_BRAM_27_DEPTH(S_AXIS_BRAM_27_DEPTH),
        .S_AXIS_BRAM_28_DEPTH(S_AXIS_BRAM_28_DEPTH),
        .S_AXIS_BRAM_29_DEPTH(S_AXIS_BRAM_29_DEPTH),
        .S_AXIS_BRAM_30_DEPTH(S_AXIS_BRAM_30_DEPTH),
        .S_AXIS_BRAM_31_DEPTH(S_AXIS_BRAM_31_DEPTH),
        .S_AXIS_BRAM_32_DEPTH(S_AXIS_BRAM_32_DEPTH),
        .S_AXIS_BRAM_33_DEPTH(S_AXIS_BRAM_33_DEPTH),
        .S_AXIS_BRAM_34_DEPTH(S_AXIS_BRAM_34_DEPTH),
        .S_AXIS_BRAM_35_DEPTH(S_AXIS_BRAM_35_DEPTH),
        .S_AXIS_BRAM_36_DEPTH(S_AXIS_BRAM_36_DEPTH),
        .S_AXIS_BRAM_37_DEPTH(S_AXIS_BRAM_37_DEPTH),
        .S_AXIS_BRAM_38_DEPTH(S_AXIS_BRAM_38_DEPTH),
        .S_AXIS_BRAM_39_DEPTH(S_AXIS_BRAM_39_DEPTH),
        .S_AXIS_BRAM_40_DEPTH(S_AXIS_BRAM_40_DEPTH),
        .S_AXIS_BRAM_41_DEPTH(S_AXIS_BRAM_41_DEPTH),
        .S_AXIS_BRAM_42_DEPTH(S_AXIS_BRAM_42_DEPTH),
        .S_AXIS_BRAM_43_DEPTH(S_AXIS_BRAM_43_DEPTH),
        .S_AXIS_BRAM_44_DEPTH(S_AXIS_BRAM_44_DEPTH),
        .S_AXIS_BRAM_45_DEPTH(S_AXIS_BRAM_45_DEPTH),
        .S_AXIS_BRAM_46_DEPTH(S_AXIS_BRAM_46_DEPTH),
        .S_AXIS_BRAM_47_DEPTH(S_AXIS_BRAM_47_DEPTH),
        .S_AXIS_BRAM_48_DEPTH(S_AXIS_BRAM_48_DEPTH),
        .S_AXIS_BRAM_49_DEPTH(S_AXIS_BRAM_49_DEPTH),
        .S_AXIS_BRAM_50_DEPTH(S_AXIS_BRAM_50_DEPTH),
        .S_AXIS_BRAM_51_DEPTH(S_AXIS_BRAM_51_DEPTH),
        .S_AXIS_BRAM_52_DEPTH(S_AXIS_BRAM_52_DEPTH),
        .S_AXIS_BRAM_53_DEPTH(S_AXIS_BRAM_53_DEPTH),
        .S_AXIS_BRAM_54_DEPTH(S_AXIS_BRAM_54_DEPTH),
        .S_AXIS_BRAM_55_DEPTH(S_AXIS_BRAM_55_DEPTH),
        .S_AXIS_BRAM_56_DEPTH(S_AXIS_BRAM_56_DEPTH),
        .S_AXIS_BRAM_57_DEPTH(S_AXIS_BRAM_57_DEPTH),
        .S_AXIS_BRAM_58_DEPTH(S_AXIS_BRAM_58_DEPTH),
        .S_AXIS_BRAM_59_DEPTH(S_AXIS_BRAM_59_DEPTH),
        .S_AXIS_BRAM_60_DEPTH(S_AXIS_BRAM_60_DEPTH),
        .S_AXIS_BRAM_61_DEPTH(S_AXIS_BRAM_61_DEPTH),
        .S_AXIS_BRAM_62_DEPTH(S_AXIS_BRAM_62_DEPTH),
        .S_AXIS_BRAM_63_DEPTH(S_AXIS_BRAM_63_DEPTH),
        .S_AXIS_BRAM_64_DEPTH(S_AXIS_BRAM_64_DEPTH),
        .S_AXIS_BRAM_65_DEPTH(S_AXIS_BRAM_65_DEPTH),
        .S_AXIS_BRAM_66_DEPTH(S_AXIS_BRAM_66_DEPTH),
        .S_AXIS_BRAM_67_DEPTH(S_AXIS_BRAM_67_DEPTH),
        .S_AXIS_BRAM_68_DEPTH(S_AXIS_BRAM_68_DEPTH),
        .S_AXIS_BRAM_69_DEPTH(S_AXIS_BRAM_69_DEPTH),
        .S_AXIS_BRAM_70_DEPTH(S_AXIS_BRAM_70_DEPTH),
        .S_AXIS_BRAM_71_DEPTH(S_AXIS_BRAM_71_DEPTH),
        .S_AXIS_BRAM_72_DEPTH(S_AXIS_BRAM_72_DEPTH),
        .S_AXIS_BRAM_73_DEPTH(S_AXIS_BRAM_73_DEPTH),
        .S_AXIS_BRAM_74_DEPTH(S_AXIS_BRAM_74_DEPTH),
        .S_AXIS_BRAM_75_DEPTH(S_AXIS_BRAM_75_DEPTH),
        .S_AXIS_BRAM_76_DEPTH(S_AXIS_BRAM_76_DEPTH),
        .S_AXIS_BRAM_77_DEPTH(S_AXIS_BRAM_77_DEPTH),
        .S_AXIS_BRAM_78_DEPTH(S_AXIS_BRAM_78_DEPTH),
        .S_AXIS_BRAM_79_DEPTH(S_AXIS_BRAM_79_DEPTH),
        .S_AXIS_BRAM_80_DEPTH(S_AXIS_BRAM_80_DEPTH),
        .S_AXIS_BRAM_81_DEPTH(S_AXIS_BRAM_81_DEPTH),
        .S_AXIS_BRAM_82_DEPTH(S_AXIS_BRAM_82_DEPTH),
        .S_AXIS_BRAM_83_DEPTH(S_AXIS_BRAM_83_DEPTH),
        .S_AXIS_BRAM_84_DEPTH(S_AXIS_BRAM_84_DEPTH),
        .S_AXIS_BRAM_85_DEPTH(S_AXIS_BRAM_85_DEPTH),
        .S_AXIS_BRAM_86_DEPTH(S_AXIS_BRAM_86_DEPTH),
        .S_AXIS_BRAM_87_DEPTH(S_AXIS_BRAM_87_DEPTH),
        .S_AXIS_BRAM_88_DEPTH(S_AXIS_BRAM_88_DEPTH),
        .S_AXIS_BRAM_89_DEPTH(S_AXIS_BRAM_89_DEPTH),
        .S_AXIS_BRAM_90_DEPTH(S_AXIS_BRAM_90_DEPTH),
        .S_AXIS_BRAM_91_DEPTH(S_AXIS_BRAM_91_DEPTH),
        .S_AXIS_BRAM_92_DEPTH(S_AXIS_BRAM_92_DEPTH),
        .S_AXIS_BRAM_93_DEPTH(S_AXIS_BRAM_93_DEPTH),
        .S_AXIS_BRAM_94_DEPTH(S_AXIS_BRAM_94_DEPTH),
        .S_AXIS_BRAM_95_DEPTH(S_AXIS_BRAM_95_DEPTH),
        .S_AXIS_BRAM_96_DEPTH(S_AXIS_BRAM_96_DEPTH),
        .S_AXIS_BRAM_97_DEPTH(S_AXIS_BRAM_97_DEPTH),
        .S_AXIS_BRAM_98_DEPTH(S_AXIS_BRAM_98_DEPTH),
        .S_AXIS_BRAM_99_DEPTH(S_AXIS_BRAM_99_DEPTH),
        .S_AXIS_BRAM_100_DEPTH(S_AXIS_BRAM_100_DEPTH),
        .S_AXIS_BRAM_101_DEPTH(S_AXIS_BRAM_101_DEPTH),
        .S_AXIS_BRAM_102_DEPTH(S_AXIS_BRAM_102_DEPTH),
        .S_AXIS_BRAM_103_DEPTH(S_AXIS_BRAM_103_DEPTH),
        .S_AXIS_BRAM_104_DEPTH(S_AXIS_BRAM_104_DEPTH),
        .S_AXIS_BRAM_105_DEPTH(S_AXIS_BRAM_105_DEPTH),
        .S_AXIS_BRAM_106_DEPTH(S_AXIS_BRAM_106_DEPTH),
        .S_AXIS_BRAM_107_DEPTH(S_AXIS_BRAM_107_DEPTH),
        .S_AXIS_BRAM_108_DEPTH(S_AXIS_BRAM_108_DEPTH),
        .S_AXIS_BRAM_109_DEPTH(S_AXIS_BRAM_109_DEPTH),
        .S_AXIS_BRAM_110_DEPTH(S_AXIS_BRAM_110_DEPTH),
        .S_AXIS_BRAM_111_DEPTH(S_AXIS_BRAM_111_DEPTH),
        .S_AXIS_BRAM_112_DEPTH(S_AXIS_BRAM_112_DEPTH),
        .S_AXIS_BRAM_113_DEPTH(S_AXIS_BRAM_113_DEPTH),
        .S_AXIS_BRAM_114_DEPTH(S_AXIS_BRAM_114_DEPTH),
        .S_AXIS_BRAM_115_DEPTH(S_AXIS_BRAM_115_DEPTH),
        .S_AXIS_BRAM_116_DEPTH(S_AXIS_BRAM_116_DEPTH),
        .S_AXIS_BRAM_117_DEPTH(S_AXIS_BRAM_117_DEPTH),
        .S_AXIS_BRAM_118_DEPTH(S_AXIS_BRAM_118_DEPTH),
        .S_AXIS_BRAM_119_DEPTH(S_AXIS_BRAM_119_DEPTH),
        .S_AXIS_BRAM_120_DEPTH(S_AXIS_BRAM_120_DEPTH),
        .S_AXIS_BRAM_121_DEPTH(S_AXIS_BRAM_121_DEPTH),
        .S_AXIS_BRAM_122_DEPTH(S_AXIS_BRAM_122_DEPTH),
        .S_AXIS_BRAM_123_DEPTH(S_AXIS_BRAM_123_DEPTH),
        .S_AXIS_BRAM_124_DEPTH(S_AXIS_BRAM_124_DEPTH),
        .S_AXIS_BRAM_125_DEPTH(S_AXIS_BRAM_125_DEPTH),
        .S_AXIS_BRAM_126_DEPTH(S_AXIS_BRAM_126_DEPTH),
        .S_AXIS_BRAM_127_DEPTH(S_AXIS_BRAM_127_DEPTH),
        .S_AXIS_BRAM_0_DMWIDTH(S_AXIS_BRAM_0_DMWIDTH),
        .S_AXIS_BRAM_1_DMWIDTH(S_AXIS_BRAM_1_DMWIDTH),
        .S_AXIS_BRAM_2_DMWIDTH(S_AXIS_BRAM_2_DMWIDTH),
        .S_AXIS_BRAM_3_DMWIDTH(S_AXIS_BRAM_3_DMWIDTH),
        .S_AXIS_BRAM_4_DMWIDTH(S_AXIS_BRAM_4_DMWIDTH),
        .S_AXIS_BRAM_5_DMWIDTH(S_AXIS_BRAM_5_DMWIDTH),
        .S_AXIS_BRAM_6_DMWIDTH(S_AXIS_BRAM_6_DMWIDTH),
        .S_AXIS_BRAM_7_DMWIDTH(S_AXIS_BRAM_7_DMWIDTH),
        .S_AXIS_BRAM_8_DMWIDTH(S_AXIS_BRAM_8_DMWIDTH),
        .S_AXIS_BRAM_9_DMWIDTH(S_AXIS_BRAM_9_DMWIDTH),
        .S_AXIS_BRAM_10_DMWIDTH(S_AXIS_BRAM_10_DMWIDTH),
        .S_AXIS_BRAM_11_DMWIDTH(S_AXIS_BRAM_11_DMWIDTH),
        .S_AXIS_BRAM_12_DMWIDTH(S_AXIS_BRAM_12_DMWIDTH),
        .S_AXIS_BRAM_13_DMWIDTH(S_AXIS_BRAM_13_DMWIDTH),
        .S_AXIS_BRAM_14_DMWIDTH(S_AXIS_BRAM_14_DMWIDTH),
        .S_AXIS_BRAM_15_DMWIDTH(S_AXIS_BRAM_15_DMWIDTH),
        .S_AXIS_BRAM_16_DMWIDTH(S_AXIS_BRAM_16_DMWIDTH),
        .S_AXIS_BRAM_17_DMWIDTH(S_AXIS_BRAM_17_DMWIDTH),
        .S_AXIS_BRAM_18_DMWIDTH(S_AXIS_BRAM_18_DMWIDTH),
        .S_AXIS_BRAM_19_DMWIDTH(S_AXIS_BRAM_19_DMWIDTH),
        .S_AXIS_BRAM_20_DMWIDTH(S_AXIS_BRAM_20_DMWIDTH),
        .S_AXIS_BRAM_21_DMWIDTH(S_AXIS_BRAM_21_DMWIDTH),
        .S_AXIS_BRAM_22_DMWIDTH(S_AXIS_BRAM_22_DMWIDTH),
        .S_AXIS_BRAM_23_DMWIDTH(S_AXIS_BRAM_23_DMWIDTH),
        .S_AXIS_BRAM_24_DMWIDTH(S_AXIS_BRAM_24_DMWIDTH),
        .S_AXIS_BRAM_25_DMWIDTH(S_AXIS_BRAM_25_DMWIDTH),
        .S_AXIS_BRAM_26_DMWIDTH(S_AXIS_BRAM_26_DMWIDTH),
        .S_AXIS_BRAM_27_DMWIDTH(S_AXIS_BRAM_27_DMWIDTH),
        .S_AXIS_BRAM_28_DMWIDTH(S_AXIS_BRAM_28_DMWIDTH),
        .S_AXIS_BRAM_29_DMWIDTH(S_AXIS_BRAM_29_DMWIDTH),
        .S_AXIS_BRAM_30_DMWIDTH(S_AXIS_BRAM_30_DMWIDTH),
        .S_AXIS_BRAM_31_DMWIDTH(S_AXIS_BRAM_31_DMWIDTH),
        .S_AXIS_BRAM_32_DMWIDTH(S_AXIS_BRAM_32_DMWIDTH),
        .S_AXIS_BRAM_33_DMWIDTH(S_AXIS_BRAM_33_DMWIDTH),
        .S_AXIS_BRAM_34_DMWIDTH(S_AXIS_BRAM_34_DMWIDTH),
        .S_AXIS_BRAM_35_DMWIDTH(S_AXIS_BRAM_35_DMWIDTH),
        .S_AXIS_BRAM_36_DMWIDTH(S_AXIS_BRAM_36_DMWIDTH),
        .S_AXIS_BRAM_37_DMWIDTH(S_AXIS_BRAM_37_DMWIDTH),
        .S_AXIS_BRAM_38_DMWIDTH(S_AXIS_BRAM_38_DMWIDTH),
        .S_AXIS_BRAM_39_DMWIDTH(S_AXIS_BRAM_39_DMWIDTH),
        .S_AXIS_BRAM_40_DMWIDTH(S_AXIS_BRAM_40_DMWIDTH),
        .S_AXIS_BRAM_41_DMWIDTH(S_AXIS_BRAM_41_DMWIDTH),
        .S_AXIS_BRAM_42_DMWIDTH(S_AXIS_BRAM_42_DMWIDTH),
        .S_AXIS_BRAM_43_DMWIDTH(S_AXIS_BRAM_43_DMWIDTH),
        .S_AXIS_BRAM_44_DMWIDTH(S_AXIS_BRAM_44_DMWIDTH),
        .S_AXIS_BRAM_45_DMWIDTH(S_AXIS_BRAM_45_DMWIDTH),
        .S_AXIS_BRAM_46_DMWIDTH(S_AXIS_BRAM_46_DMWIDTH),
        .S_AXIS_BRAM_47_DMWIDTH(S_AXIS_BRAM_47_DMWIDTH),
        .S_AXIS_BRAM_48_DMWIDTH(S_AXIS_BRAM_48_DMWIDTH),
        .S_AXIS_BRAM_49_DMWIDTH(S_AXIS_BRAM_49_DMWIDTH),
        .S_AXIS_BRAM_50_DMWIDTH(S_AXIS_BRAM_50_DMWIDTH),
        .S_AXIS_BRAM_51_DMWIDTH(S_AXIS_BRAM_51_DMWIDTH),
        .S_AXIS_BRAM_52_DMWIDTH(S_AXIS_BRAM_52_DMWIDTH),
        .S_AXIS_BRAM_53_DMWIDTH(S_AXIS_BRAM_53_DMWIDTH),
        .S_AXIS_BRAM_54_DMWIDTH(S_AXIS_BRAM_54_DMWIDTH),
        .S_AXIS_BRAM_55_DMWIDTH(S_AXIS_BRAM_55_DMWIDTH),
        .S_AXIS_BRAM_56_DMWIDTH(S_AXIS_BRAM_56_DMWIDTH),
        .S_AXIS_BRAM_57_DMWIDTH(S_AXIS_BRAM_57_DMWIDTH),
        .S_AXIS_BRAM_58_DMWIDTH(S_AXIS_BRAM_58_DMWIDTH),
        .S_AXIS_BRAM_59_DMWIDTH(S_AXIS_BRAM_59_DMWIDTH),
        .S_AXIS_BRAM_60_DMWIDTH(S_AXIS_BRAM_60_DMWIDTH),
        .S_AXIS_BRAM_61_DMWIDTH(S_AXIS_BRAM_61_DMWIDTH),
        .S_AXIS_BRAM_62_DMWIDTH(S_AXIS_BRAM_62_DMWIDTH),
        .S_AXIS_BRAM_63_DMWIDTH(S_AXIS_BRAM_63_DMWIDTH),
        .S_AXIS_BRAM_64_DMWIDTH(S_AXIS_BRAM_64_DMWIDTH),
        .S_AXIS_BRAM_65_DMWIDTH(S_AXIS_BRAM_65_DMWIDTH),
        .S_AXIS_BRAM_66_DMWIDTH(S_AXIS_BRAM_66_DMWIDTH),
        .S_AXIS_BRAM_67_DMWIDTH(S_AXIS_BRAM_67_DMWIDTH),
        .S_AXIS_BRAM_68_DMWIDTH(S_AXIS_BRAM_68_DMWIDTH),
        .S_AXIS_BRAM_69_DMWIDTH(S_AXIS_BRAM_69_DMWIDTH),
        .S_AXIS_BRAM_70_DMWIDTH(S_AXIS_BRAM_70_DMWIDTH),
        .S_AXIS_BRAM_71_DMWIDTH(S_AXIS_BRAM_71_DMWIDTH),
        .S_AXIS_BRAM_72_DMWIDTH(S_AXIS_BRAM_72_DMWIDTH),
        .S_AXIS_BRAM_73_DMWIDTH(S_AXIS_BRAM_73_DMWIDTH),
        .S_AXIS_BRAM_74_DMWIDTH(S_AXIS_BRAM_74_DMWIDTH),
        .S_AXIS_BRAM_75_DMWIDTH(S_AXIS_BRAM_75_DMWIDTH),
        .S_AXIS_BRAM_76_DMWIDTH(S_AXIS_BRAM_76_DMWIDTH),
        .S_AXIS_BRAM_77_DMWIDTH(S_AXIS_BRAM_77_DMWIDTH),
        .S_AXIS_BRAM_78_DMWIDTH(S_AXIS_BRAM_78_DMWIDTH),
        .S_AXIS_BRAM_79_DMWIDTH(S_AXIS_BRAM_79_DMWIDTH),
        .S_AXIS_BRAM_80_DMWIDTH(S_AXIS_BRAM_80_DMWIDTH),
        .S_AXIS_BRAM_81_DMWIDTH(S_AXIS_BRAM_81_DMWIDTH),
        .S_AXIS_BRAM_82_DMWIDTH(S_AXIS_BRAM_82_DMWIDTH),
        .S_AXIS_BRAM_83_DMWIDTH(S_AXIS_BRAM_83_DMWIDTH),
        .S_AXIS_BRAM_84_DMWIDTH(S_AXIS_BRAM_84_DMWIDTH),
        .S_AXIS_BRAM_85_DMWIDTH(S_AXIS_BRAM_85_DMWIDTH),
        .S_AXIS_BRAM_86_DMWIDTH(S_AXIS_BRAM_86_DMWIDTH),
        .S_AXIS_BRAM_87_DMWIDTH(S_AXIS_BRAM_87_DMWIDTH),
        .S_AXIS_BRAM_88_DMWIDTH(S_AXIS_BRAM_88_DMWIDTH),
        .S_AXIS_BRAM_89_DMWIDTH(S_AXIS_BRAM_89_DMWIDTH),
        .S_AXIS_BRAM_90_DMWIDTH(S_AXIS_BRAM_90_DMWIDTH),
        .S_AXIS_BRAM_91_DMWIDTH(S_AXIS_BRAM_91_DMWIDTH),
        .S_AXIS_BRAM_92_DMWIDTH(S_AXIS_BRAM_92_DMWIDTH),
        .S_AXIS_BRAM_93_DMWIDTH(S_AXIS_BRAM_93_DMWIDTH),
        .S_AXIS_BRAM_94_DMWIDTH(S_AXIS_BRAM_94_DMWIDTH),
        .S_AXIS_BRAM_95_DMWIDTH(S_AXIS_BRAM_95_DMWIDTH),
        .S_AXIS_BRAM_96_DMWIDTH(S_AXIS_BRAM_96_DMWIDTH),
        .S_AXIS_BRAM_97_DMWIDTH(S_AXIS_BRAM_97_DMWIDTH),
        .S_AXIS_BRAM_98_DMWIDTH(S_AXIS_BRAM_98_DMWIDTH),
        .S_AXIS_BRAM_99_DMWIDTH(S_AXIS_BRAM_99_DMWIDTH),
        .S_AXIS_BRAM_100_DMWIDTH(S_AXIS_BRAM_100_DMWIDTH),
        .S_AXIS_BRAM_101_DMWIDTH(S_AXIS_BRAM_101_DMWIDTH),
        .S_AXIS_BRAM_102_DMWIDTH(S_AXIS_BRAM_102_DMWIDTH),
        .S_AXIS_BRAM_103_DMWIDTH(S_AXIS_BRAM_103_DMWIDTH),
        .S_AXIS_BRAM_104_DMWIDTH(S_AXIS_BRAM_104_DMWIDTH),
        .S_AXIS_BRAM_105_DMWIDTH(S_AXIS_BRAM_105_DMWIDTH),
        .S_AXIS_BRAM_106_DMWIDTH(S_AXIS_BRAM_106_DMWIDTH),
        .S_AXIS_BRAM_107_DMWIDTH(S_AXIS_BRAM_107_DMWIDTH),
        .S_AXIS_BRAM_108_DMWIDTH(S_AXIS_BRAM_108_DMWIDTH),
        .S_AXIS_BRAM_109_DMWIDTH(S_AXIS_BRAM_109_DMWIDTH),
        .S_AXIS_BRAM_110_DMWIDTH(S_AXIS_BRAM_110_DMWIDTH),
        .S_AXIS_BRAM_111_DMWIDTH(S_AXIS_BRAM_111_DMWIDTH),
        .S_AXIS_BRAM_112_DMWIDTH(S_AXIS_BRAM_112_DMWIDTH),
        .S_AXIS_BRAM_113_DMWIDTH(S_AXIS_BRAM_113_DMWIDTH),
        .S_AXIS_BRAM_114_DMWIDTH(S_AXIS_BRAM_114_DMWIDTH),
        .S_AXIS_BRAM_115_DMWIDTH(S_AXIS_BRAM_115_DMWIDTH),
        .S_AXIS_BRAM_116_DMWIDTH(S_AXIS_BRAM_116_DMWIDTH),
        .S_AXIS_BRAM_117_DMWIDTH(S_AXIS_BRAM_117_DMWIDTH),
        .S_AXIS_BRAM_118_DMWIDTH(S_AXIS_BRAM_118_DMWIDTH),
        .S_AXIS_BRAM_119_DMWIDTH(S_AXIS_BRAM_119_DMWIDTH),
        .S_AXIS_BRAM_120_DMWIDTH(S_AXIS_BRAM_120_DMWIDTH),
        .S_AXIS_BRAM_121_DMWIDTH(S_AXIS_BRAM_121_DMWIDTH),
        .S_AXIS_BRAM_122_DMWIDTH(S_AXIS_BRAM_122_DMWIDTH),
        .S_AXIS_BRAM_123_DMWIDTH(S_AXIS_BRAM_123_DMWIDTH),
        .S_AXIS_BRAM_124_DMWIDTH(S_AXIS_BRAM_124_DMWIDTH),
        .S_AXIS_BRAM_125_DMWIDTH(S_AXIS_BRAM_125_DMWIDTH),
        .S_AXIS_BRAM_126_DMWIDTH(S_AXIS_BRAM_126_DMWIDTH),
        .S_AXIS_BRAM_127_DMWIDTH(S_AXIS_BRAM_127_DMWIDTH),
        .M_AXIS_BRAMIO_0_DMWIDTH(M_AXIS_BRAMIO_0_DMWIDTH),
        .M_AXIS_BRAMIO_1_DMWIDTH(M_AXIS_BRAMIO_1_DMWIDTH),
        .M_AXIS_BRAMIO_2_DMWIDTH(M_AXIS_BRAMIO_2_DMWIDTH),
        .M_AXIS_BRAMIO_3_DMWIDTH(M_AXIS_BRAMIO_3_DMWIDTH),
        .M_AXIS_BRAMIO_4_DMWIDTH(M_AXIS_BRAMIO_4_DMWIDTH),
        .M_AXIS_BRAMIO_5_DMWIDTH(M_AXIS_BRAMIO_5_DMWIDTH),
        .M_AXIS_BRAMIO_6_DMWIDTH(M_AXIS_BRAMIO_6_DMWIDTH),
        .M_AXIS_BRAMIO_7_DMWIDTH(M_AXIS_BRAMIO_7_DMWIDTH),
        .M_AXIS_BRAMIO_8_DMWIDTH(M_AXIS_BRAMIO_8_DMWIDTH),
        .M_AXIS_BRAMIO_9_DMWIDTH(M_AXIS_BRAMIO_9_DMWIDTH),
        .M_AXIS_BRAMIO_10_DMWIDTH(M_AXIS_BRAMIO_10_DMWIDTH),
        .M_AXIS_BRAMIO_11_DMWIDTH(M_AXIS_BRAMIO_11_DMWIDTH),
        .M_AXIS_BRAMIO_12_DMWIDTH(M_AXIS_BRAMIO_12_DMWIDTH),
        .M_AXIS_BRAMIO_13_DMWIDTH(M_AXIS_BRAMIO_13_DMWIDTH),
        .M_AXIS_BRAMIO_14_DMWIDTH(M_AXIS_BRAMIO_14_DMWIDTH),
        .M_AXIS_BRAMIO_15_DMWIDTH(M_AXIS_BRAMIO_15_DMWIDTH),
        .M_AXIS_BRAMIO_16_DMWIDTH(M_AXIS_BRAMIO_16_DMWIDTH),
        .M_AXIS_BRAMIO_17_DMWIDTH(M_AXIS_BRAMIO_17_DMWIDTH),
        .M_AXIS_BRAMIO_18_DMWIDTH(M_AXIS_BRAMIO_18_DMWIDTH),
        .M_AXIS_BRAMIO_19_DMWIDTH(M_AXIS_BRAMIO_19_DMWIDTH),
        .M_AXIS_BRAMIO_20_DMWIDTH(M_AXIS_BRAMIO_20_DMWIDTH),
        .M_AXIS_BRAMIO_21_DMWIDTH(M_AXIS_BRAMIO_21_DMWIDTH),
        .M_AXIS_BRAMIO_22_DMWIDTH(M_AXIS_BRAMIO_22_DMWIDTH),
        .M_AXIS_BRAMIO_23_DMWIDTH(M_AXIS_BRAMIO_23_DMWIDTH),
        .M_AXIS_BRAMIO_24_DMWIDTH(M_AXIS_BRAMIO_24_DMWIDTH),
        .M_AXIS_BRAMIO_25_DMWIDTH(M_AXIS_BRAMIO_25_DMWIDTH),
        .M_AXIS_BRAMIO_26_DMWIDTH(M_AXIS_BRAMIO_26_DMWIDTH),
        .M_AXIS_BRAMIO_27_DMWIDTH(M_AXIS_BRAMIO_27_DMWIDTH),
        .M_AXIS_BRAMIO_28_DMWIDTH(M_AXIS_BRAMIO_28_DMWIDTH),
        .M_AXIS_BRAMIO_29_DMWIDTH(M_AXIS_BRAMIO_29_DMWIDTH),
        .M_AXIS_BRAMIO_30_DMWIDTH(M_AXIS_BRAMIO_30_DMWIDTH),
        .M_AXIS_BRAMIO_31_DMWIDTH(M_AXIS_BRAMIO_31_DMWIDTH),
        .M_AXIS_BRAMIO_32_DMWIDTH(M_AXIS_BRAMIO_32_DMWIDTH),
        .M_AXIS_BRAMIO_33_DMWIDTH(M_AXIS_BRAMIO_33_DMWIDTH),
        .M_AXIS_BRAMIO_34_DMWIDTH(M_AXIS_BRAMIO_34_DMWIDTH),
        .M_AXIS_BRAMIO_35_DMWIDTH(M_AXIS_BRAMIO_35_DMWIDTH),
        .M_AXIS_BRAMIO_36_DMWIDTH(M_AXIS_BRAMIO_36_DMWIDTH),
        .M_AXIS_BRAMIO_37_DMWIDTH(M_AXIS_BRAMIO_37_DMWIDTH),
        .M_AXIS_BRAMIO_38_DMWIDTH(M_AXIS_BRAMIO_38_DMWIDTH),
        .M_AXIS_BRAMIO_39_DMWIDTH(M_AXIS_BRAMIO_39_DMWIDTH),
        .M_AXIS_BRAMIO_40_DMWIDTH(M_AXIS_BRAMIO_40_DMWIDTH),
        .M_AXIS_BRAMIO_41_DMWIDTH(M_AXIS_BRAMIO_41_DMWIDTH),
        .M_AXIS_BRAMIO_42_DMWIDTH(M_AXIS_BRAMIO_42_DMWIDTH),
        .M_AXIS_BRAMIO_43_DMWIDTH(M_AXIS_BRAMIO_43_DMWIDTH),
        .M_AXIS_BRAMIO_44_DMWIDTH(M_AXIS_BRAMIO_44_DMWIDTH),
        .M_AXIS_BRAMIO_45_DMWIDTH(M_AXIS_BRAMIO_45_DMWIDTH),
        .M_AXIS_BRAMIO_46_DMWIDTH(M_AXIS_BRAMIO_46_DMWIDTH),
        .M_AXIS_BRAMIO_47_DMWIDTH(M_AXIS_BRAMIO_47_DMWIDTH),
        .M_AXIS_BRAMIO_48_DMWIDTH(M_AXIS_BRAMIO_48_DMWIDTH),
        .M_AXIS_BRAMIO_49_DMWIDTH(M_AXIS_BRAMIO_49_DMWIDTH),
        .M_AXIS_BRAMIO_50_DMWIDTH(M_AXIS_BRAMIO_50_DMWIDTH),
        .M_AXIS_BRAMIO_51_DMWIDTH(M_AXIS_BRAMIO_51_DMWIDTH),
        .M_AXIS_BRAMIO_52_DMWIDTH(M_AXIS_BRAMIO_52_DMWIDTH),
        .M_AXIS_BRAMIO_53_DMWIDTH(M_AXIS_BRAMIO_53_DMWIDTH),
        .M_AXIS_BRAMIO_54_DMWIDTH(M_AXIS_BRAMIO_54_DMWIDTH),
        .M_AXIS_BRAMIO_55_DMWIDTH(M_AXIS_BRAMIO_55_DMWIDTH),
        .M_AXIS_BRAMIO_56_DMWIDTH(M_AXIS_BRAMIO_56_DMWIDTH),
        .M_AXIS_BRAMIO_57_DMWIDTH(M_AXIS_BRAMIO_57_DMWIDTH),
        .M_AXIS_BRAMIO_58_DMWIDTH(M_AXIS_BRAMIO_58_DMWIDTH),
        .M_AXIS_BRAMIO_59_DMWIDTH(M_AXIS_BRAMIO_59_DMWIDTH),
        .M_AXIS_BRAMIO_60_DMWIDTH(M_AXIS_BRAMIO_60_DMWIDTH),
        .M_AXIS_BRAMIO_61_DMWIDTH(M_AXIS_BRAMIO_61_DMWIDTH),
        .M_AXIS_BRAMIO_62_DMWIDTH(M_AXIS_BRAMIO_62_DMWIDTH),
        .M_AXIS_BRAMIO_63_DMWIDTH(M_AXIS_BRAMIO_63_DMWIDTH),
        .M_AXIS_BRAMIO_64_DMWIDTH(M_AXIS_BRAMIO_64_DMWIDTH),
        .M_AXIS_BRAMIO_65_DMWIDTH(M_AXIS_BRAMIO_65_DMWIDTH),
        .M_AXIS_BRAMIO_66_DMWIDTH(M_AXIS_BRAMIO_66_DMWIDTH),
        .M_AXIS_BRAMIO_67_DMWIDTH(M_AXIS_BRAMIO_67_DMWIDTH),
        .M_AXIS_BRAMIO_68_DMWIDTH(M_AXIS_BRAMIO_68_DMWIDTH),
        .M_AXIS_BRAMIO_69_DMWIDTH(M_AXIS_BRAMIO_69_DMWIDTH),
        .M_AXIS_BRAMIO_70_DMWIDTH(M_AXIS_BRAMIO_70_DMWIDTH),
        .M_AXIS_BRAMIO_71_DMWIDTH(M_AXIS_BRAMIO_71_DMWIDTH),
        .M_AXIS_BRAMIO_72_DMWIDTH(M_AXIS_BRAMIO_72_DMWIDTH),
        .M_AXIS_BRAMIO_73_DMWIDTH(M_AXIS_BRAMIO_73_DMWIDTH),
        .M_AXIS_BRAMIO_74_DMWIDTH(M_AXIS_BRAMIO_74_DMWIDTH),
        .M_AXIS_BRAMIO_75_DMWIDTH(M_AXIS_BRAMIO_75_DMWIDTH),
        .M_AXIS_BRAMIO_76_DMWIDTH(M_AXIS_BRAMIO_76_DMWIDTH),
        .M_AXIS_BRAMIO_77_DMWIDTH(M_AXIS_BRAMIO_77_DMWIDTH),
        .M_AXIS_BRAMIO_78_DMWIDTH(M_AXIS_BRAMIO_78_DMWIDTH),
        .M_AXIS_BRAMIO_79_DMWIDTH(M_AXIS_BRAMIO_79_DMWIDTH),
        .M_AXIS_BRAMIO_80_DMWIDTH(M_AXIS_BRAMIO_80_DMWIDTH),
        .M_AXIS_BRAMIO_81_DMWIDTH(M_AXIS_BRAMIO_81_DMWIDTH),
        .M_AXIS_BRAMIO_82_DMWIDTH(M_AXIS_BRAMIO_82_DMWIDTH),
        .M_AXIS_BRAMIO_83_DMWIDTH(M_AXIS_BRAMIO_83_DMWIDTH),
        .M_AXIS_BRAMIO_84_DMWIDTH(M_AXIS_BRAMIO_84_DMWIDTH),
        .M_AXIS_BRAMIO_85_DMWIDTH(M_AXIS_BRAMIO_85_DMWIDTH),
        .M_AXIS_BRAMIO_86_DMWIDTH(M_AXIS_BRAMIO_86_DMWIDTH),
        .M_AXIS_BRAMIO_87_DMWIDTH(M_AXIS_BRAMIO_87_DMWIDTH),
        .M_AXIS_BRAMIO_88_DMWIDTH(M_AXIS_BRAMIO_88_DMWIDTH),
        .M_AXIS_BRAMIO_89_DMWIDTH(M_AXIS_BRAMIO_89_DMWIDTH),
        .M_AXIS_BRAMIO_90_DMWIDTH(M_AXIS_BRAMIO_90_DMWIDTH),
        .M_AXIS_BRAMIO_91_DMWIDTH(M_AXIS_BRAMIO_91_DMWIDTH),
        .M_AXIS_BRAMIO_92_DMWIDTH(M_AXIS_BRAMIO_92_DMWIDTH),
        .M_AXIS_BRAMIO_93_DMWIDTH(M_AXIS_BRAMIO_93_DMWIDTH),
        .M_AXIS_BRAMIO_94_DMWIDTH(M_AXIS_BRAMIO_94_DMWIDTH),
        .M_AXIS_BRAMIO_95_DMWIDTH(M_AXIS_BRAMIO_95_DMWIDTH),
        .M_AXIS_BRAMIO_96_DMWIDTH(M_AXIS_BRAMIO_96_DMWIDTH),
        .M_AXIS_BRAMIO_97_DMWIDTH(M_AXIS_BRAMIO_97_DMWIDTH),
        .M_AXIS_BRAMIO_98_DMWIDTH(M_AXIS_BRAMIO_98_DMWIDTH),
        .M_AXIS_BRAMIO_99_DMWIDTH(M_AXIS_BRAMIO_99_DMWIDTH),
        .M_AXIS_BRAMIO_100_DMWIDTH(M_AXIS_BRAMIO_100_DMWIDTH),
        .M_AXIS_BRAMIO_101_DMWIDTH(M_AXIS_BRAMIO_101_DMWIDTH),
        .M_AXIS_BRAMIO_102_DMWIDTH(M_AXIS_BRAMIO_102_DMWIDTH),
        .M_AXIS_BRAMIO_103_DMWIDTH(M_AXIS_BRAMIO_103_DMWIDTH),
        .M_AXIS_BRAMIO_104_DMWIDTH(M_AXIS_BRAMIO_104_DMWIDTH),
        .M_AXIS_BRAMIO_105_DMWIDTH(M_AXIS_BRAMIO_105_DMWIDTH),
        .M_AXIS_BRAMIO_106_DMWIDTH(M_AXIS_BRAMIO_106_DMWIDTH),
        .M_AXIS_BRAMIO_107_DMWIDTH(M_AXIS_BRAMIO_107_DMWIDTH),
        .M_AXIS_BRAMIO_108_DMWIDTH(M_AXIS_BRAMIO_108_DMWIDTH),
        .M_AXIS_BRAMIO_109_DMWIDTH(M_AXIS_BRAMIO_109_DMWIDTH),
        .M_AXIS_BRAMIO_110_DMWIDTH(M_AXIS_BRAMIO_110_DMWIDTH),
        .M_AXIS_BRAMIO_111_DMWIDTH(M_AXIS_BRAMIO_111_DMWIDTH),
        .M_AXIS_BRAMIO_112_DMWIDTH(M_AXIS_BRAMIO_112_DMWIDTH),
        .M_AXIS_BRAMIO_113_DMWIDTH(M_AXIS_BRAMIO_113_DMWIDTH),
        .M_AXIS_BRAMIO_114_DMWIDTH(M_AXIS_BRAMIO_114_DMWIDTH),
        .M_AXIS_BRAMIO_115_DMWIDTH(M_AXIS_BRAMIO_115_DMWIDTH),
        .M_AXIS_BRAMIO_116_DMWIDTH(M_AXIS_BRAMIO_116_DMWIDTH),
        .M_AXIS_BRAMIO_117_DMWIDTH(M_AXIS_BRAMIO_117_DMWIDTH),
        .M_AXIS_BRAMIO_118_DMWIDTH(M_AXIS_BRAMIO_118_DMWIDTH),
        .M_AXIS_BRAMIO_119_DMWIDTH(M_AXIS_BRAMIO_119_DMWIDTH),
        .M_AXIS_BRAMIO_120_DMWIDTH(M_AXIS_BRAMIO_120_DMWIDTH),
        .M_AXIS_BRAMIO_121_DMWIDTH(M_AXIS_BRAMIO_121_DMWIDTH),
        .M_AXIS_BRAMIO_122_DMWIDTH(M_AXIS_BRAMIO_122_DMWIDTH),
        .M_AXIS_BRAMIO_123_DMWIDTH(M_AXIS_BRAMIO_123_DMWIDTH),
        .M_AXIS_BRAMIO_124_DMWIDTH(M_AXIS_BRAMIO_124_DMWIDTH),
        .M_AXIS_BRAMIO_125_DMWIDTH(M_AXIS_BRAMIO_125_DMWIDTH),
        .M_AXIS_BRAMIO_126_DMWIDTH(M_AXIS_BRAMIO_126_DMWIDTH),
        .M_AXIS_BRAMIO_127_DMWIDTH(M_AXIS_BRAMIO_127_DMWIDTH),
        .S_AXIS_BRAM_0_IS_ASYNC(S_AXIS_BRAM_0_IS_ASYNC),
        .S_AXIS_BRAM_1_IS_ASYNC(S_AXIS_BRAM_1_IS_ASYNC),
        .S_AXIS_BRAM_2_IS_ASYNC(S_AXIS_BRAM_2_IS_ASYNC),
        .S_AXIS_BRAM_3_IS_ASYNC(S_AXIS_BRAM_3_IS_ASYNC),
        .S_AXIS_BRAM_4_IS_ASYNC(S_AXIS_BRAM_4_IS_ASYNC),
        .S_AXIS_BRAM_5_IS_ASYNC(S_AXIS_BRAM_5_IS_ASYNC),
        .S_AXIS_BRAM_6_IS_ASYNC(S_AXIS_BRAM_6_IS_ASYNC),
        .S_AXIS_BRAM_7_IS_ASYNC(S_AXIS_BRAM_7_IS_ASYNC),
        .S_AXIS_BRAM_8_IS_ASYNC(S_AXIS_BRAM_8_IS_ASYNC),
        .S_AXIS_BRAM_9_IS_ASYNC(S_AXIS_BRAM_9_IS_ASYNC),
        .S_AXIS_BRAM_10_IS_ASYNC(S_AXIS_BRAM_10_IS_ASYNC),
        .S_AXIS_BRAM_11_IS_ASYNC(S_AXIS_BRAM_11_IS_ASYNC),
        .S_AXIS_BRAM_12_IS_ASYNC(S_AXIS_BRAM_12_IS_ASYNC),
        .S_AXIS_BRAM_13_IS_ASYNC(S_AXIS_BRAM_13_IS_ASYNC),
        .S_AXIS_BRAM_14_IS_ASYNC(S_AXIS_BRAM_14_IS_ASYNC),
        .S_AXIS_BRAM_15_IS_ASYNC(S_AXIS_BRAM_15_IS_ASYNC),
        .S_AXIS_BRAM_16_IS_ASYNC(S_AXIS_BRAM_16_IS_ASYNC),
        .S_AXIS_BRAM_17_IS_ASYNC(S_AXIS_BRAM_17_IS_ASYNC),
        .S_AXIS_BRAM_18_IS_ASYNC(S_AXIS_BRAM_18_IS_ASYNC),
        .S_AXIS_BRAM_19_IS_ASYNC(S_AXIS_BRAM_19_IS_ASYNC),
        .S_AXIS_BRAM_20_IS_ASYNC(S_AXIS_BRAM_20_IS_ASYNC),
        .S_AXIS_BRAM_21_IS_ASYNC(S_AXIS_BRAM_21_IS_ASYNC),
        .S_AXIS_BRAM_22_IS_ASYNC(S_AXIS_BRAM_22_IS_ASYNC),
        .S_AXIS_BRAM_23_IS_ASYNC(S_AXIS_BRAM_23_IS_ASYNC),
        .S_AXIS_BRAM_24_IS_ASYNC(S_AXIS_BRAM_24_IS_ASYNC),
        .S_AXIS_BRAM_25_IS_ASYNC(S_AXIS_BRAM_25_IS_ASYNC),
        .S_AXIS_BRAM_26_IS_ASYNC(S_AXIS_BRAM_26_IS_ASYNC),
        .S_AXIS_BRAM_27_IS_ASYNC(S_AXIS_BRAM_27_IS_ASYNC),
        .S_AXIS_BRAM_28_IS_ASYNC(S_AXIS_BRAM_28_IS_ASYNC),
        .S_AXIS_BRAM_29_IS_ASYNC(S_AXIS_BRAM_29_IS_ASYNC),
        .S_AXIS_BRAM_30_IS_ASYNC(S_AXIS_BRAM_30_IS_ASYNC),
        .S_AXIS_BRAM_31_IS_ASYNC(S_AXIS_BRAM_31_IS_ASYNC),
        .S_AXIS_BRAM_32_IS_ASYNC(S_AXIS_BRAM_32_IS_ASYNC),
        .S_AXIS_BRAM_33_IS_ASYNC(S_AXIS_BRAM_33_IS_ASYNC),
        .S_AXIS_BRAM_34_IS_ASYNC(S_AXIS_BRAM_34_IS_ASYNC),
        .S_AXIS_BRAM_35_IS_ASYNC(S_AXIS_BRAM_35_IS_ASYNC),
        .S_AXIS_BRAM_36_IS_ASYNC(S_AXIS_BRAM_36_IS_ASYNC),
        .S_AXIS_BRAM_37_IS_ASYNC(S_AXIS_BRAM_37_IS_ASYNC),
        .S_AXIS_BRAM_38_IS_ASYNC(S_AXIS_BRAM_38_IS_ASYNC),
        .S_AXIS_BRAM_39_IS_ASYNC(S_AXIS_BRAM_39_IS_ASYNC),
        .S_AXIS_BRAM_40_IS_ASYNC(S_AXIS_BRAM_40_IS_ASYNC),
        .S_AXIS_BRAM_41_IS_ASYNC(S_AXIS_BRAM_41_IS_ASYNC),
        .S_AXIS_BRAM_42_IS_ASYNC(S_AXIS_BRAM_42_IS_ASYNC),
        .S_AXIS_BRAM_43_IS_ASYNC(S_AXIS_BRAM_43_IS_ASYNC),
        .S_AXIS_BRAM_44_IS_ASYNC(S_AXIS_BRAM_44_IS_ASYNC),
        .S_AXIS_BRAM_45_IS_ASYNC(S_AXIS_BRAM_45_IS_ASYNC),
        .S_AXIS_BRAM_46_IS_ASYNC(S_AXIS_BRAM_46_IS_ASYNC),
        .S_AXIS_BRAM_47_IS_ASYNC(S_AXIS_BRAM_47_IS_ASYNC),
        .S_AXIS_BRAM_48_IS_ASYNC(S_AXIS_BRAM_48_IS_ASYNC),
        .S_AXIS_BRAM_49_IS_ASYNC(S_AXIS_BRAM_49_IS_ASYNC),
        .S_AXIS_BRAM_50_IS_ASYNC(S_AXIS_BRAM_50_IS_ASYNC),
        .S_AXIS_BRAM_51_IS_ASYNC(S_AXIS_BRAM_51_IS_ASYNC),
        .S_AXIS_BRAM_52_IS_ASYNC(S_AXIS_BRAM_52_IS_ASYNC),
        .S_AXIS_BRAM_53_IS_ASYNC(S_AXIS_BRAM_53_IS_ASYNC),
        .S_AXIS_BRAM_54_IS_ASYNC(S_AXIS_BRAM_54_IS_ASYNC),
        .S_AXIS_BRAM_55_IS_ASYNC(S_AXIS_BRAM_55_IS_ASYNC),
        .S_AXIS_BRAM_56_IS_ASYNC(S_AXIS_BRAM_56_IS_ASYNC),
        .S_AXIS_BRAM_57_IS_ASYNC(S_AXIS_BRAM_57_IS_ASYNC),
        .S_AXIS_BRAM_58_IS_ASYNC(S_AXIS_BRAM_58_IS_ASYNC),
        .S_AXIS_BRAM_59_IS_ASYNC(S_AXIS_BRAM_59_IS_ASYNC),
        .S_AXIS_BRAM_60_IS_ASYNC(S_AXIS_BRAM_60_IS_ASYNC),
        .S_AXIS_BRAM_61_IS_ASYNC(S_AXIS_BRAM_61_IS_ASYNC),
        .S_AXIS_BRAM_62_IS_ASYNC(S_AXIS_BRAM_62_IS_ASYNC),
        .S_AXIS_BRAM_63_IS_ASYNC(S_AXIS_BRAM_63_IS_ASYNC),
        .S_AXIS_BRAM_64_IS_ASYNC(S_AXIS_BRAM_64_IS_ASYNC),
        .S_AXIS_BRAM_65_IS_ASYNC(S_AXIS_BRAM_65_IS_ASYNC),
        .S_AXIS_BRAM_66_IS_ASYNC(S_AXIS_BRAM_66_IS_ASYNC),
        .S_AXIS_BRAM_67_IS_ASYNC(S_AXIS_BRAM_67_IS_ASYNC),
        .S_AXIS_BRAM_68_IS_ASYNC(S_AXIS_BRAM_68_IS_ASYNC),
        .S_AXIS_BRAM_69_IS_ASYNC(S_AXIS_BRAM_69_IS_ASYNC),
        .S_AXIS_BRAM_70_IS_ASYNC(S_AXIS_BRAM_70_IS_ASYNC),
        .S_AXIS_BRAM_71_IS_ASYNC(S_AXIS_BRAM_71_IS_ASYNC),
        .S_AXIS_BRAM_72_IS_ASYNC(S_AXIS_BRAM_72_IS_ASYNC),
        .S_AXIS_BRAM_73_IS_ASYNC(S_AXIS_BRAM_73_IS_ASYNC),
        .S_AXIS_BRAM_74_IS_ASYNC(S_AXIS_BRAM_74_IS_ASYNC),
        .S_AXIS_BRAM_75_IS_ASYNC(S_AXIS_BRAM_75_IS_ASYNC),
        .S_AXIS_BRAM_76_IS_ASYNC(S_AXIS_BRAM_76_IS_ASYNC),
        .S_AXIS_BRAM_77_IS_ASYNC(S_AXIS_BRAM_77_IS_ASYNC),
        .S_AXIS_BRAM_78_IS_ASYNC(S_AXIS_BRAM_78_IS_ASYNC),
        .S_AXIS_BRAM_79_IS_ASYNC(S_AXIS_BRAM_79_IS_ASYNC),
        .S_AXIS_BRAM_80_IS_ASYNC(S_AXIS_BRAM_80_IS_ASYNC),
        .S_AXIS_BRAM_81_IS_ASYNC(S_AXIS_BRAM_81_IS_ASYNC),
        .S_AXIS_BRAM_82_IS_ASYNC(S_AXIS_BRAM_82_IS_ASYNC),
        .S_AXIS_BRAM_83_IS_ASYNC(S_AXIS_BRAM_83_IS_ASYNC),
        .S_AXIS_BRAM_84_IS_ASYNC(S_AXIS_BRAM_84_IS_ASYNC),
        .S_AXIS_BRAM_85_IS_ASYNC(S_AXIS_BRAM_85_IS_ASYNC),
        .S_AXIS_BRAM_86_IS_ASYNC(S_AXIS_BRAM_86_IS_ASYNC),
        .S_AXIS_BRAM_87_IS_ASYNC(S_AXIS_BRAM_87_IS_ASYNC),
        .S_AXIS_BRAM_88_IS_ASYNC(S_AXIS_BRAM_88_IS_ASYNC),
        .S_AXIS_BRAM_89_IS_ASYNC(S_AXIS_BRAM_89_IS_ASYNC),
        .S_AXIS_BRAM_90_IS_ASYNC(S_AXIS_BRAM_90_IS_ASYNC),
        .S_AXIS_BRAM_91_IS_ASYNC(S_AXIS_BRAM_91_IS_ASYNC),
        .S_AXIS_BRAM_92_IS_ASYNC(S_AXIS_BRAM_92_IS_ASYNC),
        .S_AXIS_BRAM_93_IS_ASYNC(S_AXIS_BRAM_93_IS_ASYNC),
        .S_AXIS_BRAM_94_IS_ASYNC(S_AXIS_BRAM_94_IS_ASYNC),
        .S_AXIS_BRAM_95_IS_ASYNC(S_AXIS_BRAM_95_IS_ASYNC),
        .S_AXIS_BRAM_96_IS_ASYNC(S_AXIS_BRAM_96_IS_ASYNC),
        .S_AXIS_BRAM_97_IS_ASYNC(S_AXIS_BRAM_97_IS_ASYNC),
        .S_AXIS_BRAM_98_IS_ASYNC(S_AXIS_BRAM_98_IS_ASYNC),
        .S_AXIS_BRAM_99_IS_ASYNC(S_AXIS_BRAM_99_IS_ASYNC),
        .S_AXIS_BRAM_100_IS_ASYNC(S_AXIS_BRAM_100_IS_ASYNC),
        .S_AXIS_BRAM_101_IS_ASYNC(S_AXIS_BRAM_101_IS_ASYNC),
        .S_AXIS_BRAM_102_IS_ASYNC(S_AXIS_BRAM_102_IS_ASYNC),
        .S_AXIS_BRAM_103_IS_ASYNC(S_AXIS_BRAM_103_IS_ASYNC),
        .S_AXIS_BRAM_104_IS_ASYNC(S_AXIS_BRAM_104_IS_ASYNC),
        .S_AXIS_BRAM_105_IS_ASYNC(S_AXIS_BRAM_105_IS_ASYNC),
        .S_AXIS_BRAM_106_IS_ASYNC(S_AXIS_BRAM_106_IS_ASYNC),
        .S_AXIS_BRAM_107_IS_ASYNC(S_AXIS_BRAM_107_IS_ASYNC),
        .S_AXIS_BRAM_108_IS_ASYNC(S_AXIS_BRAM_108_IS_ASYNC),
        .S_AXIS_BRAM_109_IS_ASYNC(S_AXIS_BRAM_109_IS_ASYNC),
        .S_AXIS_BRAM_110_IS_ASYNC(S_AXIS_BRAM_110_IS_ASYNC),
        .S_AXIS_BRAM_111_IS_ASYNC(S_AXIS_BRAM_111_IS_ASYNC),
        .S_AXIS_BRAM_112_IS_ASYNC(S_AXIS_BRAM_112_IS_ASYNC),
        .S_AXIS_BRAM_113_IS_ASYNC(S_AXIS_BRAM_113_IS_ASYNC),
        .S_AXIS_BRAM_114_IS_ASYNC(S_AXIS_BRAM_114_IS_ASYNC),
        .S_AXIS_BRAM_115_IS_ASYNC(S_AXIS_BRAM_115_IS_ASYNC),
        .S_AXIS_BRAM_116_IS_ASYNC(S_AXIS_BRAM_116_IS_ASYNC),
        .S_AXIS_BRAM_117_IS_ASYNC(S_AXIS_BRAM_117_IS_ASYNC),
        .S_AXIS_BRAM_118_IS_ASYNC(S_AXIS_BRAM_118_IS_ASYNC),
        .S_AXIS_BRAM_119_IS_ASYNC(S_AXIS_BRAM_119_IS_ASYNC),
        .S_AXIS_BRAM_120_IS_ASYNC(S_AXIS_BRAM_120_IS_ASYNC),
        .S_AXIS_BRAM_121_IS_ASYNC(S_AXIS_BRAM_121_IS_ASYNC),
        .S_AXIS_BRAM_122_IS_ASYNC(S_AXIS_BRAM_122_IS_ASYNC),
        .S_AXIS_BRAM_123_IS_ASYNC(S_AXIS_BRAM_123_IS_ASYNC),
        .S_AXIS_BRAM_124_IS_ASYNC(S_AXIS_BRAM_124_IS_ASYNC),
        .S_AXIS_BRAM_125_IS_ASYNC(S_AXIS_BRAM_125_IS_ASYNC),
        .S_AXIS_BRAM_126_IS_ASYNC(S_AXIS_BRAM_126_IS_ASYNC),
        .S_AXIS_BRAM_127_IS_ASYNC(S_AXIS_BRAM_127_IS_ASYNC),
        .M_AXIS_BRAMIO_0_IS_ASYNC(M_AXIS_BRAMIO_0_IS_ASYNC),
        .M_AXIS_BRAMIO_1_IS_ASYNC(M_AXIS_BRAMIO_1_IS_ASYNC),
        .M_AXIS_BRAMIO_2_IS_ASYNC(M_AXIS_BRAMIO_2_IS_ASYNC),
        .M_AXIS_BRAMIO_3_IS_ASYNC(M_AXIS_BRAMIO_3_IS_ASYNC),
        .M_AXIS_BRAMIO_4_IS_ASYNC(M_AXIS_BRAMIO_4_IS_ASYNC),
        .M_AXIS_BRAMIO_5_IS_ASYNC(M_AXIS_BRAMIO_5_IS_ASYNC),
        .M_AXIS_BRAMIO_6_IS_ASYNC(M_AXIS_BRAMIO_6_IS_ASYNC),
        .M_AXIS_BRAMIO_7_IS_ASYNC(M_AXIS_BRAMIO_7_IS_ASYNC),
        .M_AXIS_BRAMIO_8_IS_ASYNC(M_AXIS_BRAMIO_8_IS_ASYNC),
        .M_AXIS_BRAMIO_9_IS_ASYNC(M_AXIS_BRAMIO_9_IS_ASYNC),
        .M_AXIS_BRAMIO_10_IS_ASYNC(M_AXIS_BRAMIO_10_IS_ASYNC),
        .M_AXIS_BRAMIO_11_IS_ASYNC(M_AXIS_BRAMIO_11_IS_ASYNC),
        .M_AXIS_BRAMIO_12_IS_ASYNC(M_AXIS_BRAMIO_12_IS_ASYNC),
        .M_AXIS_BRAMIO_13_IS_ASYNC(M_AXIS_BRAMIO_13_IS_ASYNC),
        .M_AXIS_BRAMIO_14_IS_ASYNC(M_AXIS_BRAMIO_14_IS_ASYNC),
        .M_AXIS_BRAMIO_15_IS_ASYNC(M_AXIS_BRAMIO_15_IS_ASYNC),
        .M_AXIS_BRAMIO_16_IS_ASYNC(M_AXIS_BRAMIO_16_IS_ASYNC),
        .M_AXIS_BRAMIO_17_IS_ASYNC(M_AXIS_BRAMIO_17_IS_ASYNC),
        .M_AXIS_BRAMIO_18_IS_ASYNC(M_AXIS_BRAMIO_18_IS_ASYNC),
        .M_AXIS_BRAMIO_19_IS_ASYNC(M_AXIS_BRAMIO_19_IS_ASYNC),
        .M_AXIS_BRAMIO_20_IS_ASYNC(M_AXIS_BRAMIO_20_IS_ASYNC),
        .M_AXIS_BRAMIO_21_IS_ASYNC(M_AXIS_BRAMIO_21_IS_ASYNC),
        .M_AXIS_BRAMIO_22_IS_ASYNC(M_AXIS_BRAMIO_22_IS_ASYNC),
        .M_AXIS_BRAMIO_23_IS_ASYNC(M_AXIS_BRAMIO_23_IS_ASYNC),
        .M_AXIS_BRAMIO_24_IS_ASYNC(M_AXIS_BRAMIO_24_IS_ASYNC),
        .M_AXIS_BRAMIO_25_IS_ASYNC(M_AXIS_BRAMIO_25_IS_ASYNC),
        .M_AXIS_BRAMIO_26_IS_ASYNC(M_AXIS_BRAMIO_26_IS_ASYNC),
        .M_AXIS_BRAMIO_27_IS_ASYNC(M_AXIS_BRAMIO_27_IS_ASYNC),
        .M_AXIS_BRAMIO_28_IS_ASYNC(M_AXIS_BRAMIO_28_IS_ASYNC),
        .M_AXIS_BRAMIO_29_IS_ASYNC(M_AXIS_BRAMIO_29_IS_ASYNC),
        .M_AXIS_BRAMIO_30_IS_ASYNC(M_AXIS_BRAMIO_30_IS_ASYNC),
        .M_AXIS_BRAMIO_31_IS_ASYNC(M_AXIS_BRAMIO_31_IS_ASYNC),
        .M_AXIS_BRAMIO_32_IS_ASYNC(M_AXIS_BRAMIO_32_IS_ASYNC),
        .M_AXIS_BRAMIO_33_IS_ASYNC(M_AXIS_BRAMIO_33_IS_ASYNC),
        .M_AXIS_BRAMIO_34_IS_ASYNC(M_AXIS_BRAMIO_34_IS_ASYNC),
        .M_AXIS_BRAMIO_35_IS_ASYNC(M_AXIS_BRAMIO_35_IS_ASYNC),
        .M_AXIS_BRAMIO_36_IS_ASYNC(M_AXIS_BRAMIO_36_IS_ASYNC),
        .M_AXIS_BRAMIO_37_IS_ASYNC(M_AXIS_BRAMIO_37_IS_ASYNC),
        .M_AXIS_BRAMIO_38_IS_ASYNC(M_AXIS_BRAMIO_38_IS_ASYNC),
        .M_AXIS_BRAMIO_39_IS_ASYNC(M_AXIS_BRAMIO_39_IS_ASYNC),
        .M_AXIS_BRAMIO_40_IS_ASYNC(M_AXIS_BRAMIO_40_IS_ASYNC),
        .M_AXIS_BRAMIO_41_IS_ASYNC(M_AXIS_BRAMIO_41_IS_ASYNC),
        .M_AXIS_BRAMIO_42_IS_ASYNC(M_AXIS_BRAMIO_42_IS_ASYNC),
        .M_AXIS_BRAMIO_43_IS_ASYNC(M_AXIS_BRAMIO_43_IS_ASYNC),
        .M_AXIS_BRAMIO_44_IS_ASYNC(M_AXIS_BRAMIO_44_IS_ASYNC),
        .M_AXIS_BRAMIO_45_IS_ASYNC(M_AXIS_BRAMIO_45_IS_ASYNC),
        .M_AXIS_BRAMIO_46_IS_ASYNC(M_AXIS_BRAMIO_46_IS_ASYNC),
        .M_AXIS_BRAMIO_47_IS_ASYNC(M_AXIS_BRAMIO_47_IS_ASYNC),
        .M_AXIS_BRAMIO_48_IS_ASYNC(M_AXIS_BRAMIO_48_IS_ASYNC),
        .M_AXIS_BRAMIO_49_IS_ASYNC(M_AXIS_BRAMIO_49_IS_ASYNC),
        .M_AXIS_BRAMIO_50_IS_ASYNC(M_AXIS_BRAMIO_50_IS_ASYNC),
        .M_AXIS_BRAMIO_51_IS_ASYNC(M_AXIS_BRAMIO_51_IS_ASYNC),
        .M_AXIS_BRAMIO_52_IS_ASYNC(M_AXIS_BRAMIO_52_IS_ASYNC),
        .M_AXIS_BRAMIO_53_IS_ASYNC(M_AXIS_BRAMIO_53_IS_ASYNC),
        .M_AXIS_BRAMIO_54_IS_ASYNC(M_AXIS_BRAMIO_54_IS_ASYNC),
        .M_AXIS_BRAMIO_55_IS_ASYNC(M_AXIS_BRAMIO_55_IS_ASYNC),
        .M_AXIS_BRAMIO_56_IS_ASYNC(M_AXIS_BRAMIO_56_IS_ASYNC),
        .M_AXIS_BRAMIO_57_IS_ASYNC(M_AXIS_BRAMIO_57_IS_ASYNC),
        .M_AXIS_BRAMIO_58_IS_ASYNC(M_AXIS_BRAMIO_58_IS_ASYNC),
        .M_AXIS_BRAMIO_59_IS_ASYNC(M_AXIS_BRAMIO_59_IS_ASYNC),
        .M_AXIS_BRAMIO_60_IS_ASYNC(M_AXIS_BRAMIO_60_IS_ASYNC),
        .M_AXIS_BRAMIO_61_IS_ASYNC(M_AXIS_BRAMIO_61_IS_ASYNC),
        .M_AXIS_BRAMIO_62_IS_ASYNC(M_AXIS_BRAMIO_62_IS_ASYNC),
        .M_AXIS_BRAMIO_63_IS_ASYNC(M_AXIS_BRAMIO_63_IS_ASYNC),
        .M_AXIS_BRAMIO_64_IS_ASYNC(M_AXIS_BRAMIO_64_IS_ASYNC),
        .M_AXIS_BRAMIO_65_IS_ASYNC(M_AXIS_BRAMIO_65_IS_ASYNC),
        .M_AXIS_BRAMIO_66_IS_ASYNC(M_AXIS_BRAMIO_66_IS_ASYNC),
        .M_AXIS_BRAMIO_67_IS_ASYNC(M_AXIS_BRAMIO_67_IS_ASYNC),
        .M_AXIS_BRAMIO_68_IS_ASYNC(M_AXIS_BRAMIO_68_IS_ASYNC),
        .M_AXIS_BRAMIO_69_IS_ASYNC(M_AXIS_BRAMIO_69_IS_ASYNC),
        .M_AXIS_BRAMIO_70_IS_ASYNC(M_AXIS_BRAMIO_70_IS_ASYNC),
        .M_AXIS_BRAMIO_71_IS_ASYNC(M_AXIS_BRAMIO_71_IS_ASYNC),
        .M_AXIS_BRAMIO_72_IS_ASYNC(M_AXIS_BRAMIO_72_IS_ASYNC),
        .M_AXIS_BRAMIO_73_IS_ASYNC(M_AXIS_BRAMIO_73_IS_ASYNC),
        .M_AXIS_BRAMIO_74_IS_ASYNC(M_AXIS_BRAMIO_74_IS_ASYNC),
        .M_AXIS_BRAMIO_75_IS_ASYNC(M_AXIS_BRAMIO_75_IS_ASYNC),
        .M_AXIS_BRAMIO_76_IS_ASYNC(M_AXIS_BRAMIO_76_IS_ASYNC),
        .M_AXIS_BRAMIO_77_IS_ASYNC(M_AXIS_BRAMIO_77_IS_ASYNC),
        .M_AXIS_BRAMIO_78_IS_ASYNC(M_AXIS_BRAMIO_78_IS_ASYNC),
        .M_AXIS_BRAMIO_79_IS_ASYNC(M_AXIS_BRAMIO_79_IS_ASYNC),
        .M_AXIS_BRAMIO_80_IS_ASYNC(M_AXIS_BRAMIO_80_IS_ASYNC),
        .M_AXIS_BRAMIO_81_IS_ASYNC(M_AXIS_BRAMIO_81_IS_ASYNC),
        .M_AXIS_BRAMIO_82_IS_ASYNC(M_AXIS_BRAMIO_82_IS_ASYNC),
        .M_AXIS_BRAMIO_83_IS_ASYNC(M_AXIS_BRAMIO_83_IS_ASYNC),
        .M_AXIS_BRAMIO_84_IS_ASYNC(M_AXIS_BRAMIO_84_IS_ASYNC),
        .M_AXIS_BRAMIO_85_IS_ASYNC(M_AXIS_BRAMIO_85_IS_ASYNC),
        .M_AXIS_BRAMIO_86_IS_ASYNC(M_AXIS_BRAMIO_86_IS_ASYNC),
        .M_AXIS_BRAMIO_87_IS_ASYNC(M_AXIS_BRAMIO_87_IS_ASYNC),
        .M_AXIS_BRAMIO_88_IS_ASYNC(M_AXIS_BRAMIO_88_IS_ASYNC),
        .M_AXIS_BRAMIO_89_IS_ASYNC(M_AXIS_BRAMIO_89_IS_ASYNC),
        .M_AXIS_BRAMIO_90_IS_ASYNC(M_AXIS_BRAMIO_90_IS_ASYNC),
        .M_AXIS_BRAMIO_91_IS_ASYNC(M_AXIS_BRAMIO_91_IS_ASYNC),
        .M_AXIS_BRAMIO_92_IS_ASYNC(M_AXIS_BRAMIO_92_IS_ASYNC),
        .M_AXIS_BRAMIO_93_IS_ASYNC(M_AXIS_BRAMIO_93_IS_ASYNC),
        .M_AXIS_BRAMIO_94_IS_ASYNC(M_AXIS_BRAMIO_94_IS_ASYNC),
        .M_AXIS_BRAMIO_95_IS_ASYNC(M_AXIS_BRAMIO_95_IS_ASYNC),
        .M_AXIS_BRAMIO_96_IS_ASYNC(M_AXIS_BRAMIO_96_IS_ASYNC),
        .M_AXIS_BRAMIO_97_IS_ASYNC(M_AXIS_BRAMIO_97_IS_ASYNC),
        .M_AXIS_BRAMIO_98_IS_ASYNC(M_AXIS_BRAMIO_98_IS_ASYNC),
        .M_AXIS_BRAMIO_99_IS_ASYNC(M_AXIS_BRAMIO_99_IS_ASYNC),
        .M_AXIS_BRAMIO_100_IS_ASYNC(M_AXIS_BRAMIO_100_IS_ASYNC),
        .M_AXIS_BRAMIO_101_IS_ASYNC(M_AXIS_BRAMIO_101_IS_ASYNC),
        .M_AXIS_BRAMIO_102_IS_ASYNC(M_AXIS_BRAMIO_102_IS_ASYNC),
        .M_AXIS_BRAMIO_103_IS_ASYNC(M_AXIS_BRAMIO_103_IS_ASYNC),
        .M_AXIS_BRAMIO_104_IS_ASYNC(M_AXIS_BRAMIO_104_IS_ASYNC),
        .M_AXIS_BRAMIO_105_IS_ASYNC(M_AXIS_BRAMIO_105_IS_ASYNC),
        .M_AXIS_BRAMIO_106_IS_ASYNC(M_AXIS_BRAMIO_106_IS_ASYNC),
        .M_AXIS_BRAMIO_107_IS_ASYNC(M_AXIS_BRAMIO_107_IS_ASYNC),
        .M_AXIS_BRAMIO_108_IS_ASYNC(M_AXIS_BRAMIO_108_IS_ASYNC),
        .M_AXIS_BRAMIO_109_IS_ASYNC(M_AXIS_BRAMIO_109_IS_ASYNC),
        .M_AXIS_BRAMIO_110_IS_ASYNC(M_AXIS_BRAMIO_110_IS_ASYNC),
        .M_AXIS_BRAMIO_111_IS_ASYNC(M_AXIS_BRAMIO_111_IS_ASYNC),
        .M_AXIS_BRAMIO_112_IS_ASYNC(M_AXIS_BRAMIO_112_IS_ASYNC),
        .M_AXIS_BRAMIO_113_IS_ASYNC(M_AXIS_BRAMIO_113_IS_ASYNC),
        .M_AXIS_BRAMIO_114_IS_ASYNC(M_AXIS_BRAMIO_114_IS_ASYNC),
        .M_AXIS_BRAMIO_115_IS_ASYNC(M_AXIS_BRAMIO_115_IS_ASYNC),
        .M_AXIS_BRAMIO_116_IS_ASYNC(M_AXIS_BRAMIO_116_IS_ASYNC),
        .M_AXIS_BRAMIO_117_IS_ASYNC(M_AXIS_BRAMIO_117_IS_ASYNC),
        .M_AXIS_BRAMIO_118_IS_ASYNC(M_AXIS_BRAMIO_118_IS_ASYNC),
        .M_AXIS_BRAMIO_119_IS_ASYNC(M_AXIS_BRAMIO_119_IS_ASYNC),
        .M_AXIS_BRAMIO_120_IS_ASYNC(M_AXIS_BRAMIO_120_IS_ASYNC),
        .M_AXIS_BRAMIO_121_IS_ASYNC(M_AXIS_BRAMIO_121_IS_ASYNC),
        .M_AXIS_BRAMIO_122_IS_ASYNC(M_AXIS_BRAMIO_122_IS_ASYNC),
        .M_AXIS_BRAMIO_123_IS_ASYNC(M_AXIS_BRAMIO_123_IS_ASYNC),
        .M_AXIS_BRAMIO_124_IS_ASYNC(M_AXIS_BRAMIO_124_IS_ASYNC),
        .M_AXIS_BRAMIO_125_IS_ASYNC(M_AXIS_BRAMIO_125_IS_ASYNC),
        .M_AXIS_BRAMIO_126_IS_ASYNC(M_AXIS_BRAMIO_126_IS_ASYNC),
        .M_AXIS_BRAMIO_127_IS_ASYNC(M_AXIS_BRAMIO_127_IS_ASYNC),
        .S_AXIS_BRAM_0_IS_INOUT(S_AXIS_BRAM_0_IS_INOUT),
        .S_AXIS_BRAM_1_IS_INOUT(S_AXIS_BRAM_1_IS_INOUT),
        .S_AXIS_BRAM_2_IS_INOUT(S_AXIS_BRAM_2_IS_INOUT),
        .S_AXIS_BRAM_3_IS_INOUT(S_AXIS_BRAM_3_IS_INOUT),
        .S_AXIS_BRAM_4_IS_INOUT(S_AXIS_BRAM_4_IS_INOUT),
        .S_AXIS_BRAM_5_IS_INOUT(S_AXIS_BRAM_5_IS_INOUT),
        .S_AXIS_BRAM_6_IS_INOUT(S_AXIS_BRAM_6_IS_INOUT),
        .S_AXIS_BRAM_7_IS_INOUT(S_AXIS_BRAM_7_IS_INOUT),
        .S_AXIS_BRAM_8_IS_INOUT(S_AXIS_BRAM_8_IS_INOUT),
        .S_AXIS_BRAM_9_IS_INOUT(S_AXIS_BRAM_9_IS_INOUT),
        .S_AXIS_BRAM_10_IS_INOUT(S_AXIS_BRAM_10_IS_INOUT),
        .S_AXIS_BRAM_11_IS_INOUT(S_AXIS_BRAM_11_IS_INOUT),
        .S_AXIS_BRAM_12_IS_INOUT(S_AXIS_BRAM_12_IS_INOUT),
        .S_AXIS_BRAM_13_IS_INOUT(S_AXIS_BRAM_13_IS_INOUT),
        .S_AXIS_BRAM_14_IS_INOUT(S_AXIS_BRAM_14_IS_INOUT),
        .S_AXIS_BRAM_15_IS_INOUT(S_AXIS_BRAM_15_IS_INOUT),
        .S_AXIS_BRAM_16_IS_INOUT(S_AXIS_BRAM_16_IS_INOUT),
        .S_AXIS_BRAM_17_IS_INOUT(S_AXIS_BRAM_17_IS_INOUT),
        .S_AXIS_BRAM_18_IS_INOUT(S_AXIS_BRAM_18_IS_INOUT),
        .S_AXIS_BRAM_19_IS_INOUT(S_AXIS_BRAM_19_IS_INOUT),
        .S_AXIS_BRAM_20_IS_INOUT(S_AXIS_BRAM_20_IS_INOUT),
        .S_AXIS_BRAM_21_IS_INOUT(S_AXIS_BRAM_21_IS_INOUT),
        .S_AXIS_BRAM_22_IS_INOUT(S_AXIS_BRAM_22_IS_INOUT),
        .S_AXIS_BRAM_23_IS_INOUT(S_AXIS_BRAM_23_IS_INOUT),
        .S_AXIS_BRAM_24_IS_INOUT(S_AXIS_BRAM_24_IS_INOUT),
        .S_AXIS_BRAM_25_IS_INOUT(S_AXIS_BRAM_25_IS_INOUT),
        .S_AXIS_BRAM_26_IS_INOUT(S_AXIS_BRAM_26_IS_INOUT),
        .S_AXIS_BRAM_27_IS_INOUT(S_AXIS_BRAM_27_IS_INOUT),
        .S_AXIS_BRAM_28_IS_INOUT(S_AXIS_BRAM_28_IS_INOUT),
        .S_AXIS_BRAM_29_IS_INOUT(S_AXIS_BRAM_29_IS_INOUT),
        .S_AXIS_BRAM_30_IS_INOUT(S_AXIS_BRAM_30_IS_INOUT),
        .S_AXIS_BRAM_31_IS_INOUT(S_AXIS_BRAM_31_IS_INOUT),
        .S_AXIS_BRAM_32_IS_INOUT(S_AXIS_BRAM_32_IS_INOUT),
        .S_AXIS_BRAM_33_IS_INOUT(S_AXIS_BRAM_33_IS_INOUT),
        .S_AXIS_BRAM_34_IS_INOUT(S_AXIS_BRAM_34_IS_INOUT),
        .S_AXIS_BRAM_35_IS_INOUT(S_AXIS_BRAM_35_IS_INOUT),
        .S_AXIS_BRAM_36_IS_INOUT(S_AXIS_BRAM_36_IS_INOUT),
        .S_AXIS_BRAM_37_IS_INOUT(S_AXIS_BRAM_37_IS_INOUT),
        .S_AXIS_BRAM_38_IS_INOUT(S_AXIS_BRAM_38_IS_INOUT),
        .S_AXIS_BRAM_39_IS_INOUT(S_AXIS_BRAM_39_IS_INOUT),
        .S_AXIS_BRAM_40_IS_INOUT(S_AXIS_BRAM_40_IS_INOUT),
        .S_AXIS_BRAM_41_IS_INOUT(S_AXIS_BRAM_41_IS_INOUT),
        .S_AXIS_BRAM_42_IS_INOUT(S_AXIS_BRAM_42_IS_INOUT),
        .S_AXIS_BRAM_43_IS_INOUT(S_AXIS_BRAM_43_IS_INOUT),
        .S_AXIS_BRAM_44_IS_INOUT(S_AXIS_BRAM_44_IS_INOUT),
        .S_AXIS_BRAM_45_IS_INOUT(S_AXIS_BRAM_45_IS_INOUT),
        .S_AXIS_BRAM_46_IS_INOUT(S_AXIS_BRAM_46_IS_INOUT),
        .S_AXIS_BRAM_47_IS_INOUT(S_AXIS_BRAM_47_IS_INOUT),
        .S_AXIS_BRAM_48_IS_INOUT(S_AXIS_BRAM_48_IS_INOUT),
        .S_AXIS_BRAM_49_IS_INOUT(S_AXIS_BRAM_49_IS_INOUT),
        .S_AXIS_BRAM_50_IS_INOUT(S_AXIS_BRAM_50_IS_INOUT),
        .S_AXIS_BRAM_51_IS_INOUT(S_AXIS_BRAM_51_IS_INOUT),
        .S_AXIS_BRAM_52_IS_INOUT(S_AXIS_BRAM_52_IS_INOUT),
        .S_AXIS_BRAM_53_IS_INOUT(S_AXIS_BRAM_53_IS_INOUT),
        .S_AXIS_BRAM_54_IS_INOUT(S_AXIS_BRAM_54_IS_INOUT),
        .S_AXIS_BRAM_55_IS_INOUT(S_AXIS_BRAM_55_IS_INOUT),
        .S_AXIS_BRAM_56_IS_INOUT(S_AXIS_BRAM_56_IS_INOUT),
        .S_AXIS_BRAM_57_IS_INOUT(S_AXIS_BRAM_57_IS_INOUT),
        .S_AXIS_BRAM_58_IS_INOUT(S_AXIS_BRAM_58_IS_INOUT),
        .S_AXIS_BRAM_59_IS_INOUT(S_AXIS_BRAM_59_IS_INOUT),
        .S_AXIS_BRAM_60_IS_INOUT(S_AXIS_BRAM_60_IS_INOUT),
        .S_AXIS_BRAM_61_IS_INOUT(S_AXIS_BRAM_61_IS_INOUT),
        .S_AXIS_BRAM_62_IS_INOUT(S_AXIS_BRAM_62_IS_INOUT),
        .S_AXIS_BRAM_63_IS_INOUT(S_AXIS_BRAM_63_IS_INOUT),
        .S_AXIS_BRAM_64_IS_INOUT(S_AXIS_BRAM_64_IS_INOUT),
        .S_AXIS_BRAM_65_IS_INOUT(S_AXIS_BRAM_65_IS_INOUT),
        .S_AXIS_BRAM_66_IS_INOUT(S_AXIS_BRAM_66_IS_INOUT),
        .S_AXIS_BRAM_67_IS_INOUT(S_AXIS_BRAM_67_IS_INOUT),
        .S_AXIS_BRAM_68_IS_INOUT(S_AXIS_BRAM_68_IS_INOUT),
        .S_AXIS_BRAM_69_IS_INOUT(S_AXIS_BRAM_69_IS_INOUT),
        .S_AXIS_BRAM_70_IS_INOUT(S_AXIS_BRAM_70_IS_INOUT),
        .S_AXIS_BRAM_71_IS_INOUT(S_AXIS_BRAM_71_IS_INOUT),
        .S_AXIS_BRAM_72_IS_INOUT(S_AXIS_BRAM_72_IS_INOUT),
        .S_AXIS_BRAM_73_IS_INOUT(S_AXIS_BRAM_73_IS_INOUT),
        .S_AXIS_BRAM_74_IS_INOUT(S_AXIS_BRAM_74_IS_INOUT),
        .S_AXIS_BRAM_75_IS_INOUT(S_AXIS_BRAM_75_IS_INOUT),
        .S_AXIS_BRAM_76_IS_INOUT(S_AXIS_BRAM_76_IS_INOUT),
        .S_AXIS_BRAM_77_IS_INOUT(S_AXIS_BRAM_77_IS_INOUT),
        .S_AXIS_BRAM_78_IS_INOUT(S_AXIS_BRAM_78_IS_INOUT),
        .S_AXIS_BRAM_79_IS_INOUT(S_AXIS_BRAM_79_IS_INOUT),
        .S_AXIS_BRAM_80_IS_INOUT(S_AXIS_BRAM_80_IS_INOUT),
        .S_AXIS_BRAM_81_IS_INOUT(S_AXIS_BRAM_81_IS_INOUT),
        .S_AXIS_BRAM_82_IS_INOUT(S_AXIS_BRAM_82_IS_INOUT),
        .S_AXIS_BRAM_83_IS_INOUT(S_AXIS_BRAM_83_IS_INOUT),
        .S_AXIS_BRAM_84_IS_INOUT(S_AXIS_BRAM_84_IS_INOUT),
        .S_AXIS_BRAM_85_IS_INOUT(S_AXIS_BRAM_85_IS_INOUT),
        .S_AXIS_BRAM_86_IS_INOUT(S_AXIS_BRAM_86_IS_INOUT),
        .S_AXIS_BRAM_87_IS_INOUT(S_AXIS_BRAM_87_IS_INOUT),
        .S_AXIS_BRAM_88_IS_INOUT(S_AXIS_BRAM_88_IS_INOUT),
        .S_AXIS_BRAM_89_IS_INOUT(S_AXIS_BRAM_89_IS_INOUT),
        .S_AXIS_BRAM_90_IS_INOUT(S_AXIS_BRAM_90_IS_INOUT),
        .S_AXIS_BRAM_91_IS_INOUT(S_AXIS_BRAM_91_IS_INOUT),
        .S_AXIS_BRAM_92_IS_INOUT(S_AXIS_BRAM_92_IS_INOUT),
        .S_AXIS_BRAM_93_IS_INOUT(S_AXIS_BRAM_93_IS_INOUT),
        .S_AXIS_BRAM_94_IS_INOUT(S_AXIS_BRAM_94_IS_INOUT),
        .S_AXIS_BRAM_95_IS_INOUT(S_AXIS_BRAM_95_IS_INOUT),
        .S_AXIS_BRAM_96_IS_INOUT(S_AXIS_BRAM_96_IS_INOUT),
        .S_AXIS_BRAM_97_IS_INOUT(S_AXIS_BRAM_97_IS_INOUT),
        .S_AXIS_BRAM_98_IS_INOUT(S_AXIS_BRAM_98_IS_INOUT),
        .S_AXIS_BRAM_99_IS_INOUT(S_AXIS_BRAM_99_IS_INOUT),
        .S_AXIS_BRAM_100_IS_INOUT(S_AXIS_BRAM_100_IS_INOUT),
        .S_AXIS_BRAM_101_IS_INOUT(S_AXIS_BRAM_101_IS_INOUT),
        .S_AXIS_BRAM_102_IS_INOUT(S_AXIS_BRAM_102_IS_INOUT),
        .S_AXIS_BRAM_103_IS_INOUT(S_AXIS_BRAM_103_IS_INOUT),
        .S_AXIS_BRAM_104_IS_INOUT(S_AXIS_BRAM_104_IS_INOUT),
        .S_AXIS_BRAM_105_IS_INOUT(S_AXIS_BRAM_105_IS_INOUT),
        .S_AXIS_BRAM_106_IS_INOUT(S_AXIS_BRAM_106_IS_INOUT),
        .S_AXIS_BRAM_107_IS_INOUT(S_AXIS_BRAM_107_IS_INOUT),
        .S_AXIS_BRAM_108_IS_INOUT(S_AXIS_BRAM_108_IS_INOUT),
        .S_AXIS_BRAM_109_IS_INOUT(S_AXIS_BRAM_109_IS_INOUT),
        .S_AXIS_BRAM_110_IS_INOUT(S_AXIS_BRAM_110_IS_INOUT),
        .S_AXIS_BRAM_111_IS_INOUT(S_AXIS_BRAM_111_IS_INOUT),
        .S_AXIS_BRAM_112_IS_INOUT(S_AXIS_BRAM_112_IS_INOUT),
        .S_AXIS_BRAM_113_IS_INOUT(S_AXIS_BRAM_113_IS_INOUT),
        .S_AXIS_BRAM_114_IS_INOUT(S_AXIS_BRAM_114_IS_INOUT),
        .S_AXIS_BRAM_115_IS_INOUT(S_AXIS_BRAM_115_IS_INOUT),
        .S_AXIS_BRAM_116_IS_INOUT(S_AXIS_BRAM_116_IS_INOUT),
        .S_AXIS_BRAM_117_IS_INOUT(S_AXIS_BRAM_117_IS_INOUT),
        .S_AXIS_BRAM_118_IS_INOUT(S_AXIS_BRAM_118_IS_INOUT),
        .S_AXIS_BRAM_119_IS_INOUT(S_AXIS_BRAM_119_IS_INOUT),
        .S_AXIS_BRAM_120_IS_INOUT(S_AXIS_BRAM_120_IS_INOUT),
        .S_AXIS_BRAM_121_IS_INOUT(S_AXIS_BRAM_121_IS_INOUT),
        .S_AXIS_BRAM_122_IS_INOUT(S_AXIS_BRAM_122_IS_INOUT),
        .S_AXIS_BRAM_123_IS_INOUT(S_AXIS_BRAM_123_IS_INOUT),
        .S_AXIS_BRAM_124_IS_INOUT(S_AXIS_BRAM_124_IS_INOUT),
        .S_AXIS_BRAM_125_IS_INOUT(S_AXIS_BRAM_125_IS_INOUT),
        .S_AXIS_BRAM_126_IS_INOUT(S_AXIS_BRAM_126_IS_INOUT),
        .S_AXIS_BRAM_127_IS_INOUT(S_AXIS_BRAM_127_IS_INOUT),
        .S_AXIS_BRAM_0_MB_DEPTH(S_AXIS_BRAM_0_MB_DEPTH),
        .S_AXIS_BRAM_1_MB_DEPTH(S_AXIS_BRAM_1_MB_DEPTH),
        .S_AXIS_BRAM_2_MB_DEPTH(S_AXIS_BRAM_2_MB_DEPTH),
        .S_AXIS_BRAM_3_MB_DEPTH(S_AXIS_BRAM_3_MB_DEPTH),
        .S_AXIS_BRAM_4_MB_DEPTH(S_AXIS_BRAM_4_MB_DEPTH),
        .S_AXIS_BRAM_5_MB_DEPTH(S_AXIS_BRAM_5_MB_DEPTH),
        .S_AXIS_BRAM_6_MB_DEPTH(S_AXIS_BRAM_6_MB_DEPTH),
        .S_AXIS_BRAM_7_MB_DEPTH(S_AXIS_BRAM_7_MB_DEPTH),
        .S_AXIS_BRAM_8_MB_DEPTH(S_AXIS_BRAM_8_MB_DEPTH),
        .S_AXIS_BRAM_9_MB_DEPTH(S_AXIS_BRAM_9_MB_DEPTH),
        .S_AXIS_BRAM_10_MB_DEPTH(S_AXIS_BRAM_10_MB_DEPTH),
        .S_AXIS_BRAM_11_MB_DEPTH(S_AXIS_BRAM_11_MB_DEPTH),
        .S_AXIS_BRAM_12_MB_DEPTH(S_AXIS_BRAM_12_MB_DEPTH),
        .S_AXIS_BRAM_13_MB_DEPTH(S_AXIS_BRAM_13_MB_DEPTH),
        .S_AXIS_BRAM_14_MB_DEPTH(S_AXIS_BRAM_14_MB_DEPTH),
        .S_AXIS_BRAM_15_MB_DEPTH(S_AXIS_BRAM_15_MB_DEPTH),
        .S_AXIS_BRAM_16_MB_DEPTH(S_AXIS_BRAM_16_MB_DEPTH),
        .S_AXIS_BRAM_17_MB_DEPTH(S_AXIS_BRAM_17_MB_DEPTH),
        .S_AXIS_BRAM_18_MB_DEPTH(S_AXIS_BRAM_18_MB_DEPTH),
        .S_AXIS_BRAM_19_MB_DEPTH(S_AXIS_BRAM_19_MB_DEPTH),
        .S_AXIS_BRAM_20_MB_DEPTH(S_AXIS_BRAM_20_MB_DEPTH),
        .S_AXIS_BRAM_21_MB_DEPTH(S_AXIS_BRAM_21_MB_DEPTH),
        .S_AXIS_BRAM_22_MB_DEPTH(S_AXIS_BRAM_22_MB_DEPTH),
        .S_AXIS_BRAM_23_MB_DEPTH(S_AXIS_BRAM_23_MB_DEPTH),
        .S_AXIS_BRAM_24_MB_DEPTH(S_AXIS_BRAM_24_MB_DEPTH),
        .S_AXIS_BRAM_25_MB_DEPTH(S_AXIS_BRAM_25_MB_DEPTH),
        .S_AXIS_BRAM_26_MB_DEPTH(S_AXIS_BRAM_26_MB_DEPTH),
        .S_AXIS_BRAM_27_MB_DEPTH(S_AXIS_BRAM_27_MB_DEPTH),
        .S_AXIS_BRAM_28_MB_DEPTH(S_AXIS_BRAM_28_MB_DEPTH),
        .S_AXIS_BRAM_29_MB_DEPTH(S_AXIS_BRAM_29_MB_DEPTH),
        .S_AXIS_BRAM_30_MB_DEPTH(S_AXIS_BRAM_30_MB_DEPTH),
        .S_AXIS_BRAM_31_MB_DEPTH(S_AXIS_BRAM_31_MB_DEPTH),
        .S_AXIS_BRAM_32_MB_DEPTH(S_AXIS_BRAM_32_MB_DEPTH),
        .S_AXIS_BRAM_33_MB_DEPTH(S_AXIS_BRAM_33_MB_DEPTH),
        .S_AXIS_BRAM_34_MB_DEPTH(S_AXIS_BRAM_34_MB_DEPTH),
        .S_AXIS_BRAM_35_MB_DEPTH(S_AXIS_BRAM_35_MB_DEPTH),
        .S_AXIS_BRAM_36_MB_DEPTH(S_AXIS_BRAM_36_MB_DEPTH),
        .S_AXIS_BRAM_37_MB_DEPTH(S_AXIS_BRAM_37_MB_DEPTH),
        .S_AXIS_BRAM_38_MB_DEPTH(S_AXIS_BRAM_38_MB_DEPTH),
        .S_AXIS_BRAM_39_MB_DEPTH(S_AXIS_BRAM_39_MB_DEPTH),
        .S_AXIS_BRAM_40_MB_DEPTH(S_AXIS_BRAM_40_MB_DEPTH),
        .S_AXIS_BRAM_41_MB_DEPTH(S_AXIS_BRAM_41_MB_DEPTH),
        .S_AXIS_BRAM_42_MB_DEPTH(S_AXIS_BRAM_42_MB_DEPTH),
        .S_AXIS_BRAM_43_MB_DEPTH(S_AXIS_BRAM_43_MB_DEPTH),
        .S_AXIS_BRAM_44_MB_DEPTH(S_AXIS_BRAM_44_MB_DEPTH),
        .S_AXIS_BRAM_45_MB_DEPTH(S_AXIS_BRAM_45_MB_DEPTH),
        .S_AXIS_BRAM_46_MB_DEPTH(S_AXIS_BRAM_46_MB_DEPTH),
        .S_AXIS_BRAM_47_MB_DEPTH(S_AXIS_BRAM_47_MB_DEPTH),
        .S_AXIS_BRAM_48_MB_DEPTH(S_AXIS_BRAM_48_MB_DEPTH),
        .S_AXIS_BRAM_49_MB_DEPTH(S_AXIS_BRAM_49_MB_DEPTH),
        .S_AXIS_BRAM_50_MB_DEPTH(S_AXIS_BRAM_50_MB_DEPTH),
        .S_AXIS_BRAM_51_MB_DEPTH(S_AXIS_BRAM_51_MB_DEPTH),
        .S_AXIS_BRAM_52_MB_DEPTH(S_AXIS_BRAM_52_MB_DEPTH),
        .S_AXIS_BRAM_53_MB_DEPTH(S_AXIS_BRAM_53_MB_DEPTH),
        .S_AXIS_BRAM_54_MB_DEPTH(S_AXIS_BRAM_54_MB_DEPTH),
        .S_AXIS_BRAM_55_MB_DEPTH(S_AXIS_BRAM_55_MB_DEPTH),
        .S_AXIS_BRAM_56_MB_DEPTH(S_AXIS_BRAM_56_MB_DEPTH),
        .S_AXIS_BRAM_57_MB_DEPTH(S_AXIS_BRAM_57_MB_DEPTH),
        .S_AXIS_BRAM_58_MB_DEPTH(S_AXIS_BRAM_58_MB_DEPTH),
        .S_AXIS_BRAM_59_MB_DEPTH(S_AXIS_BRAM_59_MB_DEPTH),
        .S_AXIS_BRAM_60_MB_DEPTH(S_AXIS_BRAM_60_MB_DEPTH),
        .S_AXIS_BRAM_61_MB_DEPTH(S_AXIS_BRAM_61_MB_DEPTH),
        .S_AXIS_BRAM_62_MB_DEPTH(S_AXIS_BRAM_62_MB_DEPTH),
        .S_AXIS_BRAM_63_MB_DEPTH(S_AXIS_BRAM_63_MB_DEPTH),
        .S_AXIS_BRAM_64_MB_DEPTH(S_AXIS_BRAM_64_MB_DEPTH),
        .S_AXIS_BRAM_65_MB_DEPTH(S_AXIS_BRAM_65_MB_DEPTH),
        .S_AXIS_BRAM_66_MB_DEPTH(S_AXIS_BRAM_66_MB_DEPTH),
        .S_AXIS_BRAM_67_MB_DEPTH(S_AXIS_BRAM_67_MB_DEPTH),
        .S_AXIS_BRAM_68_MB_DEPTH(S_AXIS_BRAM_68_MB_DEPTH),
        .S_AXIS_BRAM_69_MB_DEPTH(S_AXIS_BRAM_69_MB_DEPTH),
        .S_AXIS_BRAM_70_MB_DEPTH(S_AXIS_BRAM_70_MB_DEPTH),
        .S_AXIS_BRAM_71_MB_DEPTH(S_AXIS_BRAM_71_MB_DEPTH),
        .S_AXIS_BRAM_72_MB_DEPTH(S_AXIS_BRAM_72_MB_DEPTH),
        .S_AXIS_BRAM_73_MB_DEPTH(S_AXIS_BRAM_73_MB_DEPTH),
        .S_AXIS_BRAM_74_MB_DEPTH(S_AXIS_BRAM_74_MB_DEPTH),
        .S_AXIS_BRAM_75_MB_DEPTH(S_AXIS_BRAM_75_MB_DEPTH),
        .S_AXIS_BRAM_76_MB_DEPTH(S_AXIS_BRAM_76_MB_DEPTH),
        .S_AXIS_BRAM_77_MB_DEPTH(S_AXIS_BRAM_77_MB_DEPTH),
        .S_AXIS_BRAM_78_MB_DEPTH(S_AXIS_BRAM_78_MB_DEPTH),
        .S_AXIS_BRAM_79_MB_DEPTH(S_AXIS_BRAM_79_MB_DEPTH),
        .S_AXIS_BRAM_80_MB_DEPTH(S_AXIS_BRAM_80_MB_DEPTH),
        .S_AXIS_BRAM_81_MB_DEPTH(S_AXIS_BRAM_81_MB_DEPTH),
        .S_AXIS_BRAM_82_MB_DEPTH(S_AXIS_BRAM_82_MB_DEPTH),
        .S_AXIS_BRAM_83_MB_DEPTH(S_AXIS_BRAM_83_MB_DEPTH),
        .S_AXIS_BRAM_84_MB_DEPTH(S_AXIS_BRAM_84_MB_DEPTH),
        .S_AXIS_BRAM_85_MB_DEPTH(S_AXIS_BRAM_85_MB_DEPTH),
        .S_AXIS_BRAM_86_MB_DEPTH(S_AXIS_BRAM_86_MB_DEPTH),
        .S_AXIS_BRAM_87_MB_DEPTH(S_AXIS_BRAM_87_MB_DEPTH),
        .S_AXIS_BRAM_88_MB_DEPTH(S_AXIS_BRAM_88_MB_DEPTH),
        .S_AXIS_BRAM_89_MB_DEPTH(S_AXIS_BRAM_89_MB_DEPTH),
        .S_AXIS_BRAM_90_MB_DEPTH(S_AXIS_BRAM_90_MB_DEPTH),
        .S_AXIS_BRAM_91_MB_DEPTH(S_AXIS_BRAM_91_MB_DEPTH),
        .S_AXIS_BRAM_92_MB_DEPTH(S_AXIS_BRAM_92_MB_DEPTH),
        .S_AXIS_BRAM_93_MB_DEPTH(S_AXIS_BRAM_93_MB_DEPTH),
        .S_AXIS_BRAM_94_MB_DEPTH(S_AXIS_BRAM_94_MB_DEPTH),
        .S_AXIS_BRAM_95_MB_DEPTH(S_AXIS_BRAM_95_MB_DEPTH),
        .S_AXIS_BRAM_96_MB_DEPTH(S_AXIS_BRAM_96_MB_DEPTH),
        .S_AXIS_BRAM_97_MB_DEPTH(S_AXIS_BRAM_97_MB_DEPTH),
        .S_AXIS_BRAM_98_MB_DEPTH(S_AXIS_BRAM_98_MB_DEPTH),
        .S_AXIS_BRAM_99_MB_DEPTH(S_AXIS_BRAM_99_MB_DEPTH),
        .S_AXIS_BRAM_100_MB_DEPTH(S_AXIS_BRAM_100_MB_DEPTH),
        .S_AXIS_BRAM_101_MB_DEPTH(S_AXIS_BRAM_101_MB_DEPTH),
        .S_AXIS_BRAM_102_MB_DEPTH(S_AXIS_BRAM_102_MB_DEPTH),
        .S_AXIS_BRAM_103_MB_DEPTH(S_AXIS_BRAM_103_MB_DEPTH),
        .S_AXIS_BRAM_104_MB_DEPTH(S_AXIS_BRAM_104_MB_DEPTH),
        .S_AXIS_BRAM_105_MB_DEPTH(S_AXIS_BRAM_105_MB_DEPTH),
        .S_AXIS_BRAM_106_MB_DEPTH(S_AXIS_BRAM_106_MB_DEPTH),
        .S_AXIS_BRAM_107_MB_DEPTH(S_AXIS_BRAM_107_MB_DEPTH),
        .S_AXIS_BRAM_108_MB_DEPTH(S_AXIS_BRAM_108_MB_DEPTH),
        .S_AXIS_BRAM_109_MB_DEPTH(S_AXIS_BRAM_109_MB_DEPTH),
        .S_AXIS_BRAM_110_MB_DEPTH(S_AXIS_BRAM_110_MB_DEPTH),
        .S_AXIS_BRAM_111_MB_DEPTH(S_AXIS_BRAM_111_MB_DEPTH),
        .S_AXIS_BRAM_112_MB_DEPTH(S_AXIS_BRAM_112_MB_DEPTH),
        .S_AXIS_BRAM_113_MB_DEPTH(S_AXIS_BRAM_113_MB_DEPTH),
        .S_AXIS_BRAM_114_MB_DEPTH(S_AXIS_BRAM_114_MB_DEPTH),
        .S_AXIS_BRAM_115_MB_DEPTH(S_AXIS_BRAM_115_MB_DEPTH),
        .S_AXIS_BRAM_116_MB_DEPTH(S_AXIS_BRAM_116_MB_DEPTH),
        .S_AXIS_BRAM_117_MB_DEPTH(S_AXIS_BRAM_117_MB_DEPTH),
        .S_AXIS_BRAM_118_MB_DEPTH(S_AXIS_BRAM_118_MB_DEPTH),
        .S_AXIS_BRAM_119_MB_DEPTH(S_AXIS_BRAM_119_MB_DEPTH),
        .S_AXIS_BRAM_120_MB_DEPTH(S_AXIS_BRAM_120_MB_DEPTH),
        .S_AXIS_BRAM_121_MB_DEPTH(S_AXIS_BRAM_121_MB_DEPTH),
        .S_AXIS_BRAM_122_MB_DEPTH(S_AXIS_BRAM_122_MB_DEPTH),
        .S_AXIS_BRAM_123_MB_DEPTH(S_AXIS_BRAM_123_MB_DEPTH),
        .S_AXIS_BRAM_124_MB_DEPTH(S_AXIS_BRAM_124_MB_DEPTH),
        .S_AXIS_BRAM_125_MB_DEPTH(S_AXIS_BRAM_125_MB_DEPTH),
        .S_AXIS_BRAM_126_MB_DEPTH(S_AXIS_BRAM_126_MB_DEPTH),
        .S_AXIS_BRAM_127_MB_DEPTH(S_AXIS_BRAM_127_MB_DEPTH),
        .S_AXIS_BRAM_0_ADDR_WIDTH(S_AXIS_BRAM_0_ADDR_WIDTH),
        .S_AXIS_BRAM_1_ADDR_WIDTH(S_AXIS_BRAM_1_ADDR_WIDTH),
        .S_AXIS_BRAM_2_ADDR_WIDTH(S_AXIS_BRAM_2_ADDR_WIDTH),
        .S_AXIS_BRAM_3_ADDR_WIDTH(S_AXIS_BRAM_3_ADDR_WIDTH),
        .S_AXIS_BRAM_4_ADDR_WIDTH(S_AXIS_BRAM_4_ADDR_WIDTH),
        .S_AXIS_BRAM_5_ADDR_WIDTH(S_AXIS_BRAM_5_ADDR_WIDTH),
        .S_AXIS_BRAM_6_ADDR_WIDTH(S_AXIS_BRAM_6_ADDR_WIDTH),
        .S_AXIS_BRAM_7_ADDR_WIDTH(S_AXIS_BRAM_7_ADDR_WIDTH),
        .S_AXIS_BRAM_8_ADDR_WIDTH(S_AXIS_BRAM_8_ADDR_WIDTH),
        .S_AXIS_BRAM_9_ADDR_WIDTH(S_AXIS_BRAM_9_ADDR_WIDTH),
        .S_AXIS_BRAM_10_ADDR_WIDTH(S_AXIS_BRAM_10_ADDR_WIDTH),
        .S_AXIS_BRAM_11_ADDR_WIDTH(S_AXIS_BRAM_11_ADDR_WIDTH),
        .S_AXIS_BRAM_12_ADDR_WIDTH(S_AXIS_BRAM_12_ADDR_WIDTH),
        .S_AXIS_BRAM_13_ADDR_WIDTH(S_AXIS_BRAM_13_ADDR_WIDTH),
        .S_AXIS_BRAM_14_ADDR_WIDTH(S_AXIS_BRAM_14_ADDR_WIDTH),
        .S_AXIS_BRAM_15_ADDR_WIDTH(S_AXIS_BRAM_15_ADDR_WIDTH),
        .S_AXIS_BRAM_16_ADDR_WIDTH(S_AXIS_BRAM_16_ADDR_WIDTH),
        .S_AXIS_BRAM_17_ADDR_WIDTH(S_AXIS_BRAM_17_ADDR_WIDTH),
        .S_AXIS_BRAM_18_ADDR_WIDTH(S_AXIS_BRAM_18_ADDR_WIDTH),
        .S_AXIS_BRAM_19_ADDR_WIDTH(S_AXIS_BRAM_19_ADDR_WIDTH),
        .S_AXIS_BRAM_20_ADDR_WIDTH(S_AXIS_BRAM_20_ADDR_WIDTH),
        .S_AXIS_BRAM_21_ADDR_WIDTH(S_AXIS_BRAM_21_ADDR_WIDTH),
        .S_AXIS_BRAM_22_ADDR_WIDTH(S_AXIS_BRAM_22_ADDR_WIDTH),
        .S_AXIS_BRAM_23_ADDR_WIDTH(S_AXIS_BRAM_23_ADDR_WIDTH),
        .S_AXIS_BRAM_24_ADDR_WIDTH(S_AXIS_BRAM_24_ADDR_WIDTH),
        .S_AXIS_BRAM_25_ADDR_WIDTH(S_AXIS_BRAM_25_ADDR_WIDTH),
        .S_AXIS_BRAM_26_ADDR_WIDTH(S_AXIS_BRAM_26_ADDR_WIDTH),
        .S_AXIS_BRAM_27_ADDR_WIDTH(S_AXIS_BRAM_27_ADDR_WIDTH),
        .S_AXIS_BRAM_28_ADDR_WIDTH(S_AXIS_BRAM_28_ADDR_WIDTH),
        .S_AXIS_BRAM_29_ADDR_WIDTH(S_AXIS_BRAM_29_ADDR_WIDTH),
        .S_AXIS_BRAM_30_ADDR_WIDTH(S_AXIS_BRAM_30_ADDR_WIDTH),
        .S_AXIS_BRAM_31_ADDR_WIDTH(S_AXIS_BRAM_31_ADDR_WIDTH),
        .S_AXIS_BRAM_32_ADDR_WIDTH(S_AXIS_BRAM_32_ADDR_WIDTH),
        .S_AXIS_BRAM_33_ADDR_WIDTH(S_AXIS_BRAM_33_ADDR_WIDTH),
        .S_AXIS_BRAM_34_ADDR_WIDTH(S_AXIS_BRAM_34_ADDR_WIDTH),
        .S_AXIS_BRAM_35_ADDR_WIDTH(S_AXIS_BRAM_35_ADDR_WIDTH),
        .S_AXIS_BRAM_36_ADDR_WIDTH(S_AXIS_BRAM_36_ADDR_WIDTH),
        .S_AXIS_BRAM_37_ADDR_WIDTH(S_AXIS_BRAM_37_ADDR_WIDTH),
        .S_AXIS_BRAM_38_ADDR_WIDTH(S_AXIS_BRAM_38_ADDR_WIDTH),
        .S_AXIS_BRAM_39_ADDR_WIDTH(S_AXIS_BRAM_39_ADDR_WIDTH),
        .S_AXIS_BRAM_40_ADDR_WIDTH(S_AXIS_BRAM_40_ADDR_WIDTH),
        .S_AXIS_BRAM_41_ADDR_WIDTH(S_AXIS_BRAM_41_ADDR_WIDTH),
        .S_AXIS_BRAM_42_ADDR_WIDTH(S_AXIS_BRAM_42_ADDR_WIDTH),
        .S_AXIS_BRAM_43_ADDR_WIDTH(S_AXIS_BRAM_43_ADDR_WIDTH),
        .S_AXIS_BRAM_44_ADDR_WIDTH(S_AXIS_BRAM_44_ADDR_WIDTH),
        .S_AXIS_BRAM_45_ADDR_WIDTH(S_AXIS_BRAM_45_ADDR_WIDTH),
        .S_AXIS_BRAM_46_ADDR_WIDTH(S_AXIS_BRAM_46_ADDR_WIDTH),
        .S_AXIS_BRAM_47_ADDR_WIDTH(S_AXIS_BRAM_47_ADDR_WIDTH),
        .S_AXIS_BRAM_48_ADDR_WIDTH(S_AXIS_BRAM_48_ADDR_WIDTH),
        .S_AXIS_BRAM_49_ADDR_WIDTH(S_AXIS_BRAM_49_ADDR_WIDTH),
        .S_AXIS_BRAM_50_ADDR_WIDTH(S_AXIS_BRAM_50_ADDR_WIDTH),
        .S_AXIS_BRAM_51_ADDR_WIDTH(S_AXIS_BRAM_51_ADDR_WIDTH),
        .S_AXIS_BRAM_52_ADDR_WIDTH(S_AXIS_BRAM_52_ADDR_WIDTH),
        .S_AXIS_BRAM_53_ADDR_WIDTH(S_AXIS_BRAM_53_ADDR_WIDTH),
        .S_AXIS_BRAM_54_ADDR_WIDTH(S_AXIS_BRAM_54_ADDR_WIDTH),
        .S_AXIS_BRAM_55_ADDR_WIDTH(S_AXIS_BRAM_55_ADDR_WIDTH),
        .S_AXIS_BRAM_56_ADDR_WIDTH(S_AXIS_BRAM_56_ADDR_WIDTH),
        .S_AXIS_BRAM_57_ADDR_WIDTH(S_AXIS_BRAM_57_ADDR_WIDTH),
        .S_AXIS_BRAM_58_ADDR_WIDTH(S_AXIS_BRAM_58_ADDR_WIDTH),
        .S_AXIS_BRAM_59_ADDR_WIDTH(S_AXIS_BRAM_59_ADDR_WIDTH),
        .S_AXIS_BRAM_60_ADDR_WIDTH(S_AXIS_BRAM_60_ADDR_WIDTH),
        .S_AXIS_BRAM_61_ADDR_WIDTH(S_AXIS_BRAM_61_ADDR_WIDTH),
        .S_AXIS_BRAM_62_ADDR_WIDTH(S_AXIS_BRAM_62_ADDR_WIDTH),
        .S_AXIS_BRAM_63_ADDR_WIDTH(S_AXIS_BRAM_63_ADDR_WIDTH),
        .S_AXIS_BRAM_64_ADDR_WIDTH(S_AXIS_BRAM_64_ADDR_WIDTH),
        .S_AXIS_BRAM_65_ADDR_WIDTH(S_AXIS_BRAM_65_ADDR_WIDTH),
        .S_AXIS_BRAM_66_ADDR_WIDTH(S_AXIS_BRAM_66_ADDR_WIDTH),
        .S_AXIS_BRAM_67_ADDR_WIDTH(S_AXIS_BRAM_67_ADDR_WIDTH),
        .S_AXIS_BRAM_68_ADDR_WIDTH(S_AXIS_BRAM_68_ADDR_WIDTH),
        .S_AXIS_BRAM_69_ADDR_WIDTH(S_AXIS_BRAM_69_ADDR_WIDTH),
        .S_AXIS_BRAM_70_ADDR_WIDTH(S_AXIS_BRAM_70_ADDR_WIDTH),
        .S_AXIS_BRAM_71_ADDR_WIDTH(S_AXIS_BRAM_71_ADDR_WIDTH),
        .S_AXIS_BRAM_72_ADDR_WIDTH(S_AXIS_BRAM_72_ADDR_WIDTH),
        .S_AXIS_BRAM_73_ADDR_WIDTH(S_AXIS_BRAM_73_ADDR_WIDTH),
        .S_AXIS_BRAM_74_ADDR_WIDTH(S_AXIS_BRAM_74_ADDR_WIDTH),
        .S_AXIS_BRAM_75_ADDR_WIDTH(S_AXIS_BRAM_75_ADDR_WIDTH),
        .S_AXIS_BRAM_76_ADDR_WIDTH(S_AXIS_BRAM_76_ADDR_WIDTH),
        .S_AXIS_BRAM_77_ADDR_WIDTH(S_AXIS_BRAM_77_ADDR_WIDTH),
        .S_AXIS_BRAM_78_ADDR_WIDTH(S_AXIS_BRAM_78_ADDR_WIDTH),
        .S_AXIS_BRAM_79_ADDR_WIDTH(S_AXIS_BRAM_79_ADDR_WIDTH),
        .S_AXIS_BRAM_80_ADDR_WIDTH(S_AXIS_BRAM_80_ADDR_WIDTH),
        .S_AXIS_BRAM_81_ADDR_WIDTH(S_AXIS_BRAM_81_ADDR_WIDTH),
        .S_AXIS_BRAM_82_ADDR_WIDTH(S_AXIS_BRAM_82_ADDR_WIDTH),
        .S_AXIS_BRAM_83_ADDR_WIDTH(S_AXIS_BRAM_83_ADDR_WIDTH),
        .S_AXIS_BRAM_84_ADDR_WIDTH(S_AXIS_BRAM_84_ADDR_WIDTH),
        .S_AXIS_BRAM_85_ADDR_WIDTH(S_AXIS_BRAM_85_ADDR_WIDTH),
        .S_AXIS_BRAM_86_ADDR_WIDTH(S_AXIS_BRAM_86_ADDR_WIDTH),
        .S_AXIS_BRAM_87_ADDR_WIDTH(S_AXIS_BRAM_87_ADDR_WIDTH),
        .S_AXIS_BRAM_88_ADDR_WIDTH(S_AXIS_BRAM_88_ADDR_WIDTH),
        .S_AXIS_BRAM_89_ADDR_WIDTH(S_AXIS_BRAM_89_ADDR_WIDTH),
        .S_AXIS_BRAM_90_ADDR_WIDTH(S_AXIS_BRAM_90_ADDR_WIDTH),
        .S_AXIS_BRAM_91_ADDR_WIDTH(S_AXIS_BRAM_91_ADDR_WIDTH),
        .S_AXIS_BRAM_92_ADDR_WIDTH(S_AXIS_BRAM_92_ADDR_WIDTH),
        .S_AXIS_BRAM_93_ADDR_WIDTH(S_AXIS_BRAM_93_ADDR_WIDTH),
        .S_AXIS_BRAM_94_ADDR_WIDTH(S_AXIS_BRAM_94_ADDR_WIDTH),
        .S_AXIS_BRAM_95_ADDR_WIDTH(S_AXIS_BRAM_95_ADDR_WIDTH),
        .S_AXIS_BRAM_96_ADDR_WIDTH(S_AXIS_BRAM_96_ADDR_WIDTH),
        .S_AXIS_BRAM_97_ADDR_WIDTH(S_AXIS_BRAM_97_ADDR_WIDTH),
        .S_AXIS_BRAM_98_ADDR_WIDTH(S_AXIS_BRAM_98_ADDR_WIDTH),
        .S_AXIS_BRAM_99_ADDR_WIDTH(S_AXIS_BRAM_99_ADDR_WIDTH),
        .S_AXIS_BRAM_100_ADDR_WIDTH(S_AXIS_BRAM_100_ADDR_WIDTH),
        .S_AXIS_BRAM_101_ADDR_WIDTH(S_AXIS_BRAM_101_ADDR_WIDTH),
        .S_AXIS_BRAM_102_ADDR_WIDTH(S_AXIS_BRAM_102_ADDR_WIDTH),
        .S_AXIS_BRAM_103_ADDR_WIDTH(S_AXIS_BRAM_103_ADDR_WIDTH),
        .S_AXIS_BRAM_104_ADDR_WIDTH(S_AXIS_BRAM_104_ADDR_WIDTH),
        .S_AXIS_BRAM_105_ADDR_WIDTH(S_AXIS_BRAM_105_ADDR_WIDTH),
        .S_AXIS_BRAM_106_ADDR_WIDTH(S_AXIS_BRAM_106_ADDR_WIDTH),
        .S_AXIS_BRAM_107_ADDR_WIDTH(S_AXIS_BRAM_107_ADDR_WIDTH),
        .S_AXIS_BRAM_108_ADDR_WIDTH(S_AXIS_BRAM_108_ADDR_WIDTH),
        .S_AXIS_BRAM_109_ADDR_WIDTH(S_AXIS_BRAM_109_ADDR_WIDTH),
        .S_AXIS_BRAM_110_ADDR_WIDTH(S_AXIS_BRAM_110_ADDR_WIDTH),
        .S_AXIS_BRAM_111_ADDR_WIDTH(S_AXIS_BRAM_111_ADDR_WIDTH),
        .S_AXIS_BRAM_112_ADDR_WIDTH(S_AXIS_BRAM_112_ADDR_WIDTH),
        .S_AXIS_BRAM_113_ADDR_WIDTH(S_AXIS_BRAM_113_ADDR_WIDTH),
        .S_AXIS_BRAM_114_ADDR_WIDTH(S_AXIS_BRAM_114_ADDR_WIDTH),
        .S_AXIS_BRAM_115_ADDR_WIDTH(S_AXIS_BRAM_115_ADDR_WIDTH),
        .S_AXIS_BRAM_116_ADDR_WIDTH(S_AXIS_BRAM_116_ADDR_WIDTH),
        .S_AXIS_BRAM_117_ADDR_WIDTH(S_AXIS_BRAM_117_ADDR_WIDTH),
        .S_AXIS_BRAM_118_ADDR_WIDTH(S_AXIS_BRAM_118_ADDR_WIDTH),
        .S_AXIS_BRAM_119_ADDR_WIDTH(S_AXIS_BRAM_119_ADDR_WIDTH),
        .S_AXIS_BRAM_120_ADDR_WIDTH(S_AXIS_BRAM_120_ADDR_WIDTH),
        .S_AXIS_BRAM_121_ADDR_WIDTH(S_AXIS_BRAM_121_ADDR_WIDTH),
        .S_AXIS_BRAM_122_ADDR_WIDTH(S_AXIS_BRAM_122_ADDR_WIDTH),
        .S_AXIS_BRAM_123_ADDR_WIDTH(S_AXIS_BRAM_123_ADDR_WIDTH),
        .S_AXIS_BRAM_124_ADDR_WIDTH(S_AXIS_BRAM_124_ADDR_WIDTH),
        .S_AXIS_BRAM_125_ADDR_WIDTH(S_AXIS_BRAM_125_ADDR_WIDTH),
        .S_AXIS_BRAM_126_ADDR_WIDTH(S_AXIS_BRAM_126_ADDR_WIDTH),
        .S_AXIS_BRAM_127_ADDR_WIDTH(S_AXIS_BRAM_127_ADDR_WIDTH)
    ) in_bram_args_i (
        .acc_clk(acc_aclk),
        .acc_aresetn(acc_aresetn),
        .in_bram_allow_in(inbram_ctrl_allow),
        .in_bram_allow_out(outbram_ctrl_allow),
        .acc_start(ap_start_single),
        .acc_done(ap_done),
        .in_bram_ready(inbram_ctrl_ready),
        .inout_bram_ready(inoutbram_ctrl_ready),
        .s_axis_bram_0_aclk(s_axis_bram_0_aclk),
        .s_axis_bram_0_aresetn(s_axis_bram_0_aresetn),
        .s_axis_bram_0_tlast(s_axis_bram_0_tlast),
        .s_axis_bram_0_tvalid(s_axis_bram_0_tvalid),
        .s_axis_bram_0_tkeep(s_axis_bram_0_tkeep),
        .s_axis_bram_0_tstrb(s_axis_bram_0_tstrb),
        .s_axis_bram_0_tdata(s_axis_bram_0_tdata),
        .s_axis_bram_0_tready(s_axis_bram_0_tready),
        .ap_bram_0_addr0(ap_bram_iarg_0_addr0),
        .ap_bram_0_din0(ap_bram_iarg_0_din0),
        .ap_bram_0_dout0(ap_bram_iarg_0_dout0),
        .ap_bram_0_we0(ap_bram_iarg_0_we0),
        .ap_bram_0_en0(ap_bram_iarg_0_en0),
        .ap_bram_0_addr1(ap_bram_iarg_0_addr1),
        .ap_bram_0_din1(ap_bram_iarg_0_din1),
        .ap_bram_0_dout1(ap_bram_iarg_0_dout1),
        .ap_bram_0_we1(ap_bram_iarg_0_we1),
        .ap_bram_0_en1(ap_bram_iarg_0_en1),
        .s_axis_bram_1_aclk(s_axis_bram_1_aclk),
        .s_axis_bram_1_aresetn(s_axis_bram_1_aresetn),
        .s_axis_bram_1_tlast(s_axis_bram_1_tlast),
        .s_axis_bram_1_tvalid(s_axis_bram_1_tvalid),
        .s_axis_bram_1_tkeep(s_axis_bram_1_tkeep),
        .s_axis_bram_1_tstrb(s_axis_bram_1_tstrb),
        .s_axis_bram_1_tdata(s_axis_bram_1_tdata),
        .s_axis_bram_1_tready(s_axis_bram_1_tready),
        .ap_bram_1_addr0(ap_bram_iarg_1_addr0),
        .ap_bram_1_din0(ap_bram_iarg_1_din0),
        .ap_bram_1_dout0(ap_bram_iarg_1_dout0),
        .ap_bram_1_we0(ap_bram_iarg_1_we0),
        .ap_bram_1_en0(ap_bram_iarg_1_en0),
        .ap_bram_1_addr1(ap_bram_iarg_1_addr1),
        .ap_bram_1_din1(ap_bram_iarg_1_din1),
        .ap_bram_1_dout1(ap_bram_iarg_1_dout1),
        .ap_bram_1_we1(ap_bram_iarg_1_we1),
        .ap_bram_1_en1(ap_bram_iarg_1_en1),
        .s_axis_bram_2_aclk(s_axis_bram_2_aclk),
        .s_axis_bram_2_aresetn(s_axis_bram_2_aresetn),
        .s_axis_bram_2_tlast(s_axis_bram_2_tlast),
        .s_axis_bram_2_tvalid(s_axis_bram_2_tvalid),
        .s_axis_bram_2_tkeep(s_axis_bram_2_tkeep),
        .s_axis_bram_2_tstrb(s_axis_bram_2_tstrb),
        .s_axis_bram_2_tdata(s_axis_bram_2_tdata),
        .s_axis_bram_2_tready(s_axis_bram_2_tready),
        .ap_bram_2_addr0(ap_bram_iarg_2_addr0),
        .ap_bram_2_din0(ap_bram_iarg_2_din0),
        .ap_bram_2_dout0(ap_bram_iarg_2_dout0),
        .ap_bram_2_we0(ap_bram_iarg_2_we0),
        .ap_bram_2_en0(ap_bram_iarg_2_en0),
        .ap_bram_2_addr1(ap_bram_iarg_2_addr1),
        .ap_bram_2_din1(ap_bram_iarg_2_din1),
        .ap_bram_2_dout1(ap_bram_iarg_2_dout1),
        .ap_bram_2_we1(ap_bram_iarg_2_we1),
        .ap_bram_2_en1(ap_bram_iarg_2_en1),
        .s_axis_bram_3_aclk(s_axis_bram_3_aclk),
        .s_axis_bram_3_aresetn(s_axis_bram_3_aresetn),
        .s_axis_bram_3_tlast(s_axis_bram_3_tlast),
        .s_axis_bram_3_tvalid(s_axis_bram_3_tvalid),
        .s_axis_bram_3_tkeep(s_axis_bram_3_tkeep),
        .s_axis_bram_3_tstrb(s_axis_bram_3_tstrb),
        .s_axis_bram_3_tdata(s_axis_bram_3_tdata),
        .s_axis_bram_3_tready(s_axis_bram_3_tready),
        .ap_bram_3_addr0(ap_bram_iarg_3_addr0),
        .ap_bram_3_din0(ap_bram_iarg_3_din0),
        .ap_bram_3_dout0(ap_bram_iarg_3_dout0),
        .ap_bram_3_we0(ap_bram_iarg_3_we0),
        .ap_bram_3_en0(ap_bram_iarg_3_en0),
        .ap_bram_3_addr1(ap_bram_iarg_3_addr1),
        .ap_bram_3_din1(ap_bram_iarg_3_din1),
        .ap_bram_3_dout1(ap_bram_iarg_3_dout1),
        .ap_bram_3_we1(ap_bram_iarg_3_we1),
        .ap_bram_3_en1(ap_bram_iarg_3_en1),
        .s_axis_bram_4_aclk(s_axis_bram_4_aclk),
        .s_axis_bram_4_aresetn(s_axis_bram_4_aresetn),
        .s_axis_bram_4_tlast(s_axis_bram_4_tlast),
        .s_axis_bram_4_tvalid(s_axis_bram_4_tvalid),
        .s_axis_bram_4_tkeep(s_axis_bram_4_tkeep),
        .s_axis_bram_4_tstrb(s_axis_bram_4_tstrb),
        .s_axis_bram_4_tdata(s_axis_bram_4_tdata),
        .s_axis_bram_4_tready(s_axis_bram_4_tready),
        .ap_bram_4_addr0(ap_bram_iarg_4_addr0),
        .ap_bram_4_din0(ap_bram_iarg_4_din0),
        .ap_bram_4_dout0(ap_bram_iarg_4_dout0),
        .ap_bram_4_we0(ap_bram_iarg_4_we0),
        .ap_bram_4_en0(ap_bram_iarg_4_en0),
        .ap_bram_4_addr1(ap_bram_iarg_4_addr1),
        .ap_bram_4_din1(ap_bram_iarg_4_din1),
        .ap_bram_4_dout1(ap_bram_iarg_4_dout1),
        .ap_bram_4_we1(ap_bram_iarg_4_we1),
        .ap_bram_4_en1(ap_bram_iarg_4_en1),
        .s_axis_bram_5_aclk(s_axis_bram_5_aclk),
        .s_axis_bram_5_aresetn(s_axis_bram_5_aresetn),
        .s_axis_bram_5_tlast(s_axis_bram_5_tlast),
        .s_axis_bram_5_tvalid(s_axis_bram_5_tvalid),
        .s_axis_bram_5_tkeep(s_axis_bram_5_tkeep),
        .s_axis_bram_5_tstrb(s_axis_bram_5_tstrb),
        .s_axis_bram_5_tdata(s_axis_bram_5_tdata),
        .s_axis_bram_5_tready(s_axis_bram_5_tready),
        .ap_bram_5_addr0(ap_bram_iarg_5_addr0),
        .ap_bram_5_din0(ap_bram_iarg_5_din0),
        .ap_bram_5_dout0(ap_bram_iarg_5_dout0),
        .ap_bram_5_we0(ap_bram_iarg_5_we0),
        .ap_bram_5_en0(ap_bram_iarg_5_en0),
        .ap_bram_5_addr1(ap_bram_iarg_5_addr1),
        .ap_bram_5_din1(ap_bram_iarg_5_din1),
        .ap_bram_5_dout1(ap_bram_iarg_5_dout1),
        .ap_bram_5_we1(ap_bram_iarg_5_we1),
        .ap_bram_5_en1(ap_bram_iarg_5_en1),
        .s_axis_bram_6_aclk(s_axis_bram_6_aclk),
        .s_axis_bram_6_aresetn(s_axis_bram_6_aresetn),
        .s_axis_bram_6_tlast(s_axis_bram_6_tlast),
        .s_axis_bram_6_tvalid(s_axis_bram_6_tvalid),
        .s_axis_bram_6_tkeep(s_axis_bram_6_tkeep),
        .s_axis_bram_6_tstrb(s_axis_bram_6_tstrb),
        .s_axis_bram_6_tdata(s_axis_bram_6_tdata),
        .s_axis_bram_6_tready(s_axis_bram_6_tready),
        .ap_bram_6_addr0(ap_bram_iarg_6_addr0),
        .ap_bram_6_din0(ap_bram_iarg_6_din0),
        .ap_bram_6_dout0(ap_bram_iarg_6_dout0),
        .ap_bram_6_we0(ap_bram_iarg_6_we0),
        .ap_bram_6_en0(ap_bram_iarg_6_en0),
        .ap_bram_6_addr1(ap_bram_iarg_6_addr1),
        .ap_bram_6_din1(ap_bram_iarg_6_din1),
        .ap_bram_6_dout1(ap_bram_iarg_6_dout1),
        .ap_bram_6_we1(ap_bram_iarg_6_we1),
        .ap_bram_6_en1(ap_bram_iarg_6_en1),
        .s_axis_bram_7_aclk(s_axis_bram_7_aclk),
        .s_axis_bram_7_aresetn(s_axis_bram_7_aresetn),
        .s_axis_bram_7_tlast(s_axis_bram_7_tlast),
        .s_axis_bram_7_tvalid(s_axis_bram_7_tvalid),
        .s_axis_bram_7_tkeep(s_axis_bram_7_tkeep),
        .s_axis_bram_7_tstrb(s_axis_bram_7_tstrb),
        .s_axis_bram_7_tdata(s_axis_bram_7_tdata),
        .s_axis_bram_7_tready(s_axis_bram_7_tready),
        .ap_bram_7_addr0(ap_bram_iarg_7_addr0),
        .ap_bram_7_din0(ap_bram_iarg_7_din0),
        .ap_bram_7_dout0(ap_bram_iarg_7_dout0),
        .ap_bram_7_we0(ap_bram_iarg_7_we0),
        .ap_bram_7_en0(ap_bram_iarg_7_en0),
        .ap_bram_7_addr1(ap_bram_iarg_7_addr1),
        .ap_bram_7_din1(ap_bram_iarg_7_din1),
        .ap_bram_7_dout1(ap_bram_iarg_7_dout1),
        .ap_bram_7_we1(ap_bram_iarg_7_we1),
        .ap_bram_7_en1(ap_bram_iarg_7_en1),
        .s_axis_bram_8_aclk(s_axis_bram_8_aclk),
        .s_axis_bram_8_aresetn(s_axis_bram_8_aresetn),
        .s_axis_bram_8_tlast(s_axis_bram_8_tlast),
        .s_axis_bram_8_tvalid(s_axis_bram_8_tvalid),
        .s_axis_bram_8_tkeep(s_axis_bram_8_tkeep),
        .s_axis_bram_8_tstrb(s_axis_bram_8_tstrb),
        .s_axis_bram_8_tdata(s_axis_bram_8_tdata),
        .s_axis_bram_8_tready(s_axis_bram_8_tready),
        .ap_bram_8_addr0(ap_bram_iarg_8_addr0),
        .ap_bram_8_din0(ap_bram_iarg_8_din0),
        .ap_bram_8_dout0(ap_bram_iarg_8_dout0),
        .ap_bram_8_we0(ap_bram_iarg_8_we0),
        .ap_bram_8_en0(ap_bram_iarg_8_en0),
        .ap_bram_8_addr1(ap_bram_iarg_8_addr1),
        .ap_bram_8_din1(ap_bram_iarg_8_din1),
        .ap_bram_8_dout1(ap_bram_iarg_8_dout1),
        .ap_bram_8_we1(ap_bram_iarg_8_we1),
        .ap_bram_8_en1(ap_bram_iarg_8_en1),
        .s_axis_bram_9_aclk(s_axis_bram_9_aclk),
        .s_axis_bram_9_aresetn(s_axis_bram_9_aresetn),
        .s_axis_bram_9_tlast(s_axis_bram_9_tlast),
        .s_axis_bram_9_tvalid(s_axis_bram_9_tvalid),
        .s_axis_bram_9_tkeep(s_axis_bram_9_tkeep),
        .s_axis_bram_9_tstrb(s_axis_bram_9_tstrb),
        .s_axis_bram_9_tdata(s_axis_bram_9_tdata),
        .s_axis_bram_9_tready(s_axis_bram_9_tready),
        .ap_bram_9_addr0(ap_bram_iarg_9_addr0),
        .ap_bram_9_din0(ap_bram_iarg_9_din0),
        .ap_bram_9_dout0(ap_bram_iarg_9_dout0),
        .ap_bram_9_we0(ap_bram_iarg_9_we0),
        .ap_bram_9_en0(ap_bram_iarg_9_en0),
        .ap_bram_9_addr1(ap_bram_iarg_9_addr1),
        .ap_bram_9_din1(ap_bram_iarg_9_din1),
        .ap_bram_9_dout1(ap_bram_iarg_9_dout1),
        .ap_bram_9_we1(ap_bram_iarg_9_we1),
        .ap_bram_9_en1(ap_bram_iarg_9_en1),
        .s_axis_bram_10_aclk(s_axis_bram_10_aclk),
        .s_axis_bram_10_aresetn(s_axis_bram_10_aresetn),
        .s_axis_bram_10_tlast(s_axis_bram_10_tlast),
        .s_axis_bram_10_tvalid(s_axis_bram_10_tvalid),
        .s_axis_bram_10_tkeep(s_axis_bram_10_tkeep),
        .s_axis_bram_10_tstrb(s_axis_bram_10_tstrb),
        .s_axis_bram_10_tdata(s_axis_bram_10_tdata),
        .s_axis_bram_10_tready(s_axis_bram_10_tready),
        .ap_bram_10_addr0(ap_bram_iarg_10_addr0),
        .ap_bram_10_din0(ap_bram_iarg_10_din0),
        .ap_bram_10_dout0(ap_bram_iarg_10_dout0),
        .ap_bram_10_we0(ap_bram_iarg_10_we0),
        .ap_bram_10_en0(ap_bram_iarg_10_en0),
        .ap_bram_10_addr1(ap_bram_iarg_10_addr1),
        .ap_bram_10_din1(ap_bram_iarg_10_din1),
        .ap_bram_10_dout1(ap_bram_iarg_10_dout1),
        .ap_bram_10_we1(ap_bram_iarg_10_we1),
        .ap_bram_10_en1(ap_bram_iarg_10_en1),
        .s_axis_bram_11_aclk(s_axis_bram_11_aclk),
        .s_axis_bram_11_aresetn(s_axis_bram_11_aresetn),
        .s_axis_bram_11_tlast(s_axis_bram_11_tlast),
        .s_axis_bram_11_tvalid(s_axis_bram_11_tvalid),
        .s_axis_bram_11_tkeep(s_axis_bram_11_tkeep),
        .s_axis_bram_11_tstrb(s_axis_bram_11_tstrb),
        .s_axis_bram_11_tdata(s_axis_bram_11_tdata),
        .s_axis_bram_11_tready(s_axis_bram_11_tready),
        .ap_bram_11_addr0(ap_bram_iarg_11_addr0),
        .ap_bram_11_din0(ap_bram_iarg_11_din0),
        .ap_bram_11_dout0(ap_bram_iarg_11_dout0),
        .ap_bram_11_we0(ap_bram_iarg_11_we0),
        .ap_bram_11_en0(ap_bram_iarg_11_en0),
        .ap_bram_11_addr1(ap_bram_iarg_11_addr1),
        .ap_bram_11_din1(ap_bram_iarg_11_din1),
        .ap_bram_11_dout1(ap_bram_iarg_11_dout1),
        .ap_bram_11_we1(ap_bram_iarg_11_we1),
        .ap_bram_11_en1(ap_bram_iarg_11_en1),
        .s_axis_bram_12_aclk(s_axis_bram_12_aclk),
        .s_axis_bram_12_aresetn(s_axis_bram_12_aresetn),
        .s_axis_bram_12_tlast(s_axis_bram_12_tlast),
        .s_axis_bram_12_tvalid(s_axis_bram_12_tvalid),
        .s_axis_bram_12_tkeep(s_axis_bram_12_tkeep),
        .s_axis_bram_12_tstrb(s_axis_bram_12_tstrb),
        .s_axis_bram_12_tdata(s_axis_bram_12_tdata),
        .s_axis_bram_12_tready(s_axis_bram_12_tready),
        .ap_bram_12_addr0(ap_bram_iarg_12_addr0),
        .ap_bram_12_din0(ap_bram_iarg_12_din0),
        .ap_bram_12_dout0(ap_bram_iarg_12_dout0),
        .ap_bram_12_we0(ap_bram_iarg_12_we0),
        .ap_bram_12_en0(ap_bram_iarg_12_en0),
        .ap_bram_12_addr1(ap_bram_iarg_12_addr1),
        .ap_bram_12_din1(ap_bram_iarg_12_din1),
        .ap_bram_12_dout1(ap_bram_iarg_12_dout1),
        .ap_bram_12_we1(ap_bram_iarg_12_we1),
        .ap_bram_12_en1(ap_bram_iarg_12_en1),
        .s_axis_bram_13_aclk(s_axis_bram_13_aclk),
        .s_axis_bram_13_aresetn(s_axis_bram_13_aresetn),
        .s_axis_bram_13_tlast(s_axis_bram_13_tlast),
        .s_axis_bram_13_tvalid(s_axis_bram_13_tvalid),
        .s_axis_bram_13_tkeep(s_axis_bram_13_tkeep),
        .s_axis_bram_13_tstrb(s_axis_bram_13_tstrb),
        .s_axis_bram_13_tdata(s_axis_bram_13_tdata),
        .s_axis_bram_13_tready(s_axis_bram_13_tready),
        .ap_bram_13_addr0(ap_bram_iarg_13_addr0),
        .ap_bram_13_din0(ap_bram_iarg_13_din0),
        .ap_bram_13_dout0(ap_bram_iarg_13_dout0),
        .ap_bram_13_we0(ap_bram_iarg_13_we0),
        .ap_bram_13_en0(ap_bram_iarg_13_en0),
        .ap_bram_13_addr1(ap_bram_iarg_13_addr1),
        .ap_bram_13_din1(ap_bram_iarg_13_din1),
        .ap_bram_13_dout1(ap_bram_iarg_13_dout1),
        .ap_bram_13_we1(ap_bram_iarg_13_we1),
        .ap_bram_13_en1(ap_bram_iarg_13_en1),
        .s_axis_bram_14_aclk(s_axis_bram_14_aclk),
        .s_axis_bram_14_aresetn(s_axis_bram_14_aresetn),
        .s_axis_bram_14_tlast(s_axis_bram_14_tlast),
        .s_axis_bram_14_tvalid(s_axis_bram_14_tvalid),
        .s_axis_bram_14_tkeep(s_axis_bram_14_tkeep),
        .s_axis_bram_14_tstrb(s_axis_bram_14_tstrb),
        .s_axis_bram_14_tdata(s_axis_bram_14_tdata),
        .s_axis_bram_14_tready(s_axis_bram_14_tready),
        .ap_bram_14_addr0(ap_bram_iarg_14_addr0),
        .ap_bram_14_din0(ap_bram_iarg_14_din0),
        .ap_bram_14_dout0(ap_bram_iarg_14_dout0),
        .ap_bram_14_we0(ap_bram_iarg_14_we0),
        .ap_bram_14_en0(ap_bram_iarg_14_en0),
        .ap_bram_14_addr1(ap_bram_iarg_14_addr1),
        .ap_bram_14_din1(ap_bram_iarg_14_din1),
        .ap_bram_14_dout1(ap_bram_iarg_14_dout1),
        .ap_bram_14_we1(ap_bram_iarg_14_we1),
        .ap_bram_14_en1(ap_bram_iarg_14_en1),
        .s_axis_bram_15_aclk(s_axis_bram_15_aclk),
        .s_axis_bram_15_aresetn(s_axis_bram_15_aresetn),
        .s_axis_bram_15_tlast(s_axis_bram_15_tlast),
        .s_axis_bram_15_tvalid(s_axis_bram_15_tvalid),
        .s_axis_bram_15_tkeep(s_axis_bram_15_tkeep),
        .s_axis_bram_15_tstrb(s_axis_bram_15_tstrb),
        .s_axis_bram_15_tdata(s_axis_bram_15_tdata),
        .s_axis_bram_15_tready(s_axis_bram_15_tready),
        .ap_bram_15_addr0(ap_bram_iarg_15_addr0),
        .ap_bram_15_din0(ap_bram_iarg_15_din0),
        .ap_bram_15_dout0(ap_bram_iarg_15_dout0),
        .ap_bram_15_we0(ap_bram_iarg_15_we0),
        .ap_bram_15_en0(ap_bram_iarg_15_en0),
        .ap_bram_15_addr1(ap_bram_iarg_15_addr1),
        .ap_bram_15_din1(ap_bram_iarg_15_din1),
        .ap_bram_15_dout1(ap_bram_iarg_15_dout1),
        .ap_bram_15_we1(ap_bram_iarg_15_we1),
        .ap_bram_15_en1(ap_bram_iarg_15_en1),
        .s_axis_bram_16_aclk(s_axis_bram_16_aclk),
        .s_axis_bram_16_aresetn(s_axis_bram_16_aresetn),
        .s_axis_bram_16_tlast(s_axis_bram_16_tlast),
        .s_axis_bram_16_tvalid(s_axis_bram_16_tvalid),
        .s_axis_bram_16_tkeep(s_axis_bram_16_tkeep),
        .s_axis_bram_16_tstrb(s_axis_bram_16_tstrb),
        .s_axis_bram_16_tdata(s_axis_bram_16_tdata),
        .s_axis_bram_16_tready(s_axis_bram_16_tready),
        .ap_bram_16_addr0(ap_bram_iarg_16_addr0),
        .ap_bram_16_din0(ap_bram_iarg_16_din0),
        .ap_bram_16_dout0(ap_bram_iarg_16_dout0),
        .ap_bram_16_we0(ap_bram_iarg_16_we0),
        .ap_bram_16_en0(ap_bram_iarg_16_en0),
        .ap_bram_16_addr1(ap_bram_iarg_16_addr1),
        .ap_bram_16_din1(ap_bram_iarg_16_din1),
        .ap_bram_16_dout1(ap_bram_iarg_16_dout1),
        .ap_bram_16_we1(ap_bram_iarg_16_we1),
        .ap_bram_16_en1(ap_bram_iarg_16_en1),
        .s_axis_bram_17_aclk(s_axis_bram_17_aclk),
        .s_axis_bram_17_aresetn(s_axis_bram_17_aresetn),
        .s_axis_bram_17_tlast(s_axis_bram_17_tlast),
        .s_axis_bram_17_tvalid(s_axis_bram_17_tvalid),
        .s_axis_bram_17_tkeep(s_axis_bram_17_tkeep),
        .s_axis_bram_17_tstrb(s_axis_bram_17_tstrb),
        .s_axis_bram_17_tdata(s_axis_bram_17_tdata),
        .s_axis_bram_17_tready(s_axis_bram_17_tready),
        .ap_bram_17_addr0(ap_bram_iarg_17_addr0),
        .ap_bram_17_din0(ap_bram_iarg_17_din0),
        .ap_bram_17_dout0(ap_bram_iarg_17_dout0),
        .ap_bram_17_we0(ap_bram_iarg_17_we0),
        .ap_bram_17_en0(ap_bram_iarg_17_en0),
        .ap_bram_17_addr1(ap_bram_iarg_17_addr1),
        .ap_bram_17_din1(ap_bram_iarg_17_din1),
        .ap_bram_17_dout1(ap_bram_iarg_17_dout1),
        .ap_bram_17_we1(ap_bram_iarg_17_we1),
        .ap_bram_17_en1(ap_bram_iarg_17_en1),
        .s_axis_bram_18_aclk(s_axis_bram_18_aclk),
        .s_axis_bram_18_aresetn(s_axis_bram_18_aresetn),
        .s_axis_bram_18_tlast(s_axis_bram_18_tlast),
        .s_axis_bram_18_tvalid(s_axis_bram_18_tvalid),
        .s_axis_bram_18_tkeep(s_axis_bram_18_tkeep),
        .s_axis_bram_18_tstrb(s_axis_bram_18_tstrb),
        .s_axis_bram_18_tdata(s_axis_bram_18_tdata),
        .s_axis_bram_18_tready(s_axis_bram_18_tready),
        .ap_bram_18_addr0(ap_bram_iarg_18_addr0),
        .ap_bram_18_din0(ap_bram_iarg_18_din0),
        .ap_bram_18_dout0(ap_bram_iarg_18_dout0),
        .ap_bram_18_we0(ap_bram_iarg_18_we0),
        .ap_bram_18_en0(ap_bram_iarg_18_en0),
        .ap_bram_18_addr1(ap_bram_iarg_18_addr1),
        .ap_bram_18_din1(ap_bram_iarg_18_din1),
        .ap_bram_18_dout1(ap_bram_iarg_18_dout1),
        .ap_bram_18_we1(ap_bram_iarg_18_we1),
        .ap_bram_18_en1(ap_bram_iarg_18_en1),
        .s_axis_bram_19_aclk(s_axis_bram_19_aclk),
        .s_axis_bram_19_aresetn(s_axis_bram_19_aresetn),
        .s_axis_bram_19_tlast(s_axis_bram_19_tlast),
        .s_axis_bram_19_tvalid(s_axis_bram_19_tvalid),
        .s_axis_bram_19_tkeep(s_axis_bram_19_tkeep),
        .s_axis_bram_19_tstrb(s_axis_bram_19_tstrb),
        .s_axis_bram_19_tdata(s_axis_bram_19_tdata),
        .s_axis_bram_19_tready(s_axis_bram_19_tready),
        .ap_bram_19_addr0(ap_bram_iarg_19_addr0),
        .ap_bram_19_din0(ap_bram_iarg_19_din0),
        .ap_bram_19_dout0(ap_bram_iarg_19_dout0),
        .ap_bram_19_we0(ap_bram_iarg_19_we0),
        .ap_bram_19_en0(ap_bram_iarg_19_en0),
        .ap_bram_19_addr1(ap_bram_iarg_19_addr1),
        .ap_bram_19_din1(ap_bram_iarg_19_din1),
        .ap_bram_19_dout1(ap_bram_iarg_19_dout1),
        .ap_bram_19_we1(ap_bram_iarg_19_we1),
        .ap_bram_19_en1(ap_bram_iarg_19_en1),
        .s_axis_bram_20_aclk(s_axis_bram_20_aclk),
        .s_axis_bram_20_aresetn(s_axis_bram_20_aresetn),
        .s_axis_bram_20_tlast(s_axis_bram_20_tlast),
        .s_axis_bram_20_tvalid(s_axis_bram_20_tvalid),
        .s_axis_bram_20_tkeep(s_axis_bram_20_tkeep),
        .s_axis_bram_20_tstrb(s_axis_bram_20_tstrb),
        .s_axis_bram_20_tdata(s_axis_bram_20_tdata),
        .s_axis_bram_20_tready(s_axis_bram_20_tready),
        .ap_bram_20_addr0(ap_bram_iarg_20_addr0),
        .ap_bram_20_din0(ap_bram_iarg_20_din0),
        .ap_bram_20_dout0(ap_bram_iarg_20_dout0),
        .ap_bram_20_we0(ap_bram_iarg_20_we0),
        .ap_bram_20_en0(ap_bram_iarg_20_en0),
        .ap_bram_20_addr1(ap_bram_iarg_20_addr1),
        .ap_bram_20_din1(ap_bram_iarg_20_din1),
        .ap_bram_20_dout1(ap_bram_iarg_20_dout1),
        .ap_bram_20_we1(ap_bram_iarg_20_we1),
        .ap_bram_20_en1(ap_bram_iarg_20_en1),
        .s_axis_bram_21_aclk(s_axis_bram_21_aclk),
        .s_axis_bram_21_aresetn(s_axis_bram_21_aresetn),
        .s_axis_bram_21_tlast(s_axis_bram_21_tlast),
        .s_axis_bram_21_tvalid(s_axis_bram_21_tvalid),
        .s_axis_bram_21_tkeep(s_axis_bram_21_tkeep),
        .s_axis_bram_21_tstrb(s_axis_bram_21_tstrb),
        .s_axis_bram_21_tdata(s_axis_bram_21_tdata),
        .s_axis_bram_21_tready(s_axis_bram_21_tready),
        .ap_bram_21_addr0(ap_bram_iarg_21_addr0),
        .ap_bram_21_din0(ap_bram_iarg_21_din0),
        .ap_bram_21_dout0(ap_bram_iarg_21_dout0),
        .ap_bram_21_we0(ap_bram_iarg_21_we0),
        .ap_bram_21_en0(ap_bram_iarg_21_en0),
        .ap_bram_21_addr1(ap_bram_iarg_21_addr1),
        .ap_bram_21_din1(ap_bram_iarg_21_din1),
        .ap_bram_21_dout1(ap_bram_iarg_21_dout1),
        .ap_bram_21_we1(ap_bram_iarg_21_we1),
        .ap_bram_21_en1(ap_bram_iarg_21_en1),
        .s_axis_bram_22_aclk(s_axis_bram_22_aclk),
        .s_axis_bram_22_aresetn(s_axis_bram_22_aresetn),
        .s_axis_bram_22_tlast(s_axis_bram_22_tlast),
        .s_axis_bram_22_tvalid(s_axis_bram_22_tvalid),
        .s_axis_bram_22_tkeep(s_axis_bram_22_tkeep),
        .s_axis_bram_22_tstrb(s_axis_bram_22_tstrb),
        .s_axis_bram_22_tdata(s_axis_bram_22_tdata),
        .s_axis_bram_22_tready(s_axis_bram_22_tready),
        .ap_bram_22_addr0(ap_bram_iarg_22_addr0),
        .ap_bram_22_din0(ap_bram_iarg_22_din0),
        .ap_bram_22_dout0(ap_bram_iarg_22_dout0),
        .ap_bram_22_we0(ap_bram_iarg_22_we0),
        .ap_bram_22_en0(ap_bram_iarg_22_en0),
        .ap_bram_22_addr1(ap_bram_iarg_22_addr1),
        .ap_bram_22_din1(ap_bram_iarg_22_din1),
        .ap_bram_22_dout1(ap_bram_iarg_22_dout1),
        .ap_bram_22_we1(ap_bram_iarg_22_we1),
        .ap_bram_22_en1(ap_bram_iarg_22_en1),
        .s_axis_bram_23_aclk(s_axis_bram_23_aclk),
        .s_axis_bram_23_aresetn(s_axis_bram_23_aresetn),
        .s_axis_bram_23_tlast(s_axis_bram_23_tlast),
        .s_axis_bram_23_tvalid(s_axis_bram_23_tvalid),
        .s_axis_bram_23_tkeep(s_axis_bram_23_tkeep),
        .s_axis_bram_23_tstrb(s_axis_bram_23_tstrb),
        .s_axis_bram_23_tdata(s_axis_bram_23_tdata),
        .s_axis_bram_23_tready(s_axis_bram_23_tready),
        .ap_bram_23_addr0(ap_bram_iarg_23_addr0),
        .ap_bram_23_din0(ap_bram_iarg_23_din0),
        .ap_bram_23_dout0(ap_bram_iarg_23_dout0),
        .ap_bram_23_we0(ap_bram_iarg_23_we0),
        .ap_bram_23_en0(ap_bram_iarg_23_en0),
        .ap_bram_23_addr1(ap_bram_iarg_23_addr1),
        .ap_bram_23_din1(ap_bram_iarg_23_din1),
        .ap_bram_23_dout1(ap_bram_iarg_23_dout1),
        .ap_bram_23_we1(ap_bram_iarg_23_we1),
        .ap_bram_23_en1(ap_bram_iarg_23_en1),
        .s_axis_bram_24_aclk(s_axis_bram_24_aclk),
        .s_axis_bram_24_aresetn(s_axis_bram_24_aresetn),
        .s_axis_bram_24_tlast(s_axis_bram_24_tlast),
        .s_axis_bram_24_tvalid(s_axis_bram_24_tvalid),
        .s_axis_bram_24_tkeep(s_axis_bram_24_tkeep),
        .s_axis_bram_24_tstrb(s_axis_bram_24_tstrb),
        .s_axis_bram_24_tdata(s_axis_bram_24_tdata),
        .s_axis_bram_24_tready(s_axis_bram_24_tready),
        .ap_bram_24_addr0(ap_bram_iarg_24_addr0),
        .ap_bram_24_din0(ap_bram_iarg_24_din0),
        .ap_bram_24_dout0(ap_bram_iarg_24_dout0),
        .ap_bram_24_we0(ap_bram_iarg_24_we0),
        .ap_bram_24_en0(ap_bram_iarg_24_en0),
        .ap_bram_24_addr1(ap_bram_iarg_24_addr1),
        .ap_bram_24_din1(ap_bram_iarg_24_din1),
        .ap_bram_24_dout1(ap_bram_iarg_24_dout1),
        .ap_bram_24_we1(ap_bram_iarg_24_we1),
        .ap_bram_24_en1(ap_bram_iarg_24_en1),
        .s_axis_bram_25_aclk(s_axis_bram_25_aclk),
        .s_axis_bram_25_aresetn(s_axis_bram_25_aresetn),
        .s_axis_bram_25_tlast(s_axis_bram_25_tlast),
        .s_axis_bram_25_tvalid(s_axis_bram_25_tvalid),
        .s_axis_bram_25_tkeep(s_axis_bram_25_tkeep),
        .s_axis_bram_25_tstrb(s_axis_bram_25_tstrb),
        .s_axis_bram_25_tdata(s_axis_bram_25_tdata),
        .s_axis_bram_25_tready(s_axis_bram_25_tready),
        .ap_bram_25_addr0(ap_bram_iarg_25_addr0),
        .ap_bram_25_din0(ap_bram_iarg_25_din0),
        .ap_bram_25_dout0(ap_bram_iarg_25_dout0),
        .ap_bram_25_we0(ap_bram_iarg_25_we0),
        .ap_bram_25_en0(ap_bram_iarg_25_en0),
        .ap_bram_25_addr1(ap_bram_iarg_25_addr1),
        .ap_bram_25_din1(ap_bram_iarg_25_din1),
        .ap_bram_25_dout1(ap_bram_iarg_25_dout1),
        .ap_bram_25_we1(ap_bram_iarg_25_we1),
        .ap_bram_25_en1(ap_bram_iarg_25_en1),
        .s_axis_bram_26_aclk(s_axis_bram_26_aclk),
        .s_axis_bram_26_aresetn(s_axis_bram_26_aresetn),
        .s_axis_bram_26_tlast(s_axis_bram_26_tlast),
        .s_axis_bram_26_tvalid(s_axis_bram_26_tvalid),
        .s_axis_bram_26_tkeep(s_axis_bram_26_tkeep),
        .s_axis_bram_26_tstrb(s_axis_bram_26_tstrb),
        .s_axis_bram_26_tdata(s_axis_bram_26_tdata),
        .s_axis_bram_26_tready(s_axis_bram_26_tready),
        .ap_bram_26_addr0(ap_bram_iarg_26_addr0),
        .ap_bram_26_din0(ap_bram_iarg_26_din0),
        .ap_bram_26_dout0(ap_bram_iarg_26_dout0),
        .ap_bram_26_we0(ap_bram_iarg_26_we0),
        .ap_bram_26_en0(ap_bram_iarg_26_en0),
        .ap_bram_26_addr1(ap_bram_iarg_26_addr1),
        .ap_bram_26_din1(ap_bram_iarg_26_din1),
        .ap_bram_26_dout1(ap_bram_iarg_26_dout1),
        .ap_bram_26_we1(ap_bram_iarg_26_we1),
        .ap_bram_26_en1(ap_bram_iarg_26_en1),
        .s_axis_bram_27_aclk(s_axis_bram_27_aclk),
        .s_axis_bram_27_aresetn(s_axis_bram_27_aresetn),
        .s_axis_bram_27_tlast(s_axis_bram_27_tlast),
        .s_axis_bram_27_tvalid(s_axis_bram_27_tvalid),
        .s_axis_bram_27_tkeep(s_axis_bram_27_tkeep),
        .s_axis_bram_27_tstrb(s_axis_bram_27_tstrb),
        .s_axis_bram_27_tdata(s_axis_bram_27_tdata),
        .s_axis_bram_27_tready(s_axis_bram_27_tready),
        .ap_bram_27_addr0(ap_bram_iarg_27_addr0),
        .ap_bram_27_din0(ap_bram_iarg_27_din0),
        .ap_bram_27_dout0(ap_bram_iarg_27_dout0),
        .ap_bram_27_we0(ap_bram_iarg_27_we0),
        .ap_bram_27_en0(ap_bram_iarg_27_en0),
        .ap_bram_27_addr1(ap_bram_iarg_27_addr1),
        .ap_bram_27_din1(ap_bram_iarg_27_din1),
        .ap_bram_27_dout1(ap_bram_iarg_27_dout1),
        .ap_bram_27_we1(ap_bram_iarg_27_we1),
        .ap_bram_27_en1(ap_bram_iarg_27_en1),
        .s_axis_bram_28_aclk(s_axis_bram_28_aclk),
        .s_axis_bram_28_aresetn(s_axis_bram_28_aresetn),
        .s_axis_bram_28_tlast(s_axis_bram_28_tlast),
        .s_axis_bram_28_tvalid(s_axis_bram_28_tvalid),
        .s_axis_bram_28_tkeep(s_axis_bram_28_tkeep),
        .s_axis_bram_28_tstrb(s_axis_bram_28_tstrb),
        .s_axis_bram_28_tdata(s_axis_bram_28_tdata),
        .s_axis_bram_28_tready(s_axis_bram_28_tready),
        .ap_bram_28_addr0(ap_bram_iarg_28_addr0),
        .ap_bram_28_din0(ap_bram_iarg_28_din0),
        .ap_bram_28_dout0(ap_bram_iarg_28_dout0),
        .ap_bram_28_we0(ap_bram_iarg_28_we0),
        .ap_bram_28_en0(ap_bram_iarg_28_en0),
        .ap_bram_28_addr1(ap_bram_iarg_28_addr1),
        .ap_bram_28_din1(ap_bram_iarg_28_din1),
        .ap_bram_28_dout1(ap_bram_iarg_28_dout1),
        .ap_bram_28_we1(ap_bram_iarg_28_we1),
        .ap_bram_28_en1(ap_bram_iarg_28_en1),
        .s_axis_bram_29_aclk(s_axis_bram_29_aclk),
        .s_axis_bram_29_aresetn(s_axis_bram_29_aresetn),
        .s_axis_bram_29_tlast(s_axis_bram_29_tlast),
        .s_axis_bram_29_tvalid(s_axis_bram_29_tvalid),
        .s_axis_bram_29_tkeep(s_axis_bram_29_tkeep),
        .s_axis_bram_29_tstrb(s_axis_bram_29_tstrb),
        .s_axis_bram_29_tdata(s_axis_bram_29_tdata),
        .s_axis_bram_29_tready(s_axis_bram_29_tready),
        .ap_bram_29_addr0(ap_bram_iarg_29_addr0),
        .ap_bram_29_din0(ap_bram_iarg_29_din0),
        .ap_bram_29_dout0(ap_bram_iarg_29_dout0),
        .ap_bram_29_we0(ap_bram_iarg_29_we0),
        .ap_bram_29_en0(ap_bram_iarg_29_en0),
        .ap_bram_29_addr1(ap_bram_iarg_29_addr1),
        .ap_bram_29_din1(ap_bram_iarg_29_din1),
        .ap_bram_29_dout1(ap_bram_iarg_29_dout1),
        .ap_bram_29_we1(ap_bram_iarg_29_we1),
        .ap_bram_29_en1(ap_bram_iarg_29_en1),
        .s_axis_bram_30_aclk(s_axis_bram_30_aclk),
        .s_axis_bram_30_aresetn(s_axis_bram_30_aresetn),
        .s_axis_bram_30_tlast(s_axis_bram_30_tlast),
        .s_axis_bram_30_tvalid(s_axis_bram_30_tvalid),
        .s_axis_bram_30_tkeep(s_axis_bram_30_tkeep),
        .s_axis_bram_30_tstrb(s_axis_bram_30_tstrb),
        .s_axis_bram_30_tdata(s_axis_bram_30_tdata),
        .s_axis_bram_30_tready(s_axis_bram_30_tready),
        .ap_bram_30_addr0(ap_bram_iarg_30_addr0),
        .ap_bram_30_din0(ap_bram_iarg_30_din0),
        .ap_bram_30_dout0(ap_bram_iarg_30_dout0),
        .ap_bram_30_we0(ap_bram_iarg_30_we0),
        .ap_bram_30_en0(ap_bram_iarg_30_en0),
        .ap_bram_30_addr1(ap_bram_iarg_30_addr1),
        .ap_bram_30_din1(ap_bram_iarg_30_din1),
        .ap_bram_30_dout1(ap_bram_iarg_30_dout1),
        .ap_bram_30_we1(ap_bram_iarg_30_we1),
        .ap_bram_30_en1(ap_bram_iarg_30_en1),
        .s_axis_bram_31_aclk(s_axis_bram_31_aclk),
        .s_axis_bram_31_aresetn(s_axis_bram_31_aresetn),
        .s_axis_bram_31_tlast(s_axis_bram_31_tlast),
        .s_axis_bram_31_tvalid(s_axis_bram_31_tvalid),
        .s_axis_bram_31_tkeep(s_axis_bram_31_tkeep),
        .s_axis_bram_31_tstrb(s_axis_bram_31_tstrb),
        .s_axis_bram_31_tdata(s_axis_bram_31_tdata),
        .s_axis_bram_31_tready(s_axis_bram_31_tready),
        .ap_bram_31_addr0(ap_bram_iarg_31_addr0),
        .ap_bram_31_din0(ap_bram_iarg_31_din0),
        .ap_bram_31_dout0(ap_bram_iarg_31_dout0),
        .ap_bram_31_we0(ap_bram_iarg_31_we0),
        .ap_bram_31_en0(ap_bram_iarg_31_en0),
        .ap_bram_31_addr1(ap_bram_iarg_31_addr1),
        .ap_bram_31_din1(ap_bram_iarg_31_din1),
        .ap_bram_31_dout1(ap_bram_iarg_31_dout1),
        .ap_bram_31_we1(ap_bram_iarg_31_we1),
        .ap_bram_31_en1(ap_bram_iarg_31_en1),
        .s_axis_bram_32_aclk(s_axis_bram_32_aclk),
        .s_axis_bram_32_aresetn(s_axis_bram_32_aresetn),
        .s_axis_bram_32_tlast(s_axis_bram_32_tlast),
        .s_axis_bram_32_tvalid(s_axis_bram_32_tvalid),
        .s_axis_bram_32_tkeep(s_axis_bram_32_tkeep),
        .s_axis_bram_32_tstrb(s_axis_bram_32_tstrb),
        .s_axis_bram_32_tdata(s_axis_bram_32_tdata),
        .s_axis_bram_32_tready(s_axis_bram_32_tready),
        .ap_bram_32_addr0(ap_bram_iarg_32_addr0),
        .ap_bram_32_din0(ap_bram_iarg_32_din0),
        .ap_bram_32_dout0(ap_bram_iarg_32_dout0),
        .ap_bram_32_we0(ap_bram_iarg_32_we0),
        .ap_bram_32_en0(ap_bram_iarg_32_en0),
        .ap_bram_32_addr1(ap_bram_iarg_32_addr1),
        .ap_bram_32_din1(ap_bram_iarg_32_din1),
        .ap_bram_32_dout1(ap_bram_iarg_32_dout1),
        .ap_bram_32_we1(ap_bram_iarg_32_we1),
        .ap_bram_32_en1(ap_bram_iarg_32_en1),
        .s_axis_bram_33_aclk(s_axis_bram_33_aclk),
        .s_axis_bram_33_aresetn(s_axis_bram_33_aresetn),
        .s_axis_bram_33_tlast(s_axis_bram_33_tlast),
        .s_axis_bram_33_tvalid(s_axis_bram_33_tvalid),
        .s_axis_bram_33_tkeep(s_axis_bram_33_tkeep),
        .s_axis_bram_33_tstrb(s_axis_bram_33_tstrb),
        .s_axis_bram_33_tdata(s_axis_bram_33_tdata),
        .s_axis_bram_33_tready(s_axis_bram_33_tready),
        .ap_bram_33_addr0(ap_bram_iarg_33_addr0),
        .ap_bram_33_din0(ap_bram_iarg_33_din0),
        .ap_bram_33_dout0(ap_bram_iarg_33_dout0),
        .ap_bram_33_we0(ap_bram_iarg_33_we0),
        .ap_bram_33_en0(ap_bram_iarg_33_en0),
        .ap_bram_33_addr1(ap_bram_iarg_33_addr1),
        .ap_bram_33_din1(ap_bram_iarg_33_din1),
        .ap_bram_33_dout1(ap_bram_iarg_33_dout1),
        .ap_bram_33_we1(ap_bram_iarg_33_we1),
        .ap_bram_33_en1(ap_bram_iarg_33_en1),
        .s_axis_bram_34_aclk(s_axis_bram_34_aclk),
        .s_axis_bram_34_aresetn(s_axis_bram_34_aresetn),
        .s_axis_bram_34_tlast(s_axis_bram_34_tlast),
        .s_axis_bram_34_tvalid(s_axis_bram_34_tvalid),
        .s_axis_bram_34_tkeep(s_axis_bram_34_tkeep),
        .s_axis_bram_34_tstrb(s_axis_bram_34_tstrb),
        .s_axis_bram_34_tdata(s_axis_bram_34_tdata),
        .s_axis_bram_34_tready(s_axis_bram_34_tready),
        .ap_bram_34_addr0(ap_bram_iarg_34_addr0),
        .ap_bram_34_din0(ap_bram_iarg_34_din0),
        .ap_bram_34_dout0(ap_bram_iarg_34_dout0),
        .ap_bram_34_we0(ap_bram_iarg_34_we0),
        .ap_bram_34_en0(ap_bram_iarg_34_en0),
        .ap_bram_34_addr1(ap_bram_iarg_34_addr1),
        .ap_bram_34_din1(ap_bram_iarg_34_din1),
        .ap_bram_34_dout1(ap_bram_iarg_34_dout1),
        .ap_bram_34_we1(ap_bram_iarg_34_we1),
        .ap_bram_34_en1(ap_bram_iarg_34_en1),
        .s_axis_bram_35_aclk(s_axis_bram_35_aclk),
        .s_axis_bram_35_aresetn(s_axis_bram_35_aresetn),
        .s_axis_bram_35_tlast(s_axis_bram_35_tlast),
        .s_axis_bram_35_tvalid(s_axis_bram_35_tvalid),
        .s_axis_bram_35_tkeep(s_axis_bram_35_tkeep),
        .s_axis_bram_35_tstrb(s_axis_bram_35_tstrb),
        .s_axis_bram_35_tdata(s_axis_bram_35_tdata),
        .s_axis_bram_35_tready(s_axis_bram_35_tready),
        .ap_bram_35_addr0(ap_bram_iarg_35_addr0),
        .ap_bram_35_din0(ap_bram_iarg_35_din0),
        .ap_bram_35_dout0(ap_bram_iarg_35_dout0),
        .ap_bram_35_we0(ap_bram_iarg_35_we0),
        .ap_bram_35_en0(ap_bram_iarg_35_en0),
        .ap_bram_35_addr1(ap_bram_iarg_35_addr1),
        .ap_bram_35_din1(ap_bram_iarg_35_din1),
        .ap_bram_35_dout1(ap_bram_iarg_35_dout1),
        .ap_bram_35_we1(ap_bram_iarg_35_we1),
        .ap_bram_35_en1(ap_bram_iarg_35_en1),
        .s_axis_bram_36_aclk(s_axis_bram_36_aclk),
        .s_axis_bram_36_aresetn(s_axis_bram_36_aresetn),
        .s_axis_bram_36_tlast(s_axis_bram_36_tlast),
        .s_axis_bram_36_tvalid(s_axis_bram_36_tvalid),
        .s_axis_bram_36_tkeep(s_axis_bram_36_tkeep),
        .s_axis_bram_36_tstrb(s_axis_bram_36_tstrb),
        .s_axis_bram_36_tdata(s_axis_bram_36_tdata),
        .s_axis_bram_36_tready(s_axis_bram_36_tready),
        .ap_bram_36_addr0(ap_bram_iarg_36_addr0),
        .ap_bram_36_din0(ap_bram_iarg_36_din0),
        .ap_bram_36_dout0(ap_bram_iarg_36_dout0),
        .ap_bram_36_we0(ap_bram_iarg_36_we0),
        .ap_bram_36_en0(ap_bram_iarg_36_en0),
        .ap_bram_36_addr1(ap_bram_iarg_36_addr1),
        .ap_bram_36_din1(ap_bram_iarg_36_din1),
        .ap_bram_36_dout1(ap_bram_iarg_36_dout1),
        .ap_bram_36_we1(ap_bram_iarg_36_we1),
        .ap_bram_36_en1(ap_bram_iarg_36_en1),
        .s_axis_bram_37_aclk(s_axis_bram_37_aclk),
        .s_axis_bram_37_aresetn(s_axis_bram_37_aresetn),
        .s_axis_bram_37_tlast(s_axis_bram_37_tlast),
        .s_axis_bram_37_tvalid(s_axis_bram_37_tvalid),
        .s_axis_bram_37_tkeep(s_axis_bram_37_tkeep),
        .s_axis_bram_37_tstrb(s_axis_bram_37_tstrb),
        .s_axis_bram_37_tdata(s_axis_bram_37_tdata),
        .s_axis_bram_37_tready(s_axis_bram_37_tready),
        .ap_bram_37_addr0(ap_bram_iarg_37_addr0),
        .ap_bram_37_din0(ap_bram_iarg_37_din0),
        .ap_bram_37_dout0(ap_bram_iarg_37_dout0),
        .ap_bram_37_we0(ap_bram_iarg_37_we0),
        .ap_bram_37_en0(ap_bram_iarg_37_en0),
        .ap_bram_37_addr1(ap_bram_iarg_37_addr1),
        .ap_bram_37_din1(ap_bram_iarg_37_din1),
        .ap_bram_37_dout1(ap_bram_iarg_37_dout1),
        .ap_bram_37_we1(ap_bram_iarg_37_we1),
        .ap_bram_37_en1(ap_bram_iarg_37_en1),
        .s_axis_bram_38_aclk(s_axis_bram_38_aclk),
        .s_axis_bram_38_aresetn(s_axis_bram_38_aresetn),
        .s_axis_bram_38_tlast(s_axis_bram_38_tlast),
        .s_axis_bram_38_tvalid(s_axis_bram_38_tvalid),
        .s_axis_bram_38_tkeep(s_axis_bram_38_tkeep),
        .s_axis_bram_38_tstrb(s_axis_bram_38_tstrb),
        .s_axis_bram_38_tdata(s_axis_bram_38_tdata),
        .s_axis_bram_38_tready(s_axis_bram_38_tready),
        .ap_bram_38_addr0(ap_bram_iarg_38_addr0),
        .ap_bram_38_din0(ap_bram_iarg_38_din0),
        .ap_bram_38_dout0(ap_bram_iarg_38_dout0),
        .ap_bram_38_we0(ap_bram_iarg_38_we0),
        .ap_bram_38_en0(ap_bram_iarg_38_en0),
        .ap_bram_38_addr1(ap_bram_iarg_38_addr1),
        .ap_bram_38_din1(ap_bram_iarg_38_din1),
        .ap_bram_38_dout1(ap_bram_iarg_38_dout1),
        .ap_bram_38_we1(ap_bram_iarg_38_we1),
        .ap_bram_38_en1(ap_bram_iarg_38_en1),
        .s_axis_bram_39_aclk(s_axis_bram_39_aclk),
        .s_axis_bram_39_aresetn(s_axis_bram_39_aresetn),
        .s_axis_bram_39_tlast(s_axis_bram_39_tlast),
        .s_axis_bram_39_tvalid(s_axis_bram_39_tvalid),
        .s_axis_bram_39_tkeep(s_axis_bram_39_tkeep),
        .s_axis_bram_39_tstrb(s_axis_bram_39_tstrb),
        .s_axis_bram_39_tdata(s_axis_bram_39_tdata),
        .s_axis_bram_39_tready(s_axis_bram_39_tready),
        .ap_bram_39_addr0(ap_bram_iarg_39_addr0),
        .ap_bram_39_din0(ap_bram_iarg_39_din0),
        .ap_bram_39_dout0(ap_bram_iarg_39_dout0),
        .ap_bram_39_we0(ap_bram_iarg_39_we0),
        .ap_bram_39_en0(ap_bram_iarg_39_en0),
        .ap_bram_39_addr1(ap_bram_iarg_39_addr1),
        .ap_bram_39_din1(ap_bram_iarg_39_din1),
        .ap_bram_39_dout1(ap_bram_iarg_39_dout1),
        .ap_bram_39_we1(ap_bram_iarg_39_we1),
        .ap_bram_39_en1(ap_bram_iarg_39_en1),
        .s_axis_bram_40_aclk(s_axis_bram_40_aclk),
        .s_axis_bram_40_aresetn(s_axis_bram_40_aresetn),
        .s_axis_bram_40_tlast(s_axis_bram_40_tlast),
        .s_axis_bram_40_tvalid(s_axis_bram_40_tvalid),
        .s_axis_bram_40_tkeep(s_axis_bram_40_tkeep),
        .s_axis_bram_40_tstrb(s_axis_bram_40_tstrb),
        .s_axis_bram_40_tdata(s_axis_bram_40_tdata),
        .s_axis_bram_40_tready(s_axis_bram_40_tready),
        .ap_bram_40_addr0(ap_bram_iarg_40_addr0),
        .ap_bram_40_din0(ap_bram_iarg_40_din0),
        .ap_bram_40_dout0(ap_bram_iarg_40_dout0),
        .ap_bram_40_we0(ap_bram_iarg_40_we0),
        .ap_bram_40_en0(ap_bram_iarg_40_en0),
        .ap_bram_40_addr1(ap_bram_iarg_40_addr1),
        .ap_bram_40_din1(ap_bram_iarg_40_din1),
        .ap_bram_40_dout1(ap_bram_iarg_40_dout1),
        .ap_bram_40_we1(ap_bram_iarg_40_we1),
        .ap_bram_40_en1(ap_bram_iarg_40_en1),
        .s_axis_bram_41_aclk(s_axis_bram_41_aclk),
        .s_axis_bram_41_aresetn(s_axis_bram_41_aresetn),
        .s_axis_bram_41_tlast(s_axis_bram_41_tlast),
        .s_axis_bram_41_tvalid(s_axis_bram_41_tvalid),
        .s_axis_bram_41_tkeep(s_axis_bram_41_tkeep),
        .s_axis_bram_41_tstrb(s_axis_bram_41_tstrb),
        .s_axis_bram_41_tdata(s_axis_bram_41_tdata),
        .s_axis_bram_41_tready(s_axis_bram_41_tready),
        .ap_bram_41_addr0(ap_bram_iarg_41_addr0),
        .ap_bram_41_din0(ap_bram_iarg_41_din0),
        .ap_bram_41_dout0(ap_bram_iarg_41_dout0),
        .ap_bram_41_we0(ap_bram_iarg_41_we0),
        .ap_bram_41_en0(ap_bram_iarg_41_en0),
        .ap_bram_41_addr1(ap_bram_iarg_41_addr1),
        .ap_bram_41_din1(ap_bram_iarg_41_din1),
        .ap_bram_41_dout1(ap_bram_iarg_41_dout1),
        .ap_bram_41_we1(ap_bram_iarg_41_we1),
        .ap_bram_41_en1(ap_bram_iarg_41_en1),
        .s_axis_bram_42_aclk(s_axis_bram_42_aclk),
        .s_axis_bram_42_aresetn(s_axis_bram_42_aresetn),
        .s_axis_bram_42_tlast(s_axis_bram_42_tlast),
        .s_axis_bram_42_tvalid(s_axis_bram_42_tvalid),
        .s_axis_bram_42_tkeep(s_axis_bram_42_tkeep),
        .s_axis_bram_42_tstrb(s_axis_bram_42_tstrb),
        .s_axis_bram_42_tdata(s_axis_bram_42_tdata),
        .s_axis_bram_42_tready(s_axis_bram_42_tready),
        .ap_bram_42_addr0(ap_bram_iarg_42_addr0),
        .ap_bram_42_din0(ap_bram_iarg_42_din0),
        .ap_bram_42_dout0(ap_bram_iarg_42_dout0),
        .ap_bram_42_we0(ap_bram_iarg_42_we0),
        .ap_bram_42_en0(ap_bram_iarg_42_en0),
        .ap_bram_42_addr1(ap_bram_iarg_42_addr1),
        .ap_bram_42_din1(ap_bram_iarg_42_din1),
        .ap_bram_42_dout1(ap_bram_iarg_42_dout1),
        .ap_bram_42_we1(ap_bram_iarg_42_we1),
        .ap_bram_42_en1(ap_bram_iarg_42_en1),
        .s_axis_bram_43_aclk(s_axis_bram_43_aclk),
        .s_axis_bram_43_aresetn(s_axis_bram_43_aresetn),
        .s_axis_bram_43_tlast(s_axis_bram_43_tlast),
        .s_axis_bram_43_tvalid(s_axis_bram_43_tvalid),
        .s_axis_bram_43_tkeep(s_axis_bram_43_tkeep),
        .s_axis_bram_43_tstrb(s_axis_bram_43_tstrb),
        .s_axis_bram_43_tdata(s_axis_bram_43_tdata),
        .s_axis_bram_43_tready(s_axis_bram_43_tready),
        .ap_bram_43_addr0(ap_bram_iarg_43_addr0),
        .ap_bram_43_din0(ap_bram_iarg_43_din0),
        .ap_bram_43_dout0(ap_bram_iarg_43_dout0),
        .ap_bram_43_we0(ap_bram_iarg_43_we0),
        .ap_bram_43_en0(ap_bram_iarg_43_en0),
        .ap_bram_43_addr1(ap_bram_iarg_43_addr1),
        .ap_bram_43_din1(ap_bram_iarg_43_din1),
        .ap_bram_43_dout1(ap_bram_iarg_43_dout1),
        .ap_bram_43_we1(ap_bram_iarg_43_we1),
        .ap_bram_43_en1(ap_bram_iarg_43_en1),
        .s_axis_bram_44_aclk(s_axis_bram_44_aclk),
        .s_axis_bram_44_aresetn(s_axis_bram_44_aresetn),
        .s_axis_bram_44_tlast(s_axis_bram_44_tlast),
        .s_axis_bram_44_tvalid(s_axis_bram_44_tvalid),
        .s_axis_bram_44_tkeep(s_axis_bram_44_tkeep),
        .s_axis_bram_44_tstrb(s_axis_bram_44_tstrb),
        .s_axis_bram_44_tdata(s_axis_bram_44_tdata),
        .s_axis_bram_44_tready(s_axis_bram_44_tready),
        .ap_bram_44_addr0(ap_bram_iarg_44_addr0),
        .ap_bram_44_din0(ap_bram_iarg_44_din0),
        .ap_bram_44_dout0(ap_bram_iarg_44_dout0),
        .ap_bram_44_we0(ap_bram_iarg_44_we0),
        .ap_bram_44_en0(ap_bram_iarg_44_en0),
        .ap_bram_44_addr1(ap_bram_iarg_44_addr1),
        .ap_bram_44_din1(ap_bram_iarg_44_din1),
        .ap_bram_44_dout1(ap_bram_iarg_44_dout1),
        .ap_bram_44_we1(ap_bram_iarg_44_we1),
        .ap_bram_44_en1(ap_bram_iarg_44_en1),
        .s_axis_bram_45_aclk(s_axis_bram_45_aclk),
        .s_axis_bram_45_aresetn(s_axis_bram_45_aresetn),
        .s_axis_bram_45_tlast(s_axis_bram_45_tlast),
        .s_axis_bram_45_tvalid(s_axis_bram_45_tvalid),
        .s_axis_bram_45_tkeep(s_axis_bram_45_tkeep),
        .s_axis_bram_45_tstrb(s_axis_bram_45_tstrb),
        .s_axis_bram_45_tdata(s_axis_bram_45_tdata),
        .s_axis_bram_45_tready(s_axis_bram_45_tready),
        .ap_bram_45_addr0(ap_bram_iarg_45_addr0),
        .ap_bram_45_din0(ap_bram_iarg_45_din0),
        .ap_bram_45_dout0(ap_bram_iarg_45_dout0),
        .ap_bram_45_we0(ap_bram_iarg_45_we0),
        .ap_bram_45_en0(ap_bram_iarg_45_en0),
        .ap_bram_45_addr1(ap_bram_iarg_45_addr1),
        .ap_bram_45_din1(ap_bram_iarg_45_din1),
        .ap_bram_45_dout1(ap_bram_iarg_45_dout1),
        .ap_bram_45_we1(ap_bram_iarg_45_we1),
        .ap_bram_45_en1(ap_bram_iarg_45_en1),
        .s_axis_bram_46_aclk(s_axis_bram_46_aclk),
        .s_axis_bram_46_aresetn(s_axis_bram_46_aresetn),
        .s_axis_bram_46_tlast(s_axis_bram_46_tlast),
        .s_axis_bram_46_tvalid(s_axis_bram_46_tvalid),
        .s_axis_bram_46_tkeep(s_axis_bram_46_tkeep),
        .s_axis_bram_46_tstrb(s_axis_bram_46_tstrb),
        .s_axis_bram_46_tdata(s_axis_bram_46_tdata),
        .s_axis_bram_46_tready(s_axis_bram_46_tready),
        .ap_bram_46_addr0(ap_bram_iarg_46_addr0),
        .ap_bram_46_din0(ap_bram_iarg_46_din0),
        .ap_bram_46_dout0(ap_bram_iarg_46_dout0),
        .ap_bram_46_we0(ap_bram_iarg_46_we0),
        .ap_bram_46_en0(ap_bram_iarg_46_en0),
        .ap_bram_46_addr1(ap_bram_iarg_46_addr1),
        .ap_bram_46_din1(ap_bram_iarg_46_din1),
        .ap_bram_46_dout1(ap_bram_iarg_46_dout1),
        .ap_bram_46_we1(ap_bram_iarg_46_we1),
        .ap_bram_46_en1(ap_bram_iarg_46_en1),
        .s_axis_bram_47_aclk(s_axis_bram_47_aclk),
        .s_axis_bram_47_aresetn(s_axis_bram_47_aresetn),
        .s_axis_bram_47_tlast(s_axis_bram_47_tlast),
        .s_axis_bram_47_tvalid(s_axis_bram_47_tvalid),
        .s_axis_bram_47_tkeep(s_axis_bram_47_tkeep),
        .s_axis_bram_47_tstrb(s_axis_bram_47_tstrb),
        .s_axis_bram_47_tdata(s_axis_bram_47_tdata),
        .s_axis_bram_47_tready(s_axis_bram_47_tready),
        .ap_bram_47_addr0(ap_bram_iarg_47_addr0),
        .ap_bram_47_din0(ap_bram_iarg_47_din0),
        .ap_bram_47_dout0(ap_bram_iarg_47_dout0),
        .ap_bram_47_we0(ap_bram_iarg_47_we0),
        .ap_bram_47_en0(ap_bram_iarg_47_en0),
        .ap_bram_47_addr1(ap_bram_iarg_47_addr1),
        .ap_bram_47_din1(ap_bram_iarg_47_din1),
        .ap_bram_47_dout1(ap_bram_iarg_47_dout1),
        .ap_bram_47_we1(ap_bram_iarg_47_we1),
        .ap_bram_47_en1(ap_bram_iarg_47_en1),
        .s_axis_bram_48_aclk(s_axis_bram_48_aclk),
        .s_axis_bram_48_aresetn(s_axis_bram_48_aresetn),
        .s_axis_bram_48_tlast(s_axis_bram_48_tlast),
        .s_axis_bram_48_tvalid(s_axis_bram_48_tvalid),
        .s_axis_bram_48_tkeep(s_axis_bram_48_tkeep),
        .s_axis_bram_48_tstrb(s_axis_bram_48_tstrb),
        .s_axis_bram_48_tdata(s_axis_bram_48_tdata),
        .s_axis_bram_48_tready(s_axis_bram_48_tready),
        .ap_bram_48_addr0(ap_bram_iarg_48_addr0),
        .ap_bram_48_din0(ap_bram_iarg_48_din0),
        .ap_bram_48_dout0(ap_bram_iarg_48_dout0),
        .ap_bram_48_we0(ap_bram_iarg_48_we0),
        .ap_bram_48_en0(ap_bram_iarg_48_en0),
        .ap_bram_48_addr1(ap_bram_iarg_48_addr1),
        .ap_bram_48_din1(ap_bram_iarg_48_din1),
        .ap_bram_48_dout1(ap_bram_iarg_48_dout1),
        .ap_bram_48_we1(ap_bram_iarg_48_we1),
        .ap_bram_48_en1(ap_bram_iarg_48_en1),
        .s_axis_bram_49_aclk(s_axis_bram_49_aclk),
        .s_axis_bram_49_aresetn(s_axis_bram_49_aresetn),
        .s_axis_bram_49_tlast(s_axis_bram_49_tlast),
        .s_axis_bram_49_tvalid(s_axis_bram_49_tvalid),
        .s_axis_bram_49_tkeep(s_axis_bram_49_tkeep),
        .s_axis_bram_49_tstrb(s_axis_bram_49_tstrb),
        .s_axis_bram_49_tdata(s_axis_bram_49_tdata),
        .s_axis_bram_49_tready(s_axis_bram_49_tready),
        .ap_bram_49_addr0(ap_bram_iarg_49_addr0),
        .ap_bram_49_din0(ap_bram_iarg_49_din0),
        .ap_bram_49_dout0(ap_bram_iarg_49_dout0),
        .ap_bram_49_we0(ap_bram_iarg_49_we0),
        .ap_bram_49_en0(ap_bram_iarg_49_en0),
        .ap_bram_49_addr1(ap_bram_iarg_49_addr1),
        .ap_bram_49_din1(ap_bram_iarg_49_din1),
        .ap_bram_49_dout1(ap_bram_iarg_49_dout1),
        .ap_bram_49_we1(ap_bram_iarg_49_we1),
        .ap_bram_49_en1(ap_bram_iarg_49_en1),
        .s_axis_bram_50_aclk(s_axis_bram_50_aclk),
        .s_axis_bram_50_aresetn(s_axis_bram_50_aresetn),
        .s_axis_bram_50_tlast(s_axis_bram_50_tlast),
        .s_axis_bram_50_tvalid(s_axis_bram_50_tvalid),
        .s_axis_bram_50_tkeep(s_axis_bram_50_tkeep),
        .s_axis_bram_50_tstrb(s_axis_bram_50_tstrb),
        .s_axis_bram_50_tdata(s_axis_bram_50_tdata),
        .s_axis_bram_50_tready(s_axis_bram_50_tready),
        .ap_bram_50_addr0(ap_bram_iarg_50_addr0),
        .ap_bram_50_din0(ap_bram_iarg_50_din0),
        .ap_bram_50_dout0(ap_bram_iarg_50_dout0),
        .ap_bram_50_we0(ap_bram_iarg_50_we0),
        .ap_bram_50_en0(ap_bram_iarg_50_en0),
        .ap_bram_50_addr1(ap_bram_iarg_50_addr1),
        .ap_bram_50_din1(ap_bram_iarg_50_din1),
        .ap_bram_50_dout1(ap_bram_iarg_50_dout1),
        .ap_bram_50_we1(ap_bram_iarg_50_we1),
        .ap_bram_50_en1(ap_bram_iarg_50_en1),
        .s_axis_bram_51_aclk(s_axis_bram_51_aclk),
        .s_axis_bram_51_aresetn(s_axis_bram_51_aresetn),
        .s_axis_bram_51_tlast(s_axis_bram_51_tlast),
        .s_axis_bram_51_tvalid(s_axis_bram_51_tvalid),
        .s_axis_bram_51_tkeep(s_axis_bram_51_tkeep),
        .s_axis_bram_51_tstrb(s_axis_bram_51_tstrb),
        .s_axis_bram_51_tdata(s_axis_bram_51_tdata),
        .s_axis_bram_51_tready(s_axis_bram_51_tready),
        .ap_bram_51_addr0(ap_bram_iarg_51_addr0),
        .ap_bram_51_din0(ap_bram_iarg_51_din0),
        .ap_bram_51_dout0(ap_bram_iarg_51_dout0),
        .ap_bram_51_we0(ap_bram_iarg_51_we0),
        .ap_bram_51_en0(ap_bram_iarg_51_en0),
        .ap_bram_51_addr1(ap_bram_iarg_51_addr1),
        .ap_bram_51_din1(ap_bram_iarg_51_din1),
        .ap_bram_51_dout1(ap_bram_iarg_51_dout1),
        .ap_bram_51_we1(ap_bram_iarg_51_we1),
        .ap_bram_51_en1(ap_bram_iarg_51_en1),
        .s_axis_bram_52_aclk(s_axis_bram_52_aclk),
        .s_axis_bram_52_aresetn(s_axis_bram_52_aresetn),
        .s_axis_bram_52_tlast(s_axis_bram_52_tlast),
        .s_axis_bram_52_tvalid(s_axis_bram_52_tvalid),
        .s_axis_bram_52_tkeep(s_axis_bram_52_tkeep),
        .s_axis_bram_52_tstrb(s_axis_bram_52_tstrb),
        .s_axis_bram_52_tdata(s_axis_bram_52_tdata),
        .s_axis_bram_52_tready(s_axis_bram_52_tready),
        .ap_bram_52_addr0(ap_bram_iarg_52_addr0),
        .ap_bram_52_din0(ap_bram_iarg_52_din0),
        .ap_bram_52_dout0(ap_bram_iarg_52_dout0),
        .ap_bram_52_we0(ap_bram_iarg_52_we0),
        .ap_bram_52_en0(ap_bram_iarg_52_en0),
        .ap_bram_52_addr1(ap_bram_iarg_52_addr1),
        .ap_bram_52_din1(ap_bram_iarg_52_din1),
        .ap_bram_52_dout1(ap_bram_iarg_52_dout1),
        .ap_bram_52_we1(ap_bram_iarg_52_we1),
        .ap_bram_52_en1(ap_bram_iarg_52_en1),
        .s_axis_bram_53_aclk(s_axis_bram_53_aclk),
        .s_axis_bram_53_aresetn(s_axis_bram_53_aresetn),
        .s_axis_bram_53_tlast(s_axis_bram_53_tlast),
        .s_axis_bram_53_tvalid(s_axis_bram_53_tvalid),
        .s_axis_bram_53_tkeep(s_axis_bram_53_tkeep),
        .s_axis_bram_53_tstrb(s_axis_bram_53_tstrb),
        .s_axis_bram_53_tdata(s_axis_bram_53_tdata),
        .s_axis_bram_53_tready(s_axis_bram_53_tready),
        .ap_bram_53_addr0(ap_bram_iarg_53_addr0),
        .ap_bram_53_din0(ap_bram_iarg_53_din0),
        .ap_bram_53_dout0(ap_bram_iarg_53_dout0),
        .ap_bram_53_we0(ap_bram_iarg_53_we0),
        .ap_bram_53_en0(ap_bram_iarg_53_en0),
        .ap_bram_53_addr1(ap_bram_iarg_53_addr1),
        .ap_bram_53_din1(ap_bram_iarg_53_din1),
        .ap_bram_53_dout1(ap_bram_iarg_53_dout1),
        .ap_bram_53_we1(ap_bram_iarg_53_we1),
        .ap_bram_53_en1(ap_bram_iarg_53_en1),
        .s_axis_bram_54_aclk(s_axis_bram_54_aclk),
        .s_axis_bram_54_aresetn(s_axis_bram_54_aresetn),
        .s_axis_bram_54_tlast(s_axis_bram_54_tlast),
        .s_axis_bram_54_tvalid(s_axis_bram_54_tvalid),
        .s_axis_bram_54_tkeep(s_axis_bram_54_tkeep),
        .s_axis_bram_54_tstrb(s_axis_bram_54_tstrb),
        .s_axis_bram_54_tdata(s_axis_bram_54_tdata),
        .s_axis_bram_54_tready(s_axis_bram_54_tready),
        .ap_bram_54_addr0(ap_bram_iarg_54_addr0),
        .ap_bram_54_din0(ap_bram_iarg_54_din0),
        .ap_bram_54_dout0(ap_bram_iarg_54_dout0),
        .ap_bram_54_we0(ap_bram_iarg_54_we0),
        .ap_bram_54_en0(ap_bram_iarg_54_en0),
        .ap_bram_54_addr1(ap_bram_iarg_54_addr1),
        .ap_bram_54_din1(ap_bram_iarg_54_din1),
        .ap_bram_54_dout1(ap_bram_iarg_54_dout1),
        .ap_bram_54_we1(ap_bram_iarg_54_we1),
        .ap_bram_54_en1(ap_bram_iarg_54_en1),
        .s_axis_bram_55_aclk(s_axis_bram_55_aclk),
        .s_axis_bram_55_aresetn(s_axis_bram_55_aresetn),
        .s_axis_bram_55_tlast(s_axis_bram_55_tlast),
        .s_axis_bram_55_tvalid(s_axis_bram_55_tvalid),
        .s_axis_bram_55_tkeep(s_axis_bram_55_tkeep),
        .s_axis_bram_55_tstrb(s_axis_bram_55_tstrb),
        .s_axis_bram_55_tdata(s_axis_bram_55_tdata),
        .s_axis_bram_55_tready(s_axis_bram_55_tready),
        .ap_bram_55_addr0(ap_bram_iarg_55_addr0),
        .ap_bram_55_din0(ap_bram_iarg_55_din0),
        .ap_bram_55_dout0(ap_bram_iarg_55_dout0),
        .ap_bram_55_we0(ap_bram_iarg_55_we0),
        .ap_bram_55_en0(ap_bram_iarg_55_en0),
        .ap_bram_55_addr1(ap_bram_iarg_55_addr1),
        .ap_bram_55_din1(ap_bram_iarg_55_din1),
        .ap_bram_55_dout1(ap_bram_iarg_55_dout1),
        .ap_bram_55_we1(ap_bram_iarg_55_we1),
        .ap_bram_55_en1(ap_bram_iarg_55_en1),
        .s_axis_bram_56_aclk(s_axis_bram_56_aclk),
        .s_axis_bram_56_aresetn(s_axis_bram_56_aresetn),
        .s_axis_bram_56_tlast(s_axis_bram_56_tlast),
        .s_axis_bram_56_tvalid(s_axis_bram_56_tvalid),
        .s_axis_bram_56_tkeep(s_axis_bram_56_tkeep),
        .s_axis_bram_56_tstrb(s_axis_bram_56_tstrb),
        .s_axis_bram_56_tdata(s_axis_bram_56_tdata),
        .s_axis_bram_56_tready(s_axis_bram_56_tready),
        .ap_bram_56_addr0(ap_bram_iarg_56_addr0),
        .ap_bram_56_din0(ap_bram_iarg_56_din0),
        .ap_bram_56_dout0(ap_bram_iarg_56_dout0),
        .ap_bram_56_we0(ap_bram_iarg_56_we0),
        .ap_bram_56_en0(ap_bram_iarg_56_en0),
        .ap_bram_56_addr1(ap_bram_iarg_56_addr1),
        .ap_bram_56_din1(ap_bram_iarg_56_din1),
        .ap_bram_56_dout1(ap_bram_iarg_56_dout1),
        .ap_bram_56_we1(ap_bram_iarg_56_we1),
        .ap_bram_56_en1(ap_bram_iarg_56_en1),
        .s_axis_bram_57_aclk(s_axis_bram_57_aclk),
        .s_axis_bram_57_aresetn(s_axis_bram_57_aresetn),
        .s_axis_bram_57_tlast(s_axis_bram_57_tlast),
        .s_axis_bram_57_tvalid(s_axis_bram_57_tvalid),
        .s_axis_bram_57_tkeep(s_axis_bram_57_tkeep),
        .s_axis_bram_57_tstrb(s_axis_bram_57_tstrb),
        .s_axis_bram_57_tdata(s_axis_bram_57_tdata),
        .s_axis_bram_57_tready(s_axis_bram_57_tready),
        .ap_bram_57_addr0(ap_bram_iarg_57_addr0),
        .ap_bram_57_din0(ap_bram_iarg_57_din0),
        .ap_bram_57_dout0(ap_bram_iarg_57_dout0),
        .ap_bram_57_we0(ap_bram_iarg_57_we0),
        .ap_bram_57_en0(ap_bram_iarg_57_en0),
        .ap_bram_57_addr1(ap_bram_iarg_57_addr1),
        .ap_bram_57_din1(ap_bram_iarg_57_din1),
        .ap_bram_57_dout1(ap_bram_iarg_57_dout1),
        .ap_bram_57_we1(ap_bram_iarg_57_we1),
        .ap_bram_57_en1(ap_bram_iarg_57_en1),
        .s_axis_bram_58_aclk(s_axis_bram_58_aclk),
        .s_axis_bram_58_aresetn(s_axis_bram_58_aresetn),
        .s_axis_bram_58_tlast(s_axis_bram_58_tlast),
        .s_axis_bram_58_tvalid(s_axis_bram_58_tvalid),
        .s_axis_bram_58_tkeep(s_axis_bram_58_tkeep),
        .s_axis_bram_58_tstrb(s_axis_bram_58_tstrb),
        .s_axis_bram_58_tdata(s_axis_bram_58_tdata),
        .s_axis_bram_58_tready(s_axis_bram_58_tready),
        .ap_bram_58_addr0(ap_bram_iarg_58_addr0),
        .ap_bram_58_din0(ap_bram_iarg_58_din0),
        .ap_bram_58_dout0(ap_bram_iarg_58_dout0),
        .ap_bram_58_we0(ap_bram_iarg_58_we0),
        .ap_bram_58_en0(ap_bram_iarg_58_en0),
        .ap_bram_58_addr1(ap_bram_iarg_58_addr1),
        .ap_bram_58_din1(ap_bram_iarg_58_din1),
        .ap_bram_58_dout1(ap_bram_iarg_58_dout1),
        .ap_bram_58_we1(ap_bram_iarg_58_we1),
        .ap_bram_58_en1(ap_bram_iarg_58_en1),
        .s_axis_bram_59_aclk(s_axis_bram_59_aclk),
        .s_axis_bram_59_aresetn(s_axis_bram_59_aresetn),
        .s_axis_bram_59_tlast(s_axis_bram_59_tlast),
        .s_axis_bram_59_tvalid(s_axis_bram_59_tvalid),
        .s_axis_bram_59_tkeep(s_axis_bram_59_tkeep),
        .s_axis_bram_59_tstrb(s_axis_bram_59_tstrb),
        .s_axis_bram_59_tdata(s_axis_bram_59_tdata),
        .s_axis_bram_59_tready(s_axis_bram_59_tready),
        .ap_bram_59_addr0(ap_bram_iarg_59_addr0),
        .ap_bram_59_din0(ap_bram_iarg_59_din0),
        .ap_bram_59_dout0(ap_bram_iarg_59_dout0),
        .ap_bram_59_we0(ap_bram_iarg_59_we0),
        .ap_bram_59_en0(ap_bram_iarg_59_en0),
        .ap_bram_59_addr1(ap_bram_iarg_59_addr1),
        .ap_bram_59_din1(ap_bram_iarg_59_din1),
        .ap_bram_59_dout1(ap_bram_iarg_59_dout1),
        .ap_bram_59_we1(ap_bram_iarg_59_we1),
        .ap_bram_59_en1(ap_bram_iarg_59_en1),
        .s_axis_bram_60_aclk(s_axis_bram_60_aclk),
        .s_axis_bram_60_aresetn(s_axis_bram_60_aresetn),
        .s_axis_bram_60_tlast(s_axis_bram_60_tlast),
        .s_axis_bram_60_tvalid(s_axis_bram_60_tvalid),
        .s_axis_bram_60_tkeep(s_axis_bram_60_tkeep),
        .s_axis_bram_60_tstrb(s_axis_bram_60_tstrb),
        .s_axis_bram_60_tdata(s_axis_bram_60_tdata),
        .s_axis_bram_60_tready(s_axis_bram_60_tready),
        .ap_bram_60_addr0(ap_bram_iarg_60_addr0),
        .ap_bram_60_din0(ap_bram_iarg_60_din0),
        .ap_bram_60_dout0(ap_bram_iarg_60_dout0),
        .ap_bram_60_we0(ap_bram_iarg_60_we0),
        .ap_bram_60_en0(ap_bram_iarg_60_en0),
        .ap_bram_60_addr1(ap_bram_iarg_60_addr1),
        .ap_bram_60_din1(ap_bram_iarg_60_din1),
        .ap_bram_60_dout1(ap_bram_iarg_60_dout1),
        .ap_bram_60_we1(ap_bram_iarg_60_we1),
        .ap_bram_60_en1(ap_bram_iarg_60_en1),
        .s_axis_bram_61_aclk(s_axis_bram_61_aclk),
        .s_axis_bram_61_aresetn(s_axis_bram_61_aresetn),
        .s_axis_bram_61_tlast(s_axis_bram_61_tlast),
        .s_axis_bram_61_tvalid(s_axis_bram_61_tvalid),
        .s_axis_bram_61_tkeep(s_axis_bram_61_tkeep),
        .s_axis_bram_61_tstrb(s_axis_bram_61_tstrb),
        .s_axis_bram_61_tdata(s_axis_bram_61_tdata),
        .s_axis_bram_61_tready(s_axis_bram_61_tready),
        .ap_bram_61_addr0(ap_bram_iarg_61_addr0),
        .ap_bram_61_din0(ap_bram_iarg_61_din0),
        .ap_bram_61_dout0(ap_bram_iarg_61_dout0),
        .ap_bram_61_we0(ap_bram_iarg_61_we0),
        .ap_bram_61_en0(ap_bram_iarg_61_en0),
        .ap_bram_61_addr1(ap_bram_iarg_61_addr1),
        .ap_bram_61_din1(ap_bram_iarg_61_din1),
        .ap_bram_61_dout1(ap_bram_iarg_61_dout1),
        .ap_bram_61_we1(ap_bram_iarg_61_we1),
        .ap_bram_61_en1(ap_bram_iarg_61_en1),
        .s_axis_bram_62_aclk(s_axis_bram_62_aclk),
        .s_axis_bram_62_aresetn(s_axis_bram_62_aresetn),
        .s_axis_bram_62_tlast(s_axis_bram_62_tlast),
        .s_axis_bram_62_tvalid(s_axis_bram_62_tvalid),
        .s_axis_bram_62_tkeep(s_axis_bram_62_tkeep),
        .s_axis_bram_62_tstrb(s_axis_bram_62_tstrb),
        .s_axis_bram_62_tdata(s_axis_bram_62_tdata),
        .s_axis_bram_62_tready(s_axis_bram_62_tready),
        .ap_bram_62_addr0(ap_bram_iarg_62_addr0),
        .ap_bram_62_din0(ap_bram_iarg_62_din0),
        .ap_bram_62_dout0(ap_bram_iarg_62_dout0),
        .ap_bram_62_we0(ap_bram_iarg_62_we0),
        .ap_bram_62_en0(ap_bram_iarg_62_en0),
        .ap_bram_62_addr1(ap_bram_iarg_62_addr1),
        .ap_bram_62_din1(ap_bram_iarg_62_din1),
        .ap_bram_62_dout1(ap_bram_iarg_62_dout1),
        .ap_bram_62_we1(ap_bram_iarg_62_we1),
        .ap_bram_62_en1(ap_bram_iarg_62_en1),
        .s_axis_bram_63_aclk(s_axis_bram_63_aclk),
        .s_axis_bram_63_aresetn(s_axis_bram_63_aresetn),
        .s_axis_bram_63_tlast(s_axis_bram_63_tlast),
        .s_axis_bram_63_tvalid(s_axis_bram_63_tvalid),
        .s_axis_bram_63_tkeep(s_axis_bram_63_tkeep),
        .s_axis_bram_63_tstrb(s_axis_bram_63_tstrb),
        .s_axis_bram_63_tdata(s_axis_bram_63_tdata),
        .s_axis_bram_63_tready(s_axis_bram_63_tready),
        .ap_bram_63_addr0(ap_bram_iarg_63_addr0),
        .ap_bram_63_din0(ap_bram_iarg_63_din0),
        .ap_bram_63_dout0(ap_bram_iarg_63_dout0),
        .ap_bram_63_we0(ap_bram_iarg_63_we0),
        .ap_bram_63_en0(ap_bram_iarg_63_en0),
        .ap_bram_63_addr1(ap_bram_iarg_63_addr1),
        .ap_bram_63_din1(ap_bram_iarg_63_din1),
        .ap_bram_63_dout1(ap_bram_iarg_63_dout1),
        .ap_bram_63_we1(ap_bram_iarg_63_we1),
        .ap_bram_63_en1(ap_bram_iarg_63_en1),
        .s_axis_bram_64_aclk(s_axis_bram_64_aclk),
        .s_axis_bram_64_aresetn(s_axis_bram_64_aresetn),
        .s_axis_bram_64_tlast(s_axis_bram_64_tlast),
        .s_axis_bram_64_tvalid(s_axis_bram_64_tvalid),
        .s_axis_bram_64_tkeep(s_axis_bram_64_tkeep),
        .s_axis_bram_64_tstrb(s_axis_bram_64_tstrb),
        .s_axis_bram_64_tdata(s_axis_bram_64_tdata),
        .s_axis_bram_64_tready(s_axis_bram_64_tready),
        .ap_bram_64_addr0(ap_bram_iarg_64_addr0),
        .ap_bram_64_din0(ap_bram_iarg_64_din0),
        .ap_bram_64_dout0(ap_bram_iarg_64_dout0),
        .ap_bram_64_we0(ap_bram_iarg_64_we0),
        .ap_bram_64_en0(ap_bram_iarg_64_en0),
        .ap_bram_64_addr1(ap_bram_iarg_64_addr1),
        .ap_bram_64_din1(ap_bram_iarg_64_din1),
        .ap_bram_64_dout1(ap_bram_iarg_64_dout1),
        .ap_bram_64_we1(ap_bram_iarg_64_we1),
        .ap_bram_64_en1(ap_bram_iarg_64_en1),
        .s_axis_bram_65_aclk(s_axis_bram_65_aclk),
        .s_axis_bram_65_aresetn(s_axis_bram_65_aresetn),
        .s_axis_bram_65_tlast(s_axis_bram_65_tlast),
        .s_axis_bram_65_tvalid(s_axis_bram_65_tvalid),
        .s_axis_bram_65_tkeep(s_axis_bram_65_tkeep),
        .s_axis_bram_65_tstrb(s_axis_bram_65_tstrb),
        .s_axis_bram_65_tdata(s_axis_bram_65_tdata),
        .s_axis_bram_65_tready(s_axis_bram_65_tready),
        .ap_bram_65_addr0(ap_bram_iarg_65_addr0),
        .ap_bram_65_din0(ap_bram_iarg_65_din0),
        .ap_bram_65_dout0(ap_bram_iarg_65_dout0),
        .ap_bram_65_we0(ap_bram_iarg_65_we0),
        .ap_bram_65_en0(ap_bram_iarg_65_en0),
        .ap_bram_65_addr1(ap_bram_iarg_65_addr1),
        .ap_bram_65_din1(ap_bram_iarg_65_din1),
        .ap_bram_65_dout1(ap_bram_iarg_65_dout1),
        .ap_bram_65_we1(ap_bram_iarg_65_we1),
        .ap_bram_65_en1(ap_bram_iarg_65_en1),
        .s_axis_bram_66_aclk(s_axis_bram_66_aclk),
        .s_axis_bram_66_aresetn(s_axis_bram_66_aresetn),
        .s_axis_bram_66_tlast(s_axis_bram_66_tlast),
        .s_axis_bram_66_tvalid(s_axis_bram_66_tvalid),
        .s_axis_bram_66_tkeep(s_axis_bram_66_tkeep),
        .s_axis_bram_66_tstrb(s_axis_bram_66_tstrb),
        .s_axis_bram_66_tdata(s_axis_bram_66_tdata),
        .s_axis_bram_66_tready(s_axis_bram_66_tready),
        .ap_bram_66_addr0(ap_bram_iarg_66_addr0),
        .ap_bram_66_din0(ap_bram_iarg_66_din0),
        .ap_bram_66_dout0(ap_bram_iarg_66_dout0),
        .ap_bram_66_we0(ap_bram_iarg_66_we0),
        .ap_bram_66_en0(ap_bram_iarg_66_en0),
        .ap_bram_66_addr1(ap_bram_iarg_66_addr1),
        .ap_bram_66_din1(ap_bram_iarg_66_din1),
        .ap_bram_66_dout1(ap_bram_iarg_66_dout1),
        .ap_bram_66_we1(ap_bram_iarg_66_we1),
        .ap_bram_66_en1(ap_bram_iarg_66_en1),
        .s_axis_bram_67_aclk(s_axis_bram_67_aclk),
        .s_axis_bram_67_aresetn(s_axis_bram_67_aresetn),
        .s_axis_bram_67_tlast(s_axis_bram_67_tlast),
        .s_axis_bram_67_tvalid(s_axis_bram_67_tvalid),
        .s_axis_bram_67_tkeep(s_axis_bram_67_tkeep),
        .s_axis_bram_67_tstrb(s_axis_bram_67_tstrb),
        .s_axis_bram_67_tdata(s_axis_bram_67_tdata),
        .s_axis_bram_67_tready(s_axis_bram_67_tready),
        .ap_bram_67_addr0(ap_bram_iarg_67_addr0),
        .ap_bram_67_din0(ap_bram_iarg_67_din0),
        .ap_bram_67_dout0(ap_bram_iarg_67_dout0),
        .ap_bram_67_we0(ap_bram_iarg_67_we0),
        .ap_bram_67_en0(ap_bram_iarg_67_en0),
        .ap_bram_67_addr1(ap_bram_iarg_67_addr1),
        .ap_bram_67_din1(ap_bram_iarg_67_din1),
        .ap_bram_67_dout1(ap_bram_iarg_67_dout1),
        .ap_bram_67_we1(ap_bram_iarg_67_we1),
        .ap_bram_67_en1(ap_bram_iarg_67_en1),
        .s_axis_bram_68_aclk(s_axis_bram_68_aclk),
        .s_axis_bram_68_aresetn(s_axis_bram_68_aresetn),
        .s_axis_bram_68_tlast(s_axis_bram_68_tlast),
        .s_axis_bram_68_tvalid(s_axis_bram_68_tvalid),
        .s_axis_bram_68_tkeep(s_axis_bram_68_tkeep),
        .s_axis_bram_68_tstrb(s_axis_bram_68_tstrb),
        .s_axis_bram_68_tdata(s_axis_bram_68_tdata),
        .s_axis_bram_68_tready(s_axis_bram_68_tready),
        .ap_bram_68_addr0(ap_bram_iarg_68_addr0),
        .ap_bram_68_din0(ap_bram_iarg_68_din0),
        .ap_bram_68_dout0(ap_bram_iarg_68_dout0),
        .ap_bram_68_we0(ap_bram_iarg_68_we0),
        .ap_bram_68_en0(ap_bram_iarg_68_en0),
        .ap_bram_68_addr1(ap_bram_iarg_68_addr1),
        .ap_bram_68_din1(ap_bram_iarg_68_din1),
        .ap_bram_68_dout1(ap_bram_iarg_68_dout1),
        .ap_bram_68_we1(ap_bram_iarg_68_we1),
        .ap_bram_68_en1(ap_bram_iarg_68_en1),
        .s_axis_bram_69_aclk(s_axis_bram_69_aclk),
        .s_axis_bram_69_aresetn(s_axis_bram_69_aresetn),
        .s_axis_bram_69_tlast(s_axis_bram_69_tlast),
        .s_axis_bram_69_tvalid(s_axis_bram_69_tvalid),
        .s_axis_bram_69_tkeep(s_axis_bram_69_tkeep),
        .s_axis_bram_69_tstrb(s_axis_bram_69_tstrb),
        .s_axis_bram_69_tdata(s_axis_bram_69_tdata),
        .s_axis_bram_69_tready(s_axis_bram_69_tready),
        .ap_bram_69_addr0(ap_bram_iarg_69_addr0),
        .ap_bram_69_din0(ap_bram_iarg_69_din0),
        .ap_bram_69_dout0(ap_bram_iarg_69_dout0),
        .ap_bram_69_we0(ap_bram_iarg_69_we0),
        .ap_bram_69_en0(ap_bram_iarg_69_en0),
        .ap_bram_69_addr1(ap_bram_iarg_69_addr1),
        .ap_bram_69_din1(ap_bram_iarg_69_din1),
        .ap_bram_69_dout1(ap_bram_iarg_69_dout1),
        .ap_bram_69_we1(ap_bram_iarg_69_we1),
        .ap_bram_69_en1(ap_bram_iarg_69_en1),
        .s_axis_bram_70_aclk(s_axis_bram_70_aclk),
        .s_axis_bram_70_aresetn(s_axis_bram_70_aresetn),
        .s_axis_bram_70_tlast(s_axis_bram_70_tlast),
        .s_axis_bram_70_tvalid(s_axis_bram_70_tvalid),
        .s_axis_bram_70_tkeep(s_axis_bram_70_tkeep),
        .s_axis_bram_70_tstrb(s_axis_bram_70_tstrb),
        .s_axis_bram_70_tdata(s_axis_bram_70_tdata),
        .s_axis_bram_70_tready(s_axis_bram_70_tready),
        .ap_bram_70_addr0(ap_bram_iarg_70_addr0),
        .ap_bram_70_din0(ap_bram_iarg_70_din0),
        .ap_bram_70_dout0(ap_bram_iarg_70_dout0),
        .ap_bram_70_we0(ap_bram_iarg_70_we0),
        .ap_bram_70_en0(ap_bram_iarg_70_en0),
        .ap_bram_70_addr1(ap_bram_iarg_70_addr1),
        .ap_bram_70_din1(ap_bram_iarg_70_din1),
        .ap_bram_70_dout1(ap_bram_iarg_70_dout1),
        .ap_bram_70_we1(ap_bram_iarg_70_we1),
        .ap_bram_70_en1(ap_bram_iarg_70_en1),
        .s_axis_bram_71_aclk(s_axis_bram_71_aclk),
        .s_axis_bram_71_aresetn(s_axis_bram_71_aresetn),
        .s_axis_bram_71_tlast(s_axis_bram_71_tlast),
        .s_axis_bram_71_tvalid(s_axis_bram_71_tvalid),
        .s_axis_bram_71_tkeep(s_axis_bram_71_tkeep),
        .s_axis_bram_71_tstrb(s_axis_bram_71_tstrb),
        .s_axis_bram_71_tdata(s_axis_bram_71_tdata),
        .s_axis_bram_71_tready(s_axis_bram_71_tready),
        .ap_bram_71_addr0(ap_bram_iarg_71_addr0),
        .ap_bram_71_din0(ap_bram_iarg_71_din0),
        .ap_bram_71_dout0(ap_bram_iarg_71_dout0),
        .ap_bram_71_we0(ap_bram_iarg_71_we0),
        .ap_bram_71_en0(ap_bram_iarg_71_en0),
        .ap_bram_71_addr1(ap_bram_iarg_71_addr1),
        .ap_bram_71_din1(ap_bram_iarg_71_din1),
        .ap_bram_71_dout1(ap_bram_iarg_71_dout1),
        .ap_bram_71_we1(ap_bram_iarg_71_we1),
        .ap_bram_71_en1(ap_bram_iarg_71_en1),
        .s_axis_bram_72_aclk(s_axis_bram_72_aclk),
        .s_axis_bram_72_aresetn(s_axis_bram_72_aresetn),
        .s_axis_bram_72_tlast(s_axis_bram_72_tlast),
        .s_axis_bram_72_tvalid(s_axis_bram_72_tvalid),
        .s_axis_bram_72_tkeep(s_axis_bram_72_tkeep),
        .s_axis_bram_72_tstrb(s_axis_bram_72_tstrb),
        .s_axis_bram_72_tdata(s_axis_bram_72_tdata),
        .s_axis_bram_72_tready(s_axis_bram_72_tready),
        .ap_bram_72_addr0(ap_bram_iarg_72_addr0),
        .ap_bram_72_din0(ap_bram_iarg_72_din0),
        .ap_bram_72_dout0(ap_bram_iarg_72_dout0),
        .ap_bram_72_we0(ap_bram_iarg_72_we0),
        .ap_bram_72_en0(ap_bram_iarg_72_en0),
        .ap_bram_72_addr1(ap_bram_iarg_72_addr1),
        .ap_bram_72_din1(ap_bram_iarg_72_din1),
        .ap_bram_72_dout1(ap_bram_iarg_72_dout1),
        .ap_bram_72_we1(ap_bram_iarg_72_we1),
        .ap_bram_72_en1(ap_bram_iarg_72_en1),
        .s_axis_bram_73_aclk(s_axis_bram_73_aclk),
        .s_axis_bram_73_aresetn(s_axis_bram_73_aresetn),
        .s_axis_bram_73_tlast(s_axis_bram_73_tlast),
        .s_axis_bram_73_tvalid(s_axis_bram_73_tvalid),
        .s_axis_bram_73_tkeep(s_axis_bram_73_tkeep),
        .s_axis_bram_73_tstrb(s_axis_bram_73_tstrb),
        .s_axis_bram_73_tdata(s_axis_bram_73_tdata),
        .s_axis_bram_73_tready(s_axis_bram_73_tready),
        .ap_bram_73_addr0(ap_bram_iarg_73_addr0),
        .ap_bram_73_din0(ap_bram_iarg_73_din0),
        .ap_bram_73_dout0(ap_bram_iarg_73_dout0),
        .ap_bram_73_we0(ap_bram_iarg_73_we0),
        .ap_bram_73_en0(ap_bram_iarg_73_en0),
        .ap_bram_73_addr1(ap_bram_iarg_73_addr1),
        .ap_bram_73_din1(ap_bram_iarg_73_din1),
        .ap_bram_73_dout1(ap_bram_iarg_73_dout1),
        .ap_bram_73_we1(ap_bram_iarg_73_we1),
        .ap_bram_73_en1(ap_bram_iarg_73_en1),
        .s_axis_bram_74_aclk(s_axis_bram_74_aclk),
        .s_axis_bram_74_aresetn(s_axis_bram_74_aresetn),
        .s_axis_bram_74_tlast(s_axis_bram_74_tlast),
        .s_axis_bram_74_tvalid(s_axis_bram_74_tvalid),
        .s_axis_bram_74_tkeep(s_axis_bram_74_tkeep),
        .s_axis_bram_74_tstrb(s_axis_bram_74_tstrb),
        .s_axis_bram_74_tdata(s_axis_bram_74_tdata),
        .s_axis_bram_74_tready(s_axis_bram_74_tready),
        .ap_bram_74_addr0(ap_bram_iarg_74_addr0),
        .ap_bram_74_din0(ap_bram_iarg_74_din0),
        .ap_bram_74_dout0(ap_bram_iarg_74_dout0),
        .ap_bram_74_we0(ap_bram_iarg_74_we0),
        .ap_bram_74_en0(ap_bram_iarg_74_en0),
        .ap_bram_74_addr1(ap_bram_iarg_74_addr1),
        .ap_bram_74_din1(ap_bram_iarg_74_din1),
        .ap_bram_74_dout1(ap_bram_iarg_74_dout1),
        .ap_bram_74_we1(ap_bram_iarg_74_we1),
        .ap_bram_74_en1(ap_bram_iarg_74_en1),
        .s_axis_bram_75_aclk(s_axis_bram_75_aclk),
        .s_axis_bram_75_aresetn(s_axis_bram_75_aresetn),
        .s_axis_bram_75_tlast(s_axis_bram_75_tlast),
        .s_axis_bram_75_tvalid(s_axis_bram_75_tvalid),
        .s_axis_bram_75_tkeep(s_axis_bram_75_tkeep),
        .s_axis_bram_75_tstrb(s_axis_bram_75_tstrb),
        .s_axis_bram_75_tdata(s_axis_bram_75_tdata),
        .s_axis_bram_75_tready(s_axis_bram_75_tready),
        .ap_bram_75_addr0(ap_bram_iarg_75_addr0),
        .ap_bram_75_din0(ap_bram_iarg_75_din0),
        .ap_bram_75_dout0(ap_bram_iarg_75_dout0),
        .ap_bram_75_we0(ap_bram_iarg_75_we0),
        .ap_bram_75_en0(ap_bram_iarg_75_en0),
        .ap_bram_75_addr1(ap_bram_iarg_75_addr1),
        .ap_bram_75_din1(ap_bram_iarg_75_din1),
        .ap_bram_75_dout1(ap_bram_iarg_75_dout1),
        .ap_bram_75_we1(ap_bram_iarg_75_we1),
        .ap_bram_75_en1(ap_bram_iarg_75_en1),
        .s_axis_bram_76_aclk(s_axis_bram_76_aclk),
        .s_axis_bram_76_aresetn(s_axis_bram_76_aresetn),
        .s_axis_bram_76_tlast(s_axis_bram_76_tlast),
        .s_axis_bram_76_tvalid(s_axis_bram_76_tvalid),
        .s_axis_bram_76_tkeep(s_axis_bram_76_tkeep),
        .s_axis_bram_76_tstrb(s_axis_bram_76_tstrb),
        .s_axis_bram_76_tdata(s_axis_bram_76_tdata),
        .s_axis_bram_76_tready(s_axis_bram_76_tready),
        .ap_bram_76_addr0(ap_bram_iarg_76_addr0),
        .ap_bram_76_din0(ap_bram_iarg_76_din0),
        .ap_bram_76_dout0(ap_bram_iarg_76_dout0),
        .ap_bram_76_we0(ap_bram_iarg_76_we0),
        .ap_bram_76_en0(ap_bram_iarg_76_en0),
        .ap_bram_76_addr1(ap_bram_iarg_76_addr1),
        .ap_bram_76_din1(ap_bram_iarg_76_din1),
        .ap_bram_76_dout1(ap_bram_iarg_76_dout1),
        .ap_bram_76_we1(ap_bram_iarg_76_we1),
        .ap_bram_76_en1(ap_bram_iarg_76_en1),
        .s_axis_bram_77_aclk(s_axis_bram_77_aclk),
        .s_axis_bram_77_aresetn(s_axis_bram_77_aresetn),
        .s_axis_bram_77_tlast(s_axis_bram_77_tlast),
        .s_axis_bram_77_tvalid(s_axis_bram_77_tvalid),
        .s_axis_bram_77_tkeep(s_axis_bram_77_tkeep),
        .s_axis_bram_77_tstrb(s_axis_bram_77_tstrb),
        .s_axis_bram_77_tdata(s_axis_bram_77_tdata),
        .s_axis_bram_77_tready(s_axis_bram_77_tready),
        .ap_bram_77_addr0(ap_bram_iarg_77_addr0),
        .ap_bram_77_din0(ap_bram_iarg_77_din0),
        .ap_bram_77_dout0(ap_bram_iarg_77_dout0),
        .ap_bram_77_we0(ap_bram_iarg_77_we0),
        .ap_bram_77_en0(ap_bram_iarg_77_en0),
        .ap_bram_77_addr1(ap_bram_iarg_77_addr1),
        .ap_bram_77_din1(ap_bram_iarg_77_din1),
        .ap_bram_77_dout1(ap_bram_iarg_77_dout1),
        .ap_bram_77_we1(ap_bram_iarg_77_we1),
        .ap_bram_77_en1(ap_bram_iarg_77_en1),
        .s_axis_bram_78_aclk(s_axis_bram_78_aclk),
        .s_axis_bram_78_aresetn(s_axis_bram_78_aresetn),
        .s_axis_bram_78_tlast(s_axis_bram_78_tlast),
        .s_axis_bram_78_tvalid(s_axis_bram_78_tvalid),
        .s_axis_bram_78_tkeep(s_axis_bram_78_tkeep),
        .s_axis_bram_78_tstrb(s_axis_bram_78_tstrb),
        .s_axis_bram_78_tdata(s_axis_bram_78_tdata),
        .s_axis_bram_78_tready(s_axis_bram_78_tready),
        .ap_bram_78_addr0(ap_bram_iarg_78_addr0),
        .ap_bram_78_din0(ap_bram_iarg_78_din0),
        .ap_bram_78_dout0(ap_bram_iarg_78_dout0),
        .ap_bram_78_we0(ap_bram_iarg_78_we0),
        .ap_bram_78_en0(ap_bram_iarg_78_en0),
        .ap_bram_78_addr1(ap_bram_iarg_78_addr1),
        .ap_bram_78_din1(ap_bram_iarg_78_din1),
        .ap_bram_78_dout1(ap_bram_iarg_78_dout1),
        .ap_bram_78_we1(ap_bram_iarg_78_we1),
        .ap_bram_78_en1(ap_bram_iarg_78_en1),
        .s_axis_bram_79_aclk(s_axis_bram_79_aclk),
        .s_axis_bram_79_aresetn(s_axis_bram_79_aresetn),
        .s_axis_bram_79_tlast(s_axis_bram_79_tlast),
        .s_axis_bram_79_tvalid(s_axis_bram_79_tvalid),
        .s_axis_bram_79_tkeep(s_axis_bram_79_tkeep),
        .s_axis_bram_79_tstrb(s_axis_bram_79_tstrb),
        .s_axis_bram_79_tdata(s_axis_bram_79_tdata),
        .s_axis_bram_79_tready(s_axis_bram_79_tready),
        .ap_bram_79_addr0(ap_bram_iarg_79_addr0),
        .ap_bram_79_din0(ap_bram_iarg_79_din0),
        .ap_bram_79_dout0(ap_bram_iarg_79_dout0),
        .ap_bram_79_we0(ap_bram_iarg_79_we0),
        .ap_bram_79_en0(ap_bram_iarg_79_en0),
        .ap_bram_79_addr1(ap_bram_iarg_79_addr1),
        .ap_bram_79_din1(ap_bram_iarg_79_din1),
        .ap_bram_79_dout1(ap_bram_iarg_79_dout1),
        .ap_bram_79_we1(ap_bram_iarg_79_we1),
        .ap_bram_79_en1(ap_bram_iarg_79_en1),
        .s_axis_bram_80_aclk(s_axis_bram_80_aclk),
        .s_axis_bram_80_aresetn(s_axis_bram_80_aresetn),
        .s_axis_bram_80_tlast(s_axis_bram_80_tlast),
        .s_axis_bram_80_tvalid(s_axis_bram_80_tvalid),
        .s_axis_bram_80_tkeep(s_axis_bram_80_tkeep),
        .s_axis_bram_80_tstrb(s_axis_bram_80_tstrb),
        .s_axis_bram_80_tdata(s_axis_bram_80_tdata),
        .s_axis_bram_80_tready(s_axis_bram_80_tready),
        .ap_bram_80_addr0(ap_bram_iarg_80_addr0),
        .ap_bram_80_din0(ap_bram_iarg_80_din0),
        .ap_bram_80_dout0(ap_bram_iarg_80_dout0),
        .ap_bram_80_we0(ap_bram_iarg_80_we0),
        .ap_bram_80_en0(ap_bram_iarg_80_en0),
        .ap_bram_80_addr1(ap_bram_iarg_80_addr1),
        .ap_bram_80_din1(ap_bram_iarg_80_din1),
        .ap_bram_80_dout1(ap_bram_iarg_80_dout1),
        .ap_bram_80_we1(ap_bram_iarg_80_we1),
        .ap_bram_80_en1(ap_bram_iarg_80_en1),
        .s_axis_bram_81_aclk(s_axis_bram_81_aclk),
        .s_axis_bram_81_aresetn(s_axis_bram_81_aresetn),
        .s_axis_bram_81_tlast(s_axis_bram_81_tlast),
        .s_axis_bram_81_tvalid(s_axis_bram_81_tvalid),
        .s_axis_bram_81_tkeep(s_axis_bram_81_tkeep),
        .s_axis_bram_81_tstrb(s_axis_bram_81_tstrb),
        .s_axis_bram_81_tdata(s_axis_bram_81_tdata),
        .s_axis_bram_81_tready(s_axis_bram_81_tready),
        .ap_bram_81_addr0(ap_bram_iarg_81_addr0),
        .ap_bram_81_din0(ap_bram_iarg_81_din0),
        .ap_bram_81_dout0(ap_bram_iarg_81_dout0),
        .ap_bram_81_we0(ap_bram_iarg_81_we0),
        .ap_bram_81_en0(ap_bram_iarg_81_en0),
        .ap_bram_81_addr1(ap_bram_iarg_81_addr1),
        .ap_bram_81_din1(ap_bram_iarg_81_din1),
        .ap_bram_81_dout1(ap_bram_iarg_81_dout1),
        .ap_bram_81_we1(ap_bram_iarg_81_we1),
        .ap_bram_81_en1(ap_bram_iarg_81_en1),
        .s_axis_bram_82_aclk(s_axis_bram_82_aclk),
        .s_axis_bram_82_aresetn(s_axis_bram_82_aresetn),
        .s_axis_bram_82_tlast(s_axis_bram_82_tlast),
        .s_axis_bram_82_tvalid(s_axis_bram_82_tvalid),
        .s_axis_bram_82_tkeep(s_axis_bram_82_tkeep),
        .s_axis_bram_82_tstrb(s_axis_bram_82_tstrb),
        .s_axis_bram_82_tdata(s_axis_bram_82_tdata),
        .s_axis_bram_82_tready(s_axis_bram_82_tready),
        .ap_bram_82_addr0(ap_bram_iarg_82_addr0),
        .ap_bram_82_din0(ap_bram_iarg_82_din0),
        .ap_bram_82_dout0(ap_bram_iarg_82_dout0),
        .ap_bram_82_we0(ap_bram_iarg_82_we0),
        .ap_bram_82_en0(ap_bram_iarg_82_en0),
        .ap_bram_82_addr1(ap_bram_iarg_82_addr1),
        .ap_bram_82_din1(ap_bram_iarg_82_din1),
        .ap_bram_82_dout1(ap_bram_iarg_82_dout1),
        .ap_bram_82_we1(ap_bram_iarg_82_we1),
        .ap_bram_82_en1(ap_bram_iarg_82_en1),
        .s_axis_bram_83_aclk(s_axis_bram_83_aclk),
        .s_axis_bram_83_aresetn(s_axis_bram_83_aresetn),
        .s_axis_bram_83_tlast(s_axis_bram_83_tlast),
        .s_axis_bram_83_tvalid(s_axis_bram_83_tvalid),
        .s_axis_bram_83_tkeep(s_axis_bram_83_tkeep),
        .s_axis_bram_83_tstrb(s_axis_bram_83_tstrb),
        .s_axis_bram_83_tdata(s_axis_bram_83_tdata),
        .s_axis_bram_83_tready(s_axis_bram_83_tready),
        .ap_bram_83_addr0(ap_bram_iarg_83_addr0),
        .ap_bram_83_din0(ap_bram_iarg_83_din0),
        .ap_bram_83_dout0(ap_bram_iarg_83_dout0),
        .ap_bram_83_we0(ap_bram_iarg_83_we0),
        .ap_bram_83_en0(ap_bram_iarg_83_en0),
        .ap_bram_83_addr1(ap_bram_iarg_83_addr1),
        .ap_bram_83_din1(ap_bram_iarg_83_din1),
        .ap_bram_83_dout1(ap_bram_iarg_83_dout1),
        .ap_bram_83_we1(ap_bram_iarg_83_we1),
        .ap_bram_83_en1(ap_bram_iarg_83_en1),
        .s_axis_bram_84_aclk(s_axis_bram_84_aclk),
        .s_axis_bram_84_aresetn(s_axis_bram_84_aresetn),
        .s_axis_bram_84_tlast(s_axis_bram_84_tlast),
        .s_axis_bram_84_tvalid(s_axis_bram_84_tvalid),
        .s_axis_bram_84_tkeep(s_axis_bram_84_tkeep),
        .s_axis_bram_84_tstrb(s_axis_bram_84_tstrb),
        .s_axis_bram_84_tdata(s_axis_bram_84_tdata),
        .s_axis_bram_84_tready(s_axis_bram_84_tready),
        .ap_bram_84_addr0(ap_bram_iarg_84_addr0),
        .ap_bram_84_din0(ap_bram_iarg_84_din0),
        .ap_bram_84_dout0(ap_bram_iarg_84_dout0),
        .ap_bram_84_we0(ap_bram_iarg_84_we0),
        .ap_bram_84_en0(ap_bram_iarg_84_en0),
        .ap_bram_84_addr1(ap_bram_iarg_84_addr1),
        .ap_bram_84_din1(ap_bram_iarg_84_din1),
        .ap_bram_84_dout1(ap_bram_iarg_84_dout1),
        .ap_bram_84_we1(ap_bram_iarg_84_we1),
        .ap_bram_84_en1(ap_bram_iarg_84_en1),
        .s_axis_bram_85_aclk(s_axis_bram_85_aclk),
        .s_axis_bram_85_aresetn(s_axis_bram_85_aresetn),
        .s_axis_bram_85_tlast(s_axis_bram_85_tlast),
        .s_axis_bram_85_tvalid(s_axis_bram_85_tvalid),
        .s_axis_bram_85_tkeep(s_axis_bram_85_tkeep),
        .s_axis_bram_85_tstrb(s_axis_bram_85_tstrb),
        .s_axis_bram_85_tdata(s_axis_bram_85_tdata),
        .s_axis_bram_85_tready(s_axis_bram_85_tready),
        .ap_bram_85_addr0(ap_bram_iarg_85_addr0),
        .ap_bram_85_din0(ap_bram_iarg_85_din0),
        .ap_bram_85_dout0(ap_bram_iarg_85_dout0),
        .ap_bram_85_we0(ap_bram_iarg_85_we0),
        .ap_bram_85_en0(ap_bram_iarg_85_en0),
        .ap_bram_85_addr1(ap_bram_iarg_85_addr1),
        .ap_bram_85_din1(ap_bram_iarg_85_din1),
        .ap_bram_85_dout1(ap_bram_iarg_85_dout1),
        .ap_bram_85_we1(ap_bram_iarg_85_we1),
        .ap_bram_85_en1(ap_bram_iarg_85_en1),
        .s_axis_bram_86_aclk(s_axis_bram_86_aclk),
        .s_axis_bram_86_aresetn(s_axis_bram_86_aresetn),
        .s_axis_bram_86_tlast(s_axis_bram_86_tlast),
        .s_axis_bram_86_tvalid(s_axis_bram_86_tvalid),
        .s_axis_bram_86_tkeep(s_axis_bram_86_tkeep),
        .s_axis_bram_86_tstrb(s_axis_bram_86_tstrb),
        .s_axis_bram_86_tdata(s_axis_bram_86_tdata),
        .s_axis_bram_86_tready(s_axis_bram_86_tready),
        .ap_bram_86_addr0(ap_bram_iarg_86_addr0),
        .ap_bram_86_din0(ap_bram_iarg_86_din0),
        .ap_bram_86_dout0(ap_bram_iarg_86_dout0),
        .ap_bram_86_we0(ap_bram_iarg_86_we0),
        .ap_bram_86_en0(ap_bram_iarg_86_en0),
        .ap_bram_86_addr1(ap_bram_iarg_86_addr1),
        .ap_bram_86_din1(ap_bram_iarg_86_din1),
        .ap_bram_86_dout1(ap_bram_iarg_86_dout1),
        .ap_bram_86_we1(ap_bram_iarg_86_we1),
        .ap_bram_86_en1(ap_bram_iarg_86_en1),
        .s_axis_bram_87_aclk(s_axis_bram_87_aclk),
        .s_axis_bram_87_aresetn(s_axis_bram_87_aresetn),
        .s_axis_bram_87_tlast(s_axis_bram_87_tlast),
        .s_axis_bram_87_tvalid(s_axis_bram_87_tvalid),
        .s_axis_bram_87_tkeep(s_axis_bram_87_tkeep),
        .s_axis_bram_87_tstrb(s_axis_bram_87_tstrb),
        .s_axis_bram_87_tdata(s_axis_bram_87_tdata),
        .s_axis_bram_87_tready(s_axis_bram_87_tready),
        .ap_bram_87_addr0(ap_bram_iarg_87_addr0),
        .ap_bram_87_din0(ap_bram_iarg_87_din0),
        .ap_bram_87_dout0(ap_bram_iarg_87_dout0),
        .ap_bram_87_we0(ap_bram_iarg_87_we0),
        .ap_bram_87_en0(ap_bram_iarg_87_en0),
        .ap_bram_87_addr1(ap_bram_iarg_87_addr1),
        .ap_bram_87_din1(ap_bram_iarg_87_din1),
        .ap_bram_87_dout1(ap_bram_iarg_87_dout1),
        .ap_bram_87_we1(ap_bram_iarg_87_we1),
        .ap_bram_87_en1(ap_bram_iarg_87_en1),
        .s_axis_bram_88_aclk(s_axis_bram_88_aclk),
        .s_axis_bram_88_aresetn(s_axis_bram_88_aresetn),
        .s_axis_bram_88_tlast(s_axis_bram_88_tlast),
        .s_axis_bram_88_tvalid(s_axis_bram_88_tvalid),
        .s_axis_bram_88_tkeep(s_axis_bram_88_tkeep),
        .s_axis_bram_88_tstrb(s_axis_bram_88_tstrb),
        .s_axis_bram_88_tdata(s_axis_bram_88_tdata),
        .s_axis_bram_88_tready(s_axis_bram_88_tready),
        .ap_bram_88_addr0(ap_bram_iarg_88_addr0),
        .ap_bram_88_din0(ap_bram_iarg_88_din0),
        .ap_bram_88_dout0(ap_bram_iarg_88_dout0),
        .ap_bram_88_we0(ap_bram_iarg_88_we0),
        .ap_bram_88_en0(ap_bram_iarg_88_en0),
        .ap_bram_88_addr1(ap_bram_iarg_88_addr1),
        .ap_bram_88_din1(ap_bram_iarg_88_din1),
        .ap_bram_88_dout1(ap_bram_iarg_88_dout1),
        .ap_bram_88_we1(ap_bram_iarg_88_we1),
        .ap_bram_88_en1(ap_bram_iarg_88_en1),
        .s_axis_bram_89_aclk(s_axis_bram_89_aclk),
        .s_axis_bram_89_aresetn(s_axis_bram_89_aresetn),
        .s_axis_bram_89_tlast(s_axis_bram_89_tlast),
        .s_axis_bram_89_tvalid(s_axis_bram_89_tvalid),
        .s_axis_bram_89_tkeep(s_axis_bram_89_tkeep),
        .s_axis_bram_89_tstrb(s_axis_bram_89_tstrb),
        .s_axis_bram_89_tdata(s_axis_bram_89_tdata),
        .s_axis_bram_89_tready(s_axis_bram_89_tready),
        .ap_bram_89_addr0(ap_bram_iarg_89_addr0),
        .ap_bram_89_din0(ap_bram_iarg_89_din0),
        .ap_bram_89_dout0(ap_bram_iarg_89_dout0),
        .ap_bram_89_we0(ap_bram_iarg_89_we0),
        .ap_bram_89_en0(ap_bram_iarg_89_en0),
        .ap_bram_89_addr1(ap_bram_iarg_89_addr1),
        .ap_bram_89_din1(ap_bram_iarg_89_din1),
        .ap_bram_89_dout1(ap_bram_iarg_89_dout1),
        .ap_bram_89_we1(ap_bram_iarg_89_we1),
        .ap_bram_89_en1(ap_bram_iarg_89_en1),
        .s_axis_bram_90_aclk(s_axis_bram_90_aclk),
        .s_axis_bram_90_aresetn(s_axis_bram_90_aresetn),
        .s_axis_bram_90_tlast(s_axis_bram_90_tlast),
        .s_axis_bram_90_tvalid(s_axis_bram_90_tvalid),
        .s_axis_bram_90_tkeep(s_axis_bram_90_tkeep),
        .s_axis_bram_90_tstrb(s_axis_bram_90_tstrb),
        .s_axis_bram_90_tdata(s_axis_bram_90_tdata),
        .s_axis_bram_90_tready(s_axis_bram_90_tready),
        .ap_bram_90_addr0(ap_bram_iarg_90_addr0),
        .ap_bram_90_din0(ap_bram_iarg_90_din0),
        .ap_bram_90_dout0(ap_bram_iarg_90_dout0),
        .ap_bram_90_we0(ap_bram_iarg_90_we0),
        .ap_bram_90_en0(ap_bram_iarg_90_en0),
        .ap_bram_90_addr1(ap_bram_iarg_90_addr1),
        .ap_bram_90_din1(ap_bram_iarg_90_din1),
        .ap_bram_90_dout1(ap_bram_iarg_90_dout1),
        .ap_bram_90_we1(ap_bram_iarg_90_we1),
        .ap_bram_90_en1(ap_bram_iarg_90_en1),
        .s_axis_bram_91_aclk(s_axis_bram_91_aclk),
        .s_axis_bram_91_aresetn(s_axis_bram_91_aresetn),
        .s_axis_bram_91_tlast(s_axis_bram_91_tlast),
        .s_axis_bram_91_tvalid(s_axis_bram_91_tvalid),
        .s_axis_bram_91_tkeep(s_axis_bram_91_tkeep),
        .s_axis_bram_91_tstrb(s_axis_bram_91_tstrb),
        .s_axis_bram_91_tdata(s_axis_bram_91_tdata),
        .s_axis_bram_91_tready(s_axis_bram_91_tready),
        .ap_bram_91_addr0(ap_bram_iarg_91_addr0),
        .ap_bram_91_din0(ap_bram_iarg_91_din0),
        .ap_bram_91_dout0(ap_bram_iarg_91_dout0),
        .ap_bram_91_we0(ap_bram_iarg_91_we0),
        .ap_bram_91_en0(ap_bram_iarg_91_en0),
        .ap_bram_91_addr1(ap_bram_iarg_91_addr1),
        .ap_bram_91_din1(ap_bram_iarg_91_din1),
        .ap_bram_91_dout1(ap_bram_iarg_91_dout1),
        .ap_bram_91_we1(ap_bram_iarg_91_we1),
        .ap_bram_91_en1(ap_bram_iarg_91_en1),
        .s_axis_bram_92_aclk(s_axis_bram_92_aclk),
        .s_axis_bram_92_aresetn(s_axis_bram_92_aresetn),
        .s_axis_bram_92_tlast(s_axis_bram_92_tlast),
        .s_axis_bram_92_tvalid(s_axis_bram_92_tvalid),
        .s_axis_bram_92_tkeep(s_axis_bram_92_tkeep),
        .s_axis_bram_92_tstrb(s_axis_bram_92_tstrb),
        .s_axis_bram_92_tdata(s_axis_bram_92_tdata),
        .s_axis_bram_92_tready(s_axis_bram_92_tready),
        .ap_bram_92_addr0(ap_bram_iarg_92_addr0),
        .ap_bram_92_din0(ap_bram_iarg_92_din0),
        .ap_bram_92_dout0(ap_bram_iarg_92_dout0),
        .ap_bram_92_we0(ap_bram_iarg_92_we0),
        .ap_bram_92_en0(ap_bram_iarg_92_en0),
        .ap_bram_92_addr1(ap_bram_iarg_92_addr1),
        .ap_bram_92_din1(ap_bram_iarg_92_din1),
        .ap_bram_92_dout1(ap_bram_iarg_92_dout1),
        .ap_bram_92_we1(ap_bram_iarg_92_we1),
        .ap_bram_92_en1(ap_bram_iarg_92_en1),
        .s_axis_bram_93_aclk(s_axis_bram_93_aclk),
        .s_axis_bram_93_aresetn(s_axis_bram_93_aresetn),
        .s_axis_bram_93_tlast(s_axis_bram_93_tlast),
        .s_axis_bram_93_tvalid(s_axis_bram_93_tvalid),
        .s_axis_bram_93_tkeep(s_axis_bram_93_tkeep),
        .s_axis_bram_93_tstrb(s_axis_bram_93_tstrb),
        .s_axis_bram_93_tdata(s_axis_bram_93_tdata),
        .s_axis_bram_93_tready(s_axis_bram_93_tready),
        .ap_bram_93_addr0(ap_bram_iarg_93_addr0),
        .ap_bram_93_din0(ap_bram_iarg_93_din0),
        .ap_bram_93_dout0(ap_bram_iarg_93_dout0),
        .ap_bram_93_we0(ap_bram_iarg_93_we0),
        .ap_bram_93_en0(ap_bram_iarg_93_en0),
        .ap_bram_93_addr1(ap_bram_iarg_93_addr1),
        .ap_bram_93_din1(ap_bram_iarg_93_din1),
        .ap_bram_93_dout1(ap_bram_iarg_93_dout1),
        .ap_bram_93_we1(ap_bram_iarg_93_we1),
        .ap_bram_93_en1(ap_bram_iarg_93_en1),
        .s_axis_bram_94_aclk(s_axis_bram_94_aclk),
        .s_axis_bram_94_aresetn(s_axis_bram_94_aresetn),
        .s_axis_bram_94_tlast(s_axis_bram_94_tlast),
        .s_axis_bram_94_tvalid(s_axis_bram_94_tvalid),
        .s_axis_bram_94_tkeep(s_axis_bram_94_tkeep),
        .s_axis_bram_94_tstrb(s_axis_bram_94_tstrb),
        .s_axis_bram_94_tdata(s_axis_bram_94_tdata),
        .s_axis_bram_94_tready(s_axis_bram_94_tready),
        .ap_bram_94_addr0(ap_bram_iarg_94_addr0),
        .ap_bram_94_din0(ap_bram_iarg_94_din0),
        .ap_bram_94_dout0(ap_bram_iarg_94_dout0),
        .ap_bram_94_we0(ap_bram_iarg_94_we0),
        .ap_bram_94_en0(ap_bram_iarg_94_en0),
        .ap_bram_94_addr1(ap_bram_iarg_94_addr1),
        .ap_bram_94_din1(ap_bram_iarg_94_din1),
        .ap_bram_94_dout1(ap_bram_iarg_94_dout1),
        .ap_bram_94_we1(ap_bram_iarg_94_we1),
        .ap_bram_94_en1(ap_bram_iarg_94_en1),
        .s_axis_bram_95_aclk(s_axis_bram_95_aclk),
        .s_axis_bram_95_aresetn(s_axis_bram_95_aresetn),
        .s_axis_bram_95_tlast(s_axis_bram_95_tlast),
        .s_axis_bram_95_tvalid(s_axis_bram_95_tvalid),
        .s_axis_bram_95_tkeep(s_axis_bram_95_tkeep),
        .s_axis_bram_95_tstrb(s_axis_bram_95_tstrb),
        .s_axis_bram_95_tdata(s_axis_bram_95_tdata),
        .s_axis_bram_95_tready(s_axis_bram_95_tready),
        .ap_bram_95_addr0(ap_bram_iarg_95_addr0),
        .ap_bram_95_din0(ap_bram_iarg_95_din0),
        .ap_bram_95_dout0(ap_bram_iarg_95_dout0),
        .ap_bram_95_we0(ap_bram_iarg_95_we0),
        .ap_bram_95_en0(ap_bram_iarg_95_en0),
        .ap_bram_95_addr1(ap_bram_iarg_95_addr1),
        .ap_bram_95_din1(ap_bram_iarg_95_din1),
        .ap_bram_95_dout1(ap_bram_iarg_95_dout1),
        .ap_bram_95_we1(ap_bram_iarg_95_we1),
        .ap_bram_95_en1(ap_bram_iarg_95_en1),
        .s_axis_bram_96_aclk(s_axis_bram_96_aclk),
        .s_axis_bram_96_aresetn(s_axis_bram_96_aresetn),
        .s_axis_bram_96_tlast(s_axis_bram_96_tlast),
        .s_axis_bram_96_tvalid(s_axis_bram_96_tvalid),
        .s_axis_bram_96_tkeep(s_axis_bram_96_tkeep),
        .s_axis_bram_96_tstrb(s_axis_bram_96_tstrb),
        .s_axis_bram_96_tdata(s_axis_bram_96_tdata),
        .s_axis_bram_96_tready(s_axis_bram_96_tready),
        .ap_bram_96_addr0(ap_bram_iarg_96_addr0),
        .ap_bram_96_din0(ap_bram_iarg_96_din0),
        .ap_bram_96_dout0(ap_bram_iarg_96_dout0),
        .ap_bram_96_we0(ap_bram_iarg_96_we0),
        .ap_bram_96_en0(ap_bram_iarg_96_en0),
        .ap_bram_96_addr1(ap_bram_iarg_96_addr1),
        .ap_bram_96_din1(ap_bram_iarg_96_din1),
        .ap_bram_96_dout1(ap_bram_iarg_96_dout1),
        .ap_bram_96_we1(ap_bram_iarg_96_we1),
        .ap_bram_96_en1(ap_bram_iarg_96_en1),
        .s_axis_bram_97_aclk(s_axis_bram_97_aclk),
        .s_axis_bram_97_aresetn(s_axis_bram_97_aresetn),
        .s_axis_bram_97_tlast(s_axis_bram_97_tlast),
        .s_axis_bram_97_tvalid(s_axis_bram_97_tvalid),
        .s_axis_bram_97_tkeep(s_axis_bram_97_tkeep),
        .s_axis_bram_97_tstrb(s_axis_bram_97_tstrb),
        .s_axis_bram_97_tdata(s_axis_bram_97_tdata),
        .s_axis_bram_97_tready(s_axis_bram_97_tready),
        .ap_bram_97_addr0(ap_bram_iarg_97_addr0),
        .ap_bram_97_din0(ap_bram_iarg_97_din0),
        .ap_bram_97_dout0(ap_bram_iarg_97_dout0),
        .ap_bram_97_we0(ap_bram_iarg_97_we0),
        .ap_bram_97_en0(ap_bram_iarg_97_en0),
        .ap_bram_97_addr1(ap_bram_iarg_97_addr1),
        .ap_bram_97_din1(ap_bram_iarg_97_din1),
        .ap_bram_97_dout1(ap_bram_iarg_97_dout1),
        .ap_bram_97_we1(ap_bram_iarg_97_we1),
        .ap_bram_97_en1(ap_bram_iarg_97_en1),
        .s_axis_bram_98_aclk(s_axis_bram_98_aclk),
        .s_axis_bram_98_aresetn(s_axis_bram_98_aresetn),
        .s_axis_bram_98_tlast(s_axis_bram_98_tlast),
        .s_axis_bram_98_tvalid(s_axis_bram_98_tvalid),
        .s_axis_bram_98_tkeep(s_axis_bram_98_tkeep),
        .s_axis_bram_98_tstrb(s_axis_bram_98_tstrb),
        .s_axis_bram_98_tdata(s_axis_bram_98_tdata),
        .s_axis_bram_98_tready(s_axis_bram_98_tready),
        .ap_bram_98_addr0(ap_bram_iarg_98_addr0),
        .ap_bram_98_din0(ap_bram_iarg_98_din0),
        .ap_bram_98_dout0(ap_bram_iarg_98_dout0),
        .ap_bram_98_we0(ap_bram_iarg_98_we0),
        .ap_bram_98_en0(ap_bram_iarg_98_en0),
        .ap_bram_98_addr1(ap_bram_iarg_98_addr1),
        .ap_bram_98_din1(ap_bram_iarg_98_din1),
        .ap_bram_98_dout1(ap_bram_iarg_98_dout1),
        .ap_bram_98_we1(ap_bram_iarg_98_we1),
        .ap_bram_98_en1(ap_bram_iarg_98_en1),
        .s_axis_bram_99_aclk(s_axis_bram_99_aclk),
        .s_axis_bram_99_aresetn(s_axis_bram_99_aresetn),
        .s_axis_bram_99_tlast(s_axis_bram_99_tlast),
        .s_axis_bram_99_tvalid(s_axis_bram_99_tvalid),
        .s_axis_bram_99_tkeep(s_axis_bram_99_tkeep),
        .s_axis_bram_99_tstrb(s_axis_bram_99_tstrb),
        .s_axis_bram_99_tdata(s_axis_bram_99_tdata),
        .s_axis_bram_99_tready(s_axis_bram_99_tready),
        .ap_bram_99_addr0(ap_bram_iarg_99_addr0),
        .ap_bram_99_din0(ap_bram_iarg_99_din0),
        .ap_bram_99_dout0(ap_bram_iarg_99_dout0),
        .ap_bram_99_we0(ap_bram_iarg_99_we0),
        .ap_bram_99_en0(ap_bram_iarg_99_en0),
        .ap_bram_99_addr1(ap_bram_iarg_99_addr1),
        .ap_bram_99_din1(ap_bram_iarg_99_din1),
        .ap_bram_99_dout1(ap_bram_iarg_99_dout1),
        .ap_bram_99_we1(ap_bram_iarg_99_we1),
        .ap_bram_99_en1(ap_bram_iarg_99_en1),
        .s_axis_bram_100_aclk(s_axis_bram_100_aclk),
        .s_axis_bram_100_aresetn(s_axis_bram_100_aresetn),
        .s_axis_bram_100_tlast(s_axis_bram_100_tlast),
        .s_axis_bram_100_tvalid(s_axis_bram_100_tvalid),
        .s_axis_bram_100_tkeep(s_axis_bram_100_tkeep),
        .s_axis_bram_100_tstrb(s_axis_bram_100_tstrb),
        .s_axis_bram_100_tdata(s_axis_bram_100_tdata),
        .s_axis_bram_100_tready(s_axis_bram_100_tready),
        .ap_bram_100_addr0(ap_bram_iarg_100_addr0),
        .ap_bram_100_din0(ap_bram_iarg_100_din0),
        .ap_bram_100_dout0(ap_bram_iarg_100_dout0),
        .ap_bram_100_we0(ap_bram_iarg_100_we0),
        .ap_bram_100_en0(ap_bram_iarg_100_en0),
        .ap_bram_100_addr1(ap_bram_iarg_100_addr1),
        .ap_bram_100_din1(ap_bram_iarg_100_din1),
        .ap_bram_100_dout1(ap_bram_iarg_100_dout1),
        .ap_bram_100_we1(ap_bram_iarg_100_we1),
        .ap_bram_100_en1(ap_bram_iarg_100_en1),
        .s_axis_bram_101_aclk(s_axis_bram_101_aclk),
        .s_axis_bram_101_aresetn(s_axis_bram_101_aresetn),
        .s_axis_bram_101_tlast(s_axis_bram_101_tlast),
        .s_axis_bram_101_tvalid(s_axis_bram_101_tvalid),
        .s_axis_bram_101_tkeep(s_axis_bram_101_tkeep),
        .s_axis_bram_101_tstrb(s_axis_bram_101_tstrb),
        .s_axis_bram_101_tdata(s_axis_bram_101_tdata),
        .s_axis_bram_101_tready(s_axis_bram_101_tready),
        .ap_bram_101_addr0(ap_bram_iarg_101_addr0),
        .ap_bram_101_din0(ap_bram_iarg_101_din0),
        .ap_bram_101_dout0(ap_bram_iarg_101_dout0),
        .ap_bram_101_we0(ap_bram_iarg_101_we0),
        .ap_bram_101_en0(ap_bram_iarg_101_en0),
        .ap_bram_101_addr1(ap_bram_iarg_101_addr1),
        .ap_bram_101_din1(ap_bram_iarg_101_din1),
        .ap_bram_101_dout1(ap_bram_iarg_101_dout1),
        .ap_bram_101_we1(ap_bram_iarg_101_we1),
        .ap_bram_101_en1(ap_bram_iarg_101_en1),
        .s_axis_bram_102_aclk(s_axis_bram_102_aclk),
        .s_axis_bram_102_aresetn(s_axis_bram_102_aresetn),
        .s_axis_bram_102_tlast(s_axis_bram_102_tlast),
        .s_axis_bram_102_tvalid(s_axis_bram_102_tvalid),
        .s_axis_bram_102_tkeep(s_axis_bram_102_tkeep),
        .s_axis_bram_102_tstrb(s_axis_bram_102_tstrb),
        .s_axis_bram_102_tdata(s_axis_bram_102_tdata),
        .s_axis_bram_102_tready(s_axis_bram_102_tready),
        .ap_bram_102_addr0(ap_bram_iarg_102_addr0),
        .ap_bram_102_din0(ap_bram_iarg_102_din0),
        .ap_bram_102_dout0(ap_bram_iarg_102_dout0),
        .ap_bram_102_we0(ap_bram_iarg_102_we0),
        .ap_bram_102_en0(ap_bram_iarg_102_en0),
        .ap_bram_102_addr1(ap_bram_iarg_102_addr1),
        .ap_bram_102_din1(ap_bram_iarg_102_din1),
        .ap_bram_102_dout1(ap_bram_iarg_102_dout1),
        .ap_bram_102_we1(ap_bram_iarg_102_we1),
        .ap_bram_102_en1(ap_bram_iarg_102_en1),
        .s_axis_bram_103_aclk(s_axis_bram_103_aclk),
        .s_axis_bram_103_aresetn(s_axis_bram_103_aresetn),
        .s_axis_bram_103_tlast(s_axis_bram_103_tlast),
        .s_axis_bram_103_tvalid(s_axis_bram_103_tvalid),
        .s_axis_bram_103_tkeep(s_axis_bram_103_tkeep),
        .s_axis_bram_103_tstrb(s_axis_bram_103_tstrb),
        .s_axis_bram_103_tdata(s_axis_bram_103_tdata),
        .s_axis_bram_103_tready(s_axis_bram_103_tready),
        .ap_bram_103_addr0(ap_bram_iarg_103_addr0),
        .ap_bram_103_din0(ap_bram_iarg_103_din0),
        .ap_bram_103_dout0(ap_bram_iarg_103_dout0),
        .ap_bram_103_we0(ap_bram_iarg_103_we0),
        .ap_bram_103_en0(ap_bram_iarg_103_en0),
        .ap_bram_103_addr1(ap_bram_iarg_103_addr1),
        .ap_bram_103_din1(ap_bram_iarg_103_din1),
        .ap_bram_103_dout1(ap_bram_iarg_103_dout1),
        .ap_bram_103_we1(ap_bram_iarg_103_we1),
        .ap_bram_103_en1(ap_bram_iarg_103_en1),
        .s_axis_bram_104_aclk(s_axis_bram_104_aclk),
        .s_axis_bram_104_aresetn(s_axis_bram_104_aresetn),
        .s_axis_bram_104_tlast(s_axis_bram_104_tlast),
        .s_axis_bram_104_tvalid(s_axis_bram_104_tvalid),
        .s_axis_bram_104_tkeep(s_axis_bram_104_tkeep),
        .s_axis_bram_104_tstrb(s_axis_bram_104_tstrb),
        .s_axis_bram_104_tdata(s_axis_bram_104_tdata),
        .s_axis_bram_104_tready(s_axis_bram_104_tready),
        .ap_bram_104_addr0(ap_bram_iarg_104_addr0),
        .ap_bram_104_din0(ap_bram_iarg_104_din0),
        .ap_bram_104_dout0(ap_bram_iarg_104_dout0),
        .ap_bram_104_we0(ap_bram_iarg_104_we0),
        .ap_bram_104_en0(ap_bram_iarg_104_en0),
        .ap_bram_104_addr1(ap_bram_iarg_104_addr1),
        .ap_bram_104_din1(ap_bram_iarg_104_din1),
        .ap_bram_104_dout1(ap_bram_iarg_104_dout1),
        .ap_bram_104_we1(ap_bram_iarg_104_we1),
        .ap_bram_104_en1(ap_bram_iarg_104_en1),
        .s_axis_bram_105_aclk(s_axis_bram_105_aclk),
        .s_axis_bram_105_aresetn(s_axis_bram_105_aresetn),
        .s_axis_bram_105_tlast(s_axis_bram_105_tlast),
        .s_axis_bram_105_tvalid(s_axis_bram_105_tvalid),
        .s_axis_bram_105_tkeep(s_axis_bram_105_tkeep),
        .s_axis_bram_105_tstrb(s_axis_bram_105_tstrb),
        .s_axis_bram_105_tdata(s_axis_bram_105_tdata),
        .s_axis_bram_105_tready(s_axis_bram_105_tready),
        .ap_bram_105_addr0(ap_bram_iarg_105_addr0),
        .ap_bram_105_din0(ap_bram_iarg_105_din0),
        .ap_bram_105_dout0(ap_bram_iarg_105_dout0),
        .ap_bram_105_we0(ap_bram_iarg_105_we0),
        .ap_bram_105_en0(ap_bram_iarg_105_en0),
        .ap_bram_105_addr1(ap_bram_iarg_105_addr1),
        .ap_bram_105_din1(ap_bram_iarg_105_din1),
        .ap_bram_105_dout1(ap_bram_iarg_105_dout1),
        .ap_bram_105_we1(ap_bram_iarg_105_we1),
        .ap_bram_105_en1(ap_bram_iarg_105_en1),
        .s_axis_bram_106_aclk(s_axis_bram_106_aclk),
        .s_axis_bram_106_aresetn(s_axis_bram_106_aresetn),
        .s_axis_bram_106_tlast(s_axis_bram_106_tlast),
        .s_axis_bram_106_tvalid(s_axis_bram_106_tvalid),
        .s_axis_bram_106_tkeep(s_axis_bram_106_tkeep),
        .s_axis_bram_106_tstrb(s_axis_bram_106_tstrb),
        .s_axis_bram_106_tdata(s_axis_bram_106_tdata),
        .s_axis_bram_106_tready(s_axis_bram_106_tready),
        .ap_bram_106_addr0(ap_bram_iarg_106_addr0),
        .ap_bram_106_din0(ap_bram_iarg_106_din0),
        .ap_bram_106_dout0(ap_bram_iarg_106_dout0),
        .ap_bram_106_we0(ap_bram_iarg_106_we0),
        .ap_bram_106_en0(ap_bram_iarg_106_en0),
        .ap_bram_106_addr1(ap_bram_iarg_106_addr1),
        .ap_bram_106_din1(ap_bram_iarg_106_din1),
        .ap_bram_106_dout1(ap_bram_iarg_106_dout1),
        .ap_bram_106_we1(ap_bram_iarg_106_we1),
        .ap_bram_106_en1(ap_bram_iarg_106_en1),
        .s_axis_bram_107_aclk(s_axis_bram_107_aclk),
        .s_axis_bram_107_aresetn(s_axis_bram_107_aresetn),
        .s_axis_bram_107_tlast(s_axis_bram_107_tlast),
        .s_axis_bram_107_tvalid(s_axis_bram_107_tvalid),
        .s_axis_bram_107_tkeep(s_axis_bram_107_tkeep),
        .s_axis_bram_107_tstrb(s_axis_bram_107_tstrb),
        .s_axis_bram_107_tdata(s_axis_bram_107_tdata),
        .s_axis_bram_107_tready(s_axis_bram_107_tready),
        .ap_bram_107_addr0(ap_bram_iarg_107_addr0),
        .ap_bram_107_din0(ap_bram_iarg_107_din0),
        .ap_bram_107_dout0(ap_bram_iarg_107_dout0),
        .ap_bram_107_we0(ap_bram_iarg_107_we0),
        .ap_bram_107_en0(ap_bram_iarg_107_en0),
        .ap_bram_107_addr1(ap_bram_iarg_107_addr1),
        .ap_bram_107_din1(ap_bram_iarg_107_din1),
        .ap_bram_107_dout1(ap_bram_iarg_107_dout1),
        .ap_bram_107_we1(ap_bram_iarg_107_we1),
        .ap_bram_107_en1(ap_bram_iarg_107_en1),
        .s_axis_bram_108_aclk(s_axis_bram_108_aclk),
        .s_axis_bram_108_aresetn(s_axis_bram_108_aresetn),
        .s_axis_bram_108_tlast(s_axis_bram_108_tlast),
        .s_axis_bram_108_tvalid(s_axis_bram_108_tvalid),
        .s_axis_bram_108_tkeep(s_axis_bram_108_tkeep),
        .s_axis_bram_108_tstrb(s_axis_bram_108_tstrb),
        .s_axis_bram_108_tdata(s_axis_bram_108_tdata),
        .s_axis_bram_108_tready(s_axis_bram_108_tready),
        .ap_bram_108_addr0(ap_bram_iarg_108_addr0),
        .ap_bram_108_din0(ap_bram_iarg_108_din0),
        .ap_bram_108_dout0(ap_bram_iarg_108_dout0),
        .ap_bram_108_we0(ap_bram_iarg_108_we0),
        .ap_bram_108_en0(ap_bram_iarg_108_en0),
        .ap_bram_108_addr1(ap_bram_iarg_108_addr1),
        .ap_bram_108_din1(ap_bram_iarg_108_din1),
        .ap_bram_108_dout1(ap_bram_iarg_108_dout1),
        .ap_bram_108_we1(ap_bram_iarg_108_we1),
        .ap_bram_108_en1(ap_bram_iarg_108_en1),
        .s_axis_bram_109_aclk(s_axis_bram_109_aclk),
        .s_axis_bram_109_aresetn(s_axis_bram_109_aresetn),
        .s_axis_bram_109_tlast(s_axis_bram_109_tlast),
        .s_axis_bram_109_tvalid(s_axis_bram_109_tvalid),
        .s_axis_bram_109_tkeep(s_axis_bram_109_tkeep),
        .s_axis_bram_109_tstrb(s_axis_bram_109_tstrb),
        .s_axis_bram_109_tdata(s_axis_bram_109_tdata),
        .s_axis_bram_109_tready(s_axis_bram_109_tready),
        .ap_bram_109_addr0(ap_bram_iarg_109_addr0),
        .ap_bram_109_din0(ap_bram_iarg_109_din0),
        .ap_bram_109_dout0(ap_bram_iarg_109_dout0),
        .ap_bram_109_we0(ap_bram_iarg_109_we0),
        .ap_bram_109_en0(ap_bram_iarg_109_en0),
        .ap_bram_109_addr1(ap_bram_iarg_109_addr1),
        .ap_bram_109_din1(ap_bram_iarg_109_din1),
        .ap_bram_109_dout1(ap_bram_iarg_109_dout1),
        .ap_bram_109_we1(ap_bram_iarg_109_we1),
        .ap_bram_109_en1(ap_bram_iarg_109_en1),
        .s_axis_bram_110_aclk(s_axis_bram_110_aclk),
        .s_axis_bram_110_aresetn(s_axis_bram_110_aresetn),
        .s_axis_bram_110_tlast(s_axis_bram_110_tlast),
        .s_axis_bram_110_tvalid(s_axis_bram_110_tvalid),
        .s_axis_bram_110_tkeep(s_axis_bram_110_tkeep),
        .s_axis_bram_110_tstrb(s_axis_bram_110_tstrb),
        .s_axis_bram_110_tdata(s_axis_bram_110_tdata),
        .s_axis_bram_110_tready(s_axis_bram_110_tready),
        .ap_bram_110_addr0(ap_bram_iarg_110_addr0),
        .ap_bram_110_din0(ap_bram_iarg_110_din0),
        .ap_bram_110_dout0(ap_bram_iarg_110_dout0),
        .ap_bram_110_we0(ap_bram_iarg_110_we0),
        .ap_bram_110_en0(ap_bram_iarg_110_en0),
        .ap_bram_110_addr1(ap_bram_iarg_110_addr1),
        .ap_bram_110_din1(ap_bram_iarg_110_din1),
        .ap_bram_110_dout1(ap_bram_iarg_110_dout1),
        .ap_bram_110_we1(ap_bram_iarg_110_we1),
        .ap_bram_110_en1(ap_bram_iarg_110_en1),
        .s_axis_bram_111_aclk(s_axis_bram_111_aclk),
        .s_axis_bram_111_aresetn(s_axis_bram_111_aresetn),
        .s_axis_bram_111_tlast(s_axis_bram_111_tlast),
        .s_axis_bram_111_tvalid(s_axis_bram_111_tvalid),
        .s_axis_bram_111_tkeep(s_axis_bram_111_tkeep),
        .s_axis_bram_111_tstrb(s_axis_bram_111_tstrb),
        .s_axis_bram_111_tdata(s_axis_bram_111_tdata),
        .s_axis_bram_111_tready(s_axis_bram_111_tready),
        .ap_bram_111_addr0(ap_bram_iarg_111_addr0),
        .ap_bram_111_din0(ap_bram_iarg_111_din0),
        .ap_bram_111_dout0(ap_bram_iarg_111_dout0),
        .ap_bram_111_we0(ap_bram_iarg_111_we0),
        .ap_bram_111_en0(ap_bram_iarg_111_en0),
        .ap_bram_111_addr1(ap_bram_iarg_111_addr1),
        .ap_bram_111_din1(ap_bram_iarg_111_din1),
        .ap_bram_111_dout1(ap_bram_iarg_111_dout1),
        .ap_bram_111_we1(ap_bram_iarg_111_we1),
        .ap_bram_111_en1(ap_bram_iarg_111_en1),
        .s_axis_bram_112_aclk(s_axis_bram_112_aclk),
        .s_axis_bram_112_aresetn(s_axis_bram_112_aresetn),
        .s_axis_bram_112_tlast(s_axis_bram_112_tlast),
        .s_axis_bram_112_tvalid(s_axis_bram_112_tvalid),
        .s_axis_bram_112_tkeep(s_axis_bram_112_tkeep),
        .s_axis_bram_112_tstrb(s_axis_bram_112_tstrb),
        .s_axis_bram_112_tdata(s_axis_bram_112_tdata),
        .s_axis_bram_112_tready(s_axis_bram_112_tready),
        .ap_bram_112_addr0(ap_bram_iarg_112_addr0),
        .ap_bram_112_din0(ap_bram_iarg_112_din0),
        .ap_bram_112_dout0(ap_bram_iarg_112_dout0),
        .ap_bram_112_we0(ap_bram_iarg_112_we0),
        .ap_bram_112_en0(ap_bram_iarg_112_en0),
        .ap_bram_112_addr1(ap_bram_iarg_112_addr1),
        .ap_bram_112_din1(ap_bram_iarg_112_din1),
        .ap_bram_112_dout1(ap_bram_iarg_112_dout1),
        .ap_bram_112_we1(ap_bram_iarg_112_we1),
        .ap_bram_112_en1(ap_bram_iarg_112_en1),
        .s_axis_bram_113_aclk(s_axis_bram_113_aclk),
        .s_axis_bram_113_aresetn(s_axis_bram_113_aresetn),
        .s_axis_bram_113_tlast(s_axis_bram_113_tlast),
        .s_axis_bram_113_tvalid(s_axis_bram_113_tvalid),
        .s_axis_bram_113_tkeep(s_axis_bram_113_tkeep),
        .s_axis_bram_113_tstrb(s_axis_bram_113_tstrb),
        .s_axis_bram_113_tdata(s_axis_bram_113_tdata),
        .s_axis_bram_113_tready(s_axis_bram_113_tready),
        .ap_bram_113_addr0(ap_bram_iarg_113_addr0),
        .ap_bram_113_din0(ap_bram_iarg_113_din0),
        .ap_bram_113_dout0(ap_bram_iarg_113_dout0),
        .ap_bram_113_we0(ap_bram_iarg_113_we0),
        .ap_bram_113_en0(ap_bram_iarg_113_en0),
        .ap_bram_113_addr1(ap_bram_iarg_113_addr1),
        .ap_bram_113_din1(ap_bram_iarg_113_din1),
        .ap_bram_113_dout1(ap_bram_iarg_113_dout1),
        .ap_bram_113_we1(ap_bram_iarg_113_we1),
        .ap_bram_113_en1(ap_bram_iarg_113_en1),
        .s_axis_bram_114_aclk(s_axis_bram_114_aclk),
        .s_axis_bram_114_aresetn(s_axis_bram_114_aresetn),
        .s_axis_bram_114_tlast(s_axis_bram_114_tlast),
        .s_axis_bram_114_tvalid(s_axis_bram_114_tvalid),
        .s_axis_bram_114_tkeep(s_axis_bram_114_tkeep),
        .s_axis_bram_114_tstrb(s_axis_bram_114_tstrb),
        .s_axis_bram_114_tdata(s_axis_bram_114_tdata),
        .s_axis_bram_114_tready(s_axis_bram_114_tready),
        .ap_bram_114_addr0(ap_bram_iarg_114_addr0),
        .ap_bram_114_din0(ap_bram_iarg_114_din0),
        .ap_bram_114_dout0(ap_bram_iarg_114_dout0),
        .ap_bram_114_we0(ap_bram_iarg_114_we0),
        .ap_bram_114_en0(ap_bram_iarg_114_en0),
        .ap_bram_114_addr1(ap_bram_iarg_114_addr1),
        .ap_bram_114_din1(ap_bram_iarg_114_din1),
        .ap_bram_114_dout1(ap_bram_iarg_114_dout1),
        .ap_bram_114_we1(ap_bram_iarg_114_we1),
        .ap_bram_114_en1(ap_bram_iarg_114_en1),
        .s_axis_bram_115_aclk(s_axis_bram_115_aclk),
        .s_axis_bram_115_aresetn(s_axis_bram_115_aresetn),
        .s_axis_bram_115_tlast(s_axis_bram_115_tlast),
        .s_axis_bram_115_tvalid(s_axis_bram_115_tvalid),
        .s_axis_bram_115_tkeep(s_axis_bram_115_tkeep),
        .s_axis_bram_115_tstrb(s_axis_bram_115_tstrb),
        .s_axis_bram_115_tdata(s_axis_bram_115_tdata),
        .s_axis_bram_115_tready(s_axis_bram_115_tready),
        .ap_bram_115_addr0(ap_bram_iarg_115_addr0),
        .ap_bram_115_din0(ap_bram_iarg_115_din0),
        .ap_bram_115_dout0(ap_bram_iarg_115_dout0),
        .ap_bram_115_we0(ap_bram_iarg_115_we0),
        .ap_bram_115_en0(ap_bram_iarg_115_en0),
        .ap_bram_115_addr1(ap_bram_iarg_115_addr1),
        .ap_bram_115_din1(ap_bram_iarg_115_din1),
        .ap_bram_115_dout1(ap_bram_iarg_115_dout1),
        .ap_bram_115_we1(ap_bram_iarg_115_we1),
        .ap_bram_115_en1(ap_bram_iarg_115_en1),
        .s_axis_bram_116_aclk(s_axis_bram_116_aclk),
        .s_axis_bram_116_aresetn(s_axis_bram_116_aresetn),
        .s_axis_bram_116_tlast(s_axis_bram_116_tlast),
        .s_axis_bram_116_tvalid(s_axis_bram_116_tvalid),
        .s_axis_bram_116_tkeep(s_axis_bram_116_tkeep),
        .s_axis_bram_116_tstrb(s_axis_bram_116_tstrb),
        .s_axis_bram_116_tdata(s_axis_bram_116_tdata),
        .s_axis_bram_116_tready(s_axis_bram_116_tready),
        .ap_bram_116_addr0(ap_bram_iarg_116_addr0),
        .ap_bram_116_din0(ap_bram_iarg_116_din0),
        .ap_bram_116_dout0(ap_bram_iarg_116_dout0),
        .ap_bram_116_we0(ap_bram_iarg_116_we0),
        .ap_bram_116_en0(ap_bram_iarg_116_en0),
        .ap_bram_116_addr1(ap_bram_iarg_116_addr1),
        .ap_bram_116_din1(ap_bram_iarg_116_din1),
        .ap_bram_116_dout1(ap_bram_iarg_116_dout1),
        .ap_bram_116_we1(ap_bram_iarg_116_we1),
        .ap_bram_116_en1(ap_bram_iarg_116_en1),
        .s_axis_bram_117_aclk(s_axis_bram_117_aclk),
        .s_axis_bram_117_aresetn(s_axis_bram_117_aresetn),
        .s_axis_bram_117_tlast(s_axis_bram_117_tlast),
        .s_axis_bram_117_tvalid(s_axis_bram_117_tvalid),
        .s_axis_bram_117_tkeep(s_axis_bram_117_tkeep),
        .s_axis_bram_117_tstrb(s_axis_bram_117_tstrb),
        .s_axis_bram_117_tdata(s_axis_bram_117_tdata),
        .s_axis_bram_117_tready(s_axis_bram_117_tready),
        .ap_bram_117_addr0(ap_bram_iarg_117_addr0),
        .ap_bram_117_din0(ap_bram_iarg_117_din0),
        .ap_bram_117_dout0(ap_bram_iarg_117_dout0),
        .ap_bram_117_we0(ap_bram_iarg_117_we0),
        .ap_bram_117_en0(ap_bram_iarg_117_en0),
        .ap_bram_117_addr1(ap_bram_iarg_117_addr1),
        .ap_bram_117_din1(ap_bram_iarg_117_din1),
        .ap_bram_117_dout1(ap_bram_iarg_117_dout1),
        .ap_bram_117_we1(ap_bram_iarg_117_we1),
        .ap_bram_117_en1(ap_bram_iarg_117_en1),
        .s_axis_bram_118_aclk(s_axis_bram_118_aclk),
        .s_axis_bram_118_aresetn(s_axis_bram_118_aresetn),
        .s_axis_bram_118_tlast(s_axis_bram_118_tlast),
        .s_axis_bram_118_tvalid(s_axis_bram_118_tvalid),
        .s_axis_bram_118_tkeep(s_axis_bram_118_tkeep),
        .s_axis_bram_118_tstrb(s_axis_bram_118_tstrb),
        .s_axis_bram_118_tdata(s_axis_bram_118_tdata),
        .s_axis_bram_118_tready(s_axis_bram_118_tready),
        .ap_bram_118_addr0(ap_bram_iarg_118_addr0),
        .ap_bram_118_din0(ap_bram_iarg_118_din0),
        .ap_bram_118_dout0(ap_bram_iarg_118_dout0),
        .ap_bram_118_we0(ap_bram_iarg_118_we0),
        .ap_bram_118_en0(ap_bram_iarg_118_en0),
        .ap_bram_118_addr1(ap_bram_iarg_118_addr1),
        .ap_bram_118_din1(ap_bram_iarg_118_din1),
        .ap_bram_118_dout1(ap_bram_iarg_118_dout1),
        .ap_bram_118_we1(ap_bram_iarg_118_we1),
        .ap_bram_118_en1(ap_bram_iarg_118_en1),
        .s_axis_bram_119_aclk(s_axis_bram_119_aclk),
        .s_axis_bram_119_aresetn(s_axis_bram_119_aresetn),
        .s_axis_bram_119_tlast(s_axis_bram_119_tlast),
        .s_axis_bram_119_tvalid(s_axis_bram_119_tvalid),
        .s_axis_bram_119_tkeep(s_axis_bram_119_tkeep),
        .s_axis_bram_119_tstrb(s_axis_bram_119_tstrb),
        .s_axis_bram_119_tdata(s_axis_bram_119_tdata),
        .s_axis_bram_119_tready(s_axis_bram_119_tready),
        .ap_bram_119_addr0(ap_bram_iarg_119_addr0),
        .ap_bram_119_din0(ap_bram_iarg_119_din0),
        .ap_bram_119_dout0(ap_bram_iarg_119_dout0),
        .ap_bram_119_we0(ap_bram_iarg_119_we0),
        .ap_bram_119_en0(ap_bram_iarg_119_en0),
        .ap_bram_119_addr1(ap_bram_iarg_119_addr1),
        .ap_bram_119_din1(ap_bram_iarg_119_din1),
        .ap_bram_119_dout1(ap_bram_iarg_119_dout1),
        .ap_bram_119_we1(ap_bram_iarg_119_we1),
        .ap_bram_119_en1(ap_bram_iarg_119_en1),
        .s_axis_bram_120_aclk(s_axis_bram_120_aclk),
        .s_axis_bram_120_aresetn(s_axis_bram_120_aresetn),
        .s_axis_bram_120_tlast(s_axis_bram_120_tlast),
        .s_axis_bram_120_tvalid(s_axis_bram_120_tvalid),
        .s_axis_bram_120_tkeep(s_axis_bram_120_tkeep),
        .s_axis_bram_120_tstrb(s_axis_bram_120_tstrb),
        .s_axis_bram_120_tdata(s_axis_bram_120_tdata),
        .s_axis_bram_120_tready(s_axis_bram_120_tready),
        .ap_bram_120_addr0(ap_bram_iarg_120_addr0),
        .ap_bram_120_din0(ap_bram_iarg_120_din0),
        .ap_bram_120_dout0(ap_bram_iarg_120_dout0),
        .ap_bram_120_we0(ap_bram_iarg_120_we0),
        .ap_bram_120_en0(ap_bram_iarg_120_en0),
        .ap_bram_120_addr1(ap_bram_iarg_120_addr1),
        .ap_bram_120_din1(ap_bram_iarg_120_din1),
        .ap_bram_120_dout1(ap_bram_iarg_120_dout1),
        .ap_bram_120_we1(ap_bram_iarg_120_we1),
        .ap_bram_120_en1(ap_bram_iarg_120_en1),
        .s_axis_bram_121_aclk(s_axis_bram_121_aclk),
        .s_axis_bram_121_aresetn(s_axis_bram_121_aresetn),
        .s_axis_bram_121_tlast(s_axis_bram_121_tlast),
        .s_axis_bram_121_tvalid(s_axis_bram_121_tvalid),
        .s_axis_bram_121_tkeep(s_axis_bram_121_tkeep),
        .s_axis_bram_121_tstrb(s_axis_bram_121_tstrb),
        .s_axis_bram_121_tdata(s_axis_bram_121_tdata),
        .s_axis_bram_121_tready(s_axis_bram_121_tready),
        .ap_bram_121_addr0(ap_bram_iarg_121_addr0),
        .ap_bram_121_din0(ap_bram_iarg_121_din0),
        .ap_bram_121_dout0(ap_bram_iarg_121_dout0),
        .ap_bram_121_we0(ap_bram_iarg_121_we0),
        .ap_bram_121_en0(ap_bram_iarg_121_en0),
        .ap_bram_121_addr1(ap_bram_iarg_121_addr1),
        .ap_bram_121_din1(ap_bram_iarg_121_din1),
        .ap_bram_121_dout1(ap_bram_iarg_121_dout1),
        .ap_bram_121_we1(ap_bram_iarg_121_we1),
        .ap_bram_121_en1(ap_bram_iarg_121_en1),
        .s_axis_bram_122_aclk(s_axis_bram_122_aclk),
        .s_axis_bram_122_aresetn(s_axis_bram_122_aresetn),
        .s_axis_bram_122_tlast(s_axis_bram_122_tlast),
        .s_axis_bram_122_tvalid(s_axis_bram_122_tvalid),
        .s_axis_bram_122_tkeep(s_axis_bram_122_tkeep),
        .s_axis_bram_122_tstrb(s_axis_bram_122_tstrb),
        .s_axis_bram_122_tdata(s_axis_bram_122_tdata),
        .s_axis_bram_122_tready(s_axis_bram_122_tready),
        .ap_bram_122_addr0(ap_bram_iarg_122_addr0),
        .ap_bram_122_din0(ap_bram_iarg_122_din0),
        .ap_bram_122_dout0(ap_bram_iarg_122_dout0),
        .ap_bram_122_we0(ap_bram_iarg_122_we0),
        .ap_bram_122_en0(ap_bram_iarg_122_en0),
        .ap_bram_122_addr1(ap_bram_iarg_122_addr1),
        .ap_bram_122_din1(ap_bram_iarg_122_din1),
        .ap_bram_122_dout1(ap_bram_iarg_122_dout1),
        .ap_bram_122_we1(ap_bram_iarg_122_we1),
        .ap_bram_122_en1(ap_bram_iarg_122_en1),
        .s_axis_bram_123_aclk(s_axis_bram_123_aclk),
        .s_axis_bram_123_aresetn(s_axis_bram_123_aresetn),
        .s_axis_bram_123_tlast(s_axis_bram_123_tlast),
        .s_axis_bram_123_tvalid(s_axis_bram_123_tvalid),
        .s_axis_bram_123_tkeep(s_axis_bram_123_tkeep),
        .s_axis_bram_123_tstrb(s_axis_bram_123_tstrb),
        .s_axis_bram_123_tdata(s_axis_bram_123_tdata),
        .s_axis_bram_123_tready(s_axis_bram_123_tready),
        .ap_bram_123_addr0(ap_bram_iarg_123_addr0),
        .ap_bram_123_din0(ap_bram_iarg_123_din0),
        .ap_bram_123_dout0(ap_bram_iarg_123_dout0),
        .ap_bram_123_we0(ap_bram_iarg_123_we0),
        .ap_bram_123_en0(ap_bram_iarg_123_en0),
        .ap_bram_123_addr1(ap_bram_iarg_123_addr1),
        .ap_bram_123_din1(ap_bram_iarg_123_din1),
        .ap_bram_123_dout1(ap_bram_iarg_123_dout1),
        .ap_bram_123_we1(ap_bram_iarg_123_we1),
        .ap_bram_123_en1(ap_bram_iarg_123_en1),
        .s_axis_bram_124_aclk(s_axis_bram_124_aclk),
        .s_axis_bram_124_aresetn(s_axis_bram_124_aresetn),
        .s_axis_bram_124_tlast(s_axis_bram_124_tlast),
        .s_axis_bram_124_tvalid(s_axis_bram_124_tvalid),
        .s_axis_bram_124_tkeep(s_axis_bram_124_tkeep),
        .s_axis_bram_124_tstrb(s_axis_bram_124_tstrb),
        .s_axis_bram_124_tdata(s_axis_bram_124_tdata),
        .s_axis_bram_124_tready(s_axis_bram_124_tready),
        .ap_bram_124_addr0(ap_bram_iarg_124_addr0),
        .ap_bram_124_din0(ap_bram_iarg_124_din0),
        .ap_bram_124_dout0(ap_bram_iarg_124_dout0),
        .ap_bram_124_we0(ap_bram_iarg_124_we0),
        .ap_bram_124_en0(ap_bram_iarg_124_en0),
        .ap_bram_124_addr1(ap_bram_iarg_124_addr1),
        .ap_bram_124_din1(ap_bram_iarg_124_din1),
        .ap_bram_124_dout1(ap_bram_iarg_124_dout1),
        .ap_bram_124_we1(ap_bram_iarg_124_we1),
        .ap_bram_124_en1(ap_bram_iarg_124_en1),
        .s_axis_bram_125_aclk(s_axis_bram_125_aclk),
        .s_axis_bram_125_aresetn(s_axis_bram_125_aresetn),
        .s_axis_bram_125_tlast(s_axis_bram_125_tlast),
        .s_axis_bram_125_tvalid(s_axis_bram_125_tvalid),
        .s_axis_bram_125_tkeep(s_axis_bram_125_tkeep),
        .s_axis_bram_125_tstrb(s_axis_bram_125_tstrb),
        .s_axis_bram_125_tdata(s_axis_bram_125_tdata),
        .s_axis_bram_125_tready(s_axis_bram_125_tready),
        .ap_bram_125_addr0(ap_bram_iarg_125_addr0),
        .ap_bram_125_din0(ap_bram_iarg_125_din0),
        .ap_bram_125_dout0(ap_bram_iarg_125_dout0),
        .ap_bram_125_we0(ap_bram_iarg_125_we0),
        .ap_bram_125_en0(ap_bram_iarg_125_en0),
        .ap_bram_125_addr1(ap_bram_iarg_125_addr1),
        .ap_bram_125_din1(ap_bram_iarg_125_din1),
        .ap_bram_125_dout1(ap_bram_iarg_125_dout1),
        .ap_bram_125_we1(ap_bram_iarg_125_we1),
        .ap_bram_125_en1(ap_bram_iarg_125_en1),
        .s_axis_bram_126_aclk(s_axis_bram_126_aclk),
        .s_axis_bram_126_aresetn(s_axis_bram_126_aresetn),
        .s_axis_bram_126_tlast(s_axis_bram_126_tlast),
        .s_axis_bram_126_tvalid(s_axis_bram_126_tvalid),
        .s_axis_bram_126_tkeep(s_axis_bram_126_tkeep),
        .s_axis_bram_126_tstrb(s_axis_bram_126_tstrb),
        .s_axis_bram_126_tdata(s_axis_bram_126_tdata),
        .s_axis_bram_126_tready(s_axis_bram_126_tready),
        .ap_bram_126_addr0(ap_bram_iarg_126_addr0),
        .ap_bram_126_din0(ap_bram_iarg_126_din0),
        .ap_bram_126_dout0(ap_bram_iarg_126_dout0),
        .ap_bram_126_we0(ap_bram_iarg_126_we0),
        .ap_bram_126_en0(ap_bram_iarg_126_en0),
        .ap_bram_126_addr1(ap_bram_iarg_126_addr1),
        .ap_bram_126_din1(ap_bram_iarg_126_din1),
        .ap_bram_126_dout1(ap_bram_iarg_126_dout1),
        .ap_bram_126_we1(ap_bram_iarg_126_we1),
        .ap_bram_126_en1(ap_bram_iarg_126_en1),
        .s_axis_bram_127_aclk(s_axis_bram_127_aclk),
        .s_axis_bram_127_aresetn(s_axis_bram_127_aresetn),
        .s_axis_bram_127_tlast(s_axis_bram_127_tlast),
        .s_axis_bram_127_tvalid(s_axis_bram_127_tvalid),
        .s_axis_bram_127_tkeep(s_axis_bram_127_tkeep),
        .s_axis_bram_127_tstrb(s_axis_bram_127_tstrb),
        .s_axis_bram_127_tdata(s_axis_bram_127_tdata),
        .s_axis_bram_127_tready(s_axis_bram_127_tready),
        .ap_bram_127_addr0(ap_bram_iarg_127_addr0),
        .ap_bram_127_din0(ap_bram_iarg_127_din0),
        .ap_bram_127_dout0(ap_bram_iarg_127_dout0),
        .ap_bram_127_we0(ap_bram_iarg_127_we0),
        .ap_bram_127_en0(ap_bram_iarg_127_en0),
        .ap_bram_127_addr1(ap_bram_iarg_127_addr1),
        .ap_bram_127_din1(ap_bram_iarg_127_din1),
        .ap_bram_127_dout1(ap_bram_iarg_127_dout1),
        .ap_bram_127_we1(ap_bram_iarg_127_we1),
        .ap_bram_127_en1(ap_bram_iarg_127_en1),
        .m_axis_bramio_0_aclk(m_axis_bramio_0_aclk),
        .m_axis_bramio_0_aresetn(m_axis_bramio_0_aresetn),
        .m_axis_bramio_0_tlast(m_axis_bramio_0_tlast),
        .m_axis_bramio_0_tvalid(m_axis_bramio_0_tvalid),
        .m_axis_bramio_0_tkeep(m_axis_bramio_0_tkeep),
        .m_axis_bramio_0_tstrb(m_axis_bramio_0_tstrb),
        .m_axis_bramio_0_tdata(m_axis_bramio_0_tdata),
        .m_axis_bramio_0_tready(m_axis_bramio_0_tready),
        .m_axis_bramio_1_aclk(m_axis_bramio_1_aclk),
        .m_axis_bramio_1_aresetn(m_axis_bramio_1_aresetn),
        .m_axis_bramio_1_tlast(m_axis_bramio_1_tlast),
        .m_axis_bramio_1_tvalid(m_axis_bramio_1_tvalid),
        .m_axis_bramio_1_tkeep(m_axis_bramio_1_tkeep),
        .m_axis_bramio_1_tstrb(m_axis_bramio_1_tstrb),
        .m_axis_bramio_1_tdata(m_axis_bramio_1_tdata),
        .m_axis_bramio_1_tready(m_axis_bramio_1_tready),
        .m_axis_bramio_2_aclk(m_axis_bramio_2_aclk),
        .m_axis_bramio_2_aresetn(m_axis_bramio_2_aresetn),
        .m_axis_bramio_2_tlast(m_axis_bramio_2_tlast),
        .m_axis_bramio_2_tvalid(m_axis_bramio_2_tvalid),
        .m_axis_bramio_2_tkeep(m_axis_bramio_2_tkeep),
        .m_axis_bramio_2_tstrb(m_axis_bramio_2_tstrb),
        .m_axis_bramio_2_tdata(m_axis_bramio_2_tdata),
        .m_axis_bramio_2_tready(m_axis_bramio_2_tready),
        .m_axis_bramio_3_aclk(m_axis_bramio_3_aclk),
        .m_axis_bramio_3_aresetn(m_axis_bramio_3_aresetn),
        .m_axis_bramio_3_tlast(m_axis_bramio_3_tlast),
        .m_axis_bramio_3_tvalid(m_axis_bramio_3_tvalid),
        .m_axis_bramio_3_tkeep(m_axis_bramio_3_tkeep),
        .m_axis_bramio_3_tstrb(m_axis_bramio_3_tstrb),
        .m_axis_bramio_3_tdata(m_axis_bramio_3_tdata),
        .m_axis_bramio_3_tready(m_axis_bramio_3_tready),
        .m_axis_bramio_4_aclk(m_axis_bramio_4_aclk),
        .m_axis_bramio_4_aresetn(m_axis_bramio_4_aresetn),
        .m_axis_bramio_4_tlast(m_axis_bramio_4_tlast),
        .m_axis_bramio_4_tvalid(m_axis_bramio_4_tvalid),
        .m_axis_bramio_4_tkeep(m_axis_bramio_4_tkeep),
        .m_axis_bramio_4_tstrb(m_axis_bramio_4_tstrb),
        .m_axis_bramio_4_tdata(m_axis_bramio_4_tdata),
        .m_axis_bramio_4_tready(m_axis_bramio_4_tready),
        .m_axis_bramio_5_aclk(m_axis_bramio_5_aclk),
        .m_axis_bramio_5_aresetn(m_axis_bramio_5_aresetn),
        .m_axis_bramio_5_tlast(m_axis_bramio_5_tlast),
        .m_axis_bramio_5_tvalid(m_axis_bramio_5_tvalid),
        .m_axis_bramio_5_tkeep(m_axis_bramio_5_tkeep),
        .m_axis_bramio_5_tstrb(m_axis_bramio_5_tstrb),
        .m_axis_bramio_5_tdata(m_axis_bramio_5_tdata),
        .m_axis_bramio_5_tready(m_axis_bramio_5_tready),
        .m_axis_bramio_6_aclk(m_axis_bramio_6_aclk),
        .m_axis_bramio_6_aresetn(m_axis_bramio_6_aresetn),
        .m_axis_bramio_6_tlast(m_axis_bramio_6_tlast),
        .m_axis_bramio_6_tvalid(m_axis_bramio_6_tvalid),
        .m_axis_bramio_6_tkeep(m_axis_bramio_6_tkeep),
        .m_axis_bramio_6_tstrb(m_axis_bramio_6_tstrb),
        .m_axis_bramio_6_tdata(m_axis_bramio_6_tdata),
        .m_axis_bramio_6_tready(m_axis_bramio_6_tready),
        .m_axis_bramio_7_aclk(m_axis_bramio_7_aclk),
        .m_axis_bramio_7_aresetn(m_axis_bramio_7_aresetn),
        .m_axis_bramio_7_tlast(m_axis_bramio_7_tlast),
        .m_axis_bramio_7_tvalid(m_axis_bramio_7_tvalid),
        .m_axis_bramio_7_tkeep(m_axis_bramio_7_tkeep),
        .m_axis_bramio_7_tstrb(m_axis_bramio_7_tstrb),
        .m_axis_bramio_7_tdata(m_axis_bramio_7_tdata),
        .m_axis_bramio_7_tready(m_axis_bramio_7_tready),
        .m_axis_bramio_8_aclk(m_axis_bramio_8_aclk),
        .m_axis_bramio_8_aresetn(m_axis_bramio_8_aresetn),
        .m_axis_bramio_8_tlast(m_axis_bramio_8_tlast),
        .m_axis_bramio_8_tvalid(m_axis_bramio_8_tvalid),
        .m_axis_bramio_8_tkeep(m_axis_bramio_8_tkeep),
        .m_axis_bramio_8_tstrb(m_axis_bramio_8_tstrb),
        .m_axis_bramio_8_tdata(m_axis_bramio_8_tdata),
        .m_axis_bramio_8_tready(m_axis_bramio_8_tready),
        .m_axis_bramio_9_aclk(m_axis_bramio_9_aclk),
        .m_axis_bramio_9_aresetn(m_axis_bramio_9_aresetn),
        .m_axis_bramio_9_tlast(m_axis_bramio_9_tlast),
        .m_axis_bramio_9_tvalid(m_axis_bramio_9_tvalid),
        .m_axis_bramio_9_tkeep(m_axis_bramio_9_tkeep),
        .m_axis_bramio_9_tstrb(m_axis_bramio_9_tstrb),
        .m_axis_bramio_9_tdata(m_axis_bramio_9_tdata),
        .m_axis_bramio_9_tready(m_axis_bramio_9_tready),
        .m_axis_bramio_10_aclk(m_axis_bramio_10_aclk),
        .m_axis_bramio_10_aresetn(m_axis_bramio_10_aresetn),
        .m_axis_bramio_10_tlast(m_axis_bramio_10_tlast),
        .m_axis_bramio_10_tvalid(m_axis_bramio_10_tvalid),
        .m_axis_bramio_10_tkeep(m_axis_bramio_10_tkeep),
        .m_axis_bramio_10_tstrb(m_axis_bramio_10_tstrb),
        .m_axis_bramio_10_tdata(m_axis_bramio_10_tdata),
        .m_axis_bramio_10_tready(m_axis_bramio_10_tready),
        .m_axis_bramio_11_aclk(m_axis_bramio_11_aclk),
        .m_axis_bramio_11_aresetn(m_axis_bramio_11_aresetn),
        .m_axis_bramio_11_tlast(m_axis_bramio_11_tlast),
        .m_axis_bramio_11_tvalid(m_axis_bramio_11_tvalid),
        .m_axis_bramio_11_tkeep(m_axis_bramio_11_tkeep),
        .m_axis_bramio_11_tstrb(m_axis_bramio_11_tstrb),
        .m_axis_bramio_11_tdata(m_axis_bramio_11_tdata),
        .m_axis_bramio_11_tready(m_axis_bramio_11_tready),
        .m_axis_bramio_12_aclk(m_axis_bramio_12_aclk),
        .m_axis_bramio_12_aresetn(m_axis_bramio_12_aresetn),
        .m_axis_bramio_12_tlast(m_axis_bramio_12_tlast),
        .m_axis_bramio_12_tvalid(m_axis_bramio_12_tvalid),
        .m_axis_bramio_12_tkeep(m_axis_bramio_12_tkeep),
        .m_axis_bramio_12_tstrb(m_axis_bramio_12_tstrb),
        .m_axis_bramio_12_tdata(m_axis_bramio_12_tdata),
        .m_axis_bramio_12_tready(m_axis_bramio_12_tready),
        .m_axis_bramio_13_aclk(m_axis_bramio_13_aclk),
        .m_axis_bramio_13_aresetn(m_axis_bramio_13_aresetn),
        .m_axis_bramio_13_tlast(m_axis_bramio_13_tlast),
        .m_axis_bramio_13_tvalid(m_axis_bramio_13_tvalid),
        .m_axis_bramio_13_tkeep(m_axis_bramio_13_tkeep),
        .m_axis_bramio_13_tstrb(m_axis_bramio_13_tstrb),
        .m_axis_bramio_13_tdata(m_axis_bramio_13_tdata),
        .m_axis_bramio_13_tready(m_axis_bramio_13_tready),
        .m_axis_bramio_14_aclk(m_axis_bramio_14_aclk),
        .m_axis_bramio_14_aresetn(m_axis_bramio_14_aresetn),
        .m_axis_bramio_14_tlast(m_axis_bramio_14_tlast),
        .m_axis_bramio_14_tvalid(m_axis_bramio_14_tvalid),
        .m_axis_bramio_14_tkeep(m_axis_bramio_14_tkeep),
        .m_axis_bramio_14_tstrb(m_axis_bramio_14_tstrb),
        .m_axis_bramio_14_tdata(m_axis_bramio_14_tdata),
        .m_axis_bramio_14_tready(m_axis_bramio_14_tready),
        .m_axis_bramio_15_aclk(m_axis_bramio_15_aclk),
        .m_axis_bramio_15_aresetn(m_axis_bramio_15_aresetn),
        .m_axis_bramio_15_tlast(m_axis_bramio_15_tlast),
        .m_axis_bramio_15_tvalid(m_axis_bramio_15_tvalid),
        .m_axis_bramio_15_tkeep(m_axis_bramio_15_tkeep),
        .m_axis_bramio_15_tstrb(m_axis_bramio_15_tstrb),
        .m_axis_bramio_15_tdata(m_axis_bramio_15_tdata),
        .m_axis_bramio_15_tready(m_axis_bramio_15_tready),
        .m_axis_bramio_16_aclk(m_axis_bramio_16_aclk),
        .m_axis_bramio_16_aresetn(m_axis_bramio_16_aresetn),
        .m_axis_bramio_16_tlast(m_axis_bramio_16_tlast),
        .m_axis_bramio_16_tvalid(m_axis_bramio_16_tvalid),
        .m_axis_bramio_16_tkeep(m_axis_bramio_16_tkeep),
        .m_axis_bramio_16_tstrb(m_axis_bramio_16_tstrb),
        .m_axis_bramio_16_tdata(m_axis_bramio_16_tdata),
        .m_axis_bramio_16_tready(m_axis_bramio_16_tready),
        .m_axis_bramio_17_aclk(m_axis_bramio_17_aclk),
        .m_axis_bramio_17_aresetn(m_axis_bramio_17_aresetn),
        .m_axis_bramio_17_tlast(m_axis_bramio_17_tlast),
        .m_axis_bramio_17_tvalid(m_axis_bramio_17_tvalid),
        .m_axis_bramio_17_tkeep(m_axis_bramio_17_tkeep),
        .m_axis_bramio_17_tstrb(m_axis_bramio_17_tstrb),
        .m_axis_bramio_17_tdata(m_axis_bramio_17_tdata),
        .m_axis_bramio_17_tready(m_axis_bramio_17_tready),
        .m_axis_bramio_18_aclk(m_axis_bramio_18_aclk),
        .m_axis_bramio_18_aresetn(m_axis_bramio_18_aresetn),
        .m_axis_bramio_18_tlast(m_axis_bramio_18_tlast),
        .m_axis_bramio_18_tvalid(m_axis_bramio_18_tvalid),
        .m_axis_bramio_18_tkeep(m_axis_bramio_18_tkeep),
        .m_axis_bramio_18_tstrb(m_axis_bramio_18_tstrb),
        .m_axis_bramio_18_tdata(m_axis_bramio_18_tdata),
        .m_axis_bramio_18_tready(m_axis_bramio_18_tready),
        .m_axis_bramio_19_aclk(m_axis_bramio_19_aclk),
        .m_axis_bramio_19_aresetn(m_axis_bramio_19_aresetn),
        .m_axis_bramio_19_tlast(m_axis_bramio_19_tlast),
        .m_axis_bramio_19_tvalid(m_axis_bramio_19_tvalid),
        .m_axis_bramio_19_tkeep(m_axis_bramio_19_tkeep),
        .m_axis_bramio_19_tstrb(m_axis_bramio_19_tstrb),
        .m_axis_bramio_19_tdata(m_axis_bramio_19_tdata),
        .m_axis_bramio_19_tready(m_axis_bramio_19_tready),
        .m_axis_bramio_20_aclk(m_axis_bramio_20_aclk),
        .m_axis_bramio_20_aresetn(m_axis_bramio_20_aresetn),
        .m_axis_bramio_20_tlast(m_axis_bramio_20_tlast),
        .m_axis_bramio_20_tvalid(m_axis_bramio_20_tvalid),
        .m_axis_bramio_20_tkeep(m_axis_bramio_20_tkeep),
        .m_axis_bramio_20_tstrb(m_axis_bramio_20_tstrb),
        .m_axis_bramio_20_tdata(m_axis_bramio_20_tdata),
        .m_axis_bramio_20_tready(m_axis_bramio_20_tready),
        .m_axis_bramio_21_aclk(m_axis_bramio_21_aclk),
        .m_axis_bramio_21_aresetn(m_axis_bramio_21_aresetn),
        .m_axis_bramio_21_tlast(m_axis_bramio_21_tlast),
        .m_axis_bramio_21_tvalid(m_axis_bramio_21_tvalid),
        .m_axis_bramio_21_tkeep(m_axis_bramio_21_tkeep),
        .m_axis_bramio_21_tstrb(m_axis_bramio_21_tstrb),
        .m_axis_bramio_21_tdata(m_axis_bramio_21_tdata),
        .m_axis_bramio_21_tready(m_axis_bramio_21_tready),
        .m_axis_bramio_22_aclk(m_axis_bramio_22_aclk),
        .m_axis_bramio_22_aresetn(m_axis_bramio_22_aresetn),
        .m_axis_bramio_22_tlast(m_axis_bramio_22_tlast),
        .m_axis_bramio_22_tvalid(m_axis_bramio_22_tvalid),
        .m_axis_bramio_22_tkeep(m_axis_bramio_22_tkeep),
        .m_axis_bramio_22_tstrb(m_axis_bramio_22_tstrb),
        .m_axis_bramio_22_tdata(m_axis_bramio_22_tdata),
        .m_axis_bramio_22_tready(m_axis_bramio_22_tready),
        .m_axis_bramio_23_aclk(m_axis_bramio_23_aclk),
        .m_axis_bramio_23_aresetn(m_axis_bramio_23_aresetn),
        .m_axis_bramio_23_tlast(m_axis_bramio_23_tlast),
        .m_axis_bramio_23_tvalid(m_axis_bramio_23_tvalid),
        .m_axis_bramio_23_tkeep(m_axis_bramio_23_tkeep),
        .m_axis_bramio_23_tstrb(m_axis_bramio_23_tstrb),
        .m_axis_bramio_23_tdata(m_axis_bramio_23_tdata),
        .m_axis_bramio_23_tready(m_axis_bramio_23_tready),
        .m_axis_bramio_24_aclk(m_axis_bramio_24_aclk),
        .m_axis_bramio_24_aresetn(m_axis_bramio_24_aresetn),
        .m_axis_bramio_24_tlast(m_axis_bramio_24_tlast),
        .m_axis_bramio_24_tvalid(m_axis_bramio_24_tvalid),
        .m_axis_bramio_24_tkeep(m_axis_bramio_24_tkeep),
        .m_axis_bramio_24_tstrb(m_axis_bramio_24_tstrb),
        .m_axis_bramio_24_tdata(m_axis_bramio_24_tdata),
        .m_axis_bramio_24_tready(m_axis_bramio_24_tready),
        .m_axis_bramio_25_aclk(m_axis_bramio_25_aclk),
        .m_axis_bramio_25_aresetn(m_axis_bramio_25_aresetn),
        .m_axis_bramio_25_tlast(m_axis_bramio_25_tlast),
        .m_axis_bramio_25_tvalid(m_axis_bramio_25_tvalid),
        .m_axis_bramio_25_tkeep(m_axis_bramio_25_tkeep),
        .m_axis_bramio_25_tstrb(m_axis_bramio_25_tstrb),
        .m_axis_bramio_25_tdata(m_axis_bramio_25_tdata),
        .m_axis_bramio_25_tready(m_axis_bramio_25_tready),
        .m_axis_bramio_26_aclk(m_axis_bramio_26_aclk),
        .m_axis_bramio_26_aresetn(m_axis_bramio_26_aresetn),
        .m_axis_bramio_26_tlast(m_axis_bramio_26_tlast),
        .m_axis_bramio_26_tvalid(m_axis_bramio_26_tvalid),
        .m_axis_bramio_26_tkeep(m_axis_bramio_26_tkeep),
        .m_axis_bramio_26_tstrb(m_axis_bramio_26_tstrb),
        .m_axis_bramio_26_tdata(m_axis_bramio_26_tdata),
        .m_axis_bramio_26_tready(m_axis_bramio_26_tready),
        .m_axis_bramio_27_aclk(m_axis_bramio_27_aclk),
        .m_axis_bramio_27_aresetn(m_axis_bramio_27_aresetn),
        .m_axis_bramio_27_tlast(m_axis_bramio_27_tlast),
        .m_axis_bramio_27_tvalid(m_axis_bramio_27_tvalid),
        .m_axis_bramio_27_tkeep(m_axis_bramio_27_tkeep),
        .m_axis_bramio_27_tstrb(m_axis_bramio_27_tstrb),
        .m_axis_bramio_27_tdata(m_axis_bramio_27_tdata),
        .m_axis_bramio_27_tready(m_axis_bramio_27_tready),
        .m_axis_bramio_28_aclk(m_axis_bramio_28_aclk),
        .m_axis_bramio_28_aresetn(m_axis_bramio_28_aresetn),
        .m_axis_bramio_28_tlast(m_axis_bramio_28_tlast),
        .m_axis_bramio_28_tvalid(m_axis_bramio_28_tvalid),
        .m_axis_bramio_28_tkeep(m_axis_bramio_28_tkeep),
        .m_axis_bramio_28_tstrb(m_axis_bramio_28_tstrb),
        .m_axis_bramio_28_tdata(m_axis_bramio_28_tdata),
        .m_axis_bramio_28_tready(m_axis_bramio_28_tready),
        .m_axis_bramio_29_aclk(m_axis_bramio_29_aclk),
        .m_axis_bramio_29_aresetn(m_axis_bramio_29_aresetn),
        .m_axis_bramio_29_tlast(m_axis_bramio_29_tlast),
        .m_axis_bramio_29_tvalid(m_axis_bramio_29_tvalid),
        .m_axis_bramio_29_tkeep(m_axis_bramio_29_tkeep),
        .m_axis_bramio_29_tstrb(m_axis_bramio_29_tstrb),
        .m_axis_bramio_29_tdata(m_axis_bramio_29_tdata),
        .m_axis_bramio_29_tready(m_axis_bramio_29_tready),
        .m_axis_bramio_30_aclk(m_axis_bramio_30_aclk),
        .m_axis_bramio_30_aresetn(m_axis_bramio_30_aresetn),
        .m_axis_bramio_30_tlast(m_axis_bramio_30_tlast),
        .m_axis_bramio_30_tvalid(m_axis_bramio_30_tvalid),
        .m_axis_bramio_30_tkeep(m_axis_bramio_30_tkeep),
        .m_axis_bramio_30_tstrb(m_axis_bramio_30_tstrb),
        .m_axis_bramio_30_tdata(m_axis_bramio_30_tdata),
        .m_axis_bramio_30_tready(m_axis_bramio_30_tready),
        .m_axis_bramio_31_aclk(m_axis_bramio_31_aclk),
        .m_axis_bramio_31_aresetn(m_axis_bramio_31_aresetn),
        .m_axis_bramio_31_tlast(m_axis_bramio_31_tlast),
        .m_axis_bramio_31_tvalid(m_axis_bramio_31_tvalid),
        .m_axis_bramio_31_tkeep(m_axis_bramio_31_tkeep),
        .m_axis_bramio_31_tstrb(m_axis_bramio_31_tstrb),
        .m_axis_bramio_31_tdata(m_axis_bramio_31_tdata),
        .m_axis_bramio_31_tready(m_axis_bramio_31_tready),
        .m_axis_bramio_32_aclk(m_axis_bramio_32_aclk),
        .m_axis_bramio_32_aresetn(m_axis_bramio_32_aresetn),
        .m_axis_bramio_32_tlast(m_axis_bramio_32_tlast),
        .m_axis_bramio_32_tvalid(m_axis_bramio_32_tvalid),
        .m_axis_bramio_32_tkeep(m_axis_bramio_32_tkeep),
        .m_axis_bramio_32_tstrb(m_axis_bramio_32_tstrb),
        .m_axis_bramio_32_tdata(m_axis_bramio_32_tdata),
        .m_axis_bramio_32_tready(m_axis_bramio_32_tready),
        .m_axis_bramio_33_aclk(m_axis_bramio_33_aclk),
        .m_axis_bramio_33_aresetn(m_axis_bramio_33_aresetn),
        .m_axis_bramio_33_tlast(m_axis_bramio_33_tlast),
        .m_axis_bramio_33_tvalid(m_axis_bramio_33_tvalid),
        .m_axis_bramio_33_tkeep(m_axis_bramio_33_tkeep),
        .m_axis_bramio_33_tstrb(m_axis_bramio_33_tstrb),
        .m_axis_bramio_33_tdata(m_axis_bramio_33_tdata),
        .m_axis_bramio_33_tready(m_axis_bramio_33_tready),
        .m_axis_bramio_34_aclk(m_axis_bramio_34_aclk),
        .m_axis_bramio_34_aresetn(m_axis_bramio_34_aresetn),
        .m_axis_bramio_34_tlast(m_axis_bramio_34_tlast),
        .m_axis_bramio_34_tvalid(m_axis_bramio_34_tvalid),
        .m_axis_bramio_34_tkeep(m_axis_bramio_34_tkeep),
        .m_axis_bramio_34_tstrb(m_axis_bramio_34_tstrb),
        .m_axis_bramio_34_tdata(m_axis_bramio_34_tdata),
        .m_axis_bramio_34_tready(m_axis_bramio_34_tready),
        .m_axis_bramio_35_aclk(m_axis_bramio_35_aclk),
        .m_axis_bramio_35_aresetn(m_axis_bramio_35_aresetn),
        .m_axis_bramio_35_tlast(m_axis_bramio_35_tlast),
        .m_axis_bramio_35_tvalid(m_axis_bramio_35_tvalid),
        .m_axis_bramio_35_tkeep(m_axis_bramio_35_tkeep),
        .m_axis_bramio_35_tstrb(m_axis_bramio_35_tstrb),
        .m_axis_bramio_35_tdata(m_axis_bramio_35_tdata),
        .m_axis_bramio_35_tready(m_axis_bramio_35_tready),
        .m_axis_bramio_36_aclk(m_axis_bramio_36_aclk),
        .m_axis_bramio_36_aresetn(m_axis_bramio_36_aresetn),
        .m_axis_bramio_36_tlast(m_axis_bramio_36_tlast),
        .m_axis_bramio_36_tvalid(m_axis_bramio_36_tvalid),
        .m_axis_bramio_36_tkeep(m_axis_bramio_36_tkeep),
        .m_axis_bramio_36_tstrb(m_axis_bramio_36_tstrb),
        .m_axis_bramio_36_tdata(m_axis_bramio_36_tdata),
        .m_axis_bramio_36_tready(m_axis_bramio_36_tready),
        .m_axis_bramio_37_aclk(m_axis_bramio_37_aclk),
        .m_axis_bramio_37_aresetn(m_axis_bramio_37_aresetn),
        .m_axis_bramio_37_tlast(m_axis_bramio_37_tlast),
        .m_axis_bramio_37_tvalid(m_axis_bramio_37_tvalid),
        .m_axis_bramio_37_tkeep(m_axis_bramio_37_tkeep),
        .m_axis_bramio_37_tstrb(m_axis_bramio_37_tstrb),
        .m_axis_bramio_37_tdata(m_axis_bramio_37_tdata),
        .m_axis_bramio_37_tready(m_axis_bramio_37_tready),
        .m_axis_bramio_38_aclk(m_axis_bramio_38_aclk),
        .m_axis_bramio_38_aresetn(m_axis_bramio_38_aresetn),
        .m_axis_bramio_38_tlast(m_axis_bramio_38_tlast),
        .m_axis_bramio_38_tvalid(m_axis_bramio_38_tvalid),
        .m_axis_bramio_38_tkeep(m_axis_bramio_38_tkeep),
        .m_axis_bramio_38_tstrb(m_axis_bramio_38_tstrb),
        .m_axis_bramio_38_tdata(m_axis_bramio_38_tdata),
        .m_axis_bramio_38_tready(m_axis_bramio_38_tready),
        .m_axis_bramio_39_aclk(m_axis_bramio_39_aclk),
        .m_axis_bramio_39_aresetn(m_axis_bramio_39_aresetn),
        .m_axis_bramio_39_tlast(m_axis_bramio_39_tlast),
        .m_axis_bramio_39_tvalid(m_axis_bramio_39_tvalid),
        .m_axis_bramio_39_tkeep(m_axis_bramio_39_tkeep),
        .m_axis_bramio_39_tstrb(m_axis_bramio_39_tstrb),
        .m_axis_bramio_39_tdata(m_axis_bramio_39_tdata),
        .m_axis_bramio_39_tready(m_axis_bramio_39_tready),
        .m_axis_bramio_40_aclk(m_axis_bramio_40_aclk),
        .m_axis_bramio_40_aresetn(m_axis_bramio_40_aresetn),
        .m_axis_bramio_40_tlast(m_axis_bramio_40_tlast),
        .m_axis_bramio_40_tvalid(m_axis_bramio_40_tvalid),
        .m_axis_bramio_40_tkeep(m_axis_bramio_40_tkeep),
        .m_axis_bramio_40_tstrb(m_axis_bramio_40_tstrb),
        .m_axis_bramio_40_tdata(m_axis_bramio_40_tdata),
        .m_axis_bramio_40_tready(m_axis_bramio_40_tready),
        .m_axis_bramio_41_aclk(m_axis_bramio_41_aclk),
        .m_axis_bramio_41_aresetn(m_axis_bramio_41_aresetn),
        .m_axis_bramio_41_tlast(m_axis_bramio_41_tlast),
        .m_axis_bramio_41_tvalid(m_axis_bramio_41_tvalid),
        .m_axis_bramio_41_tkeep(m_axis_bramio_41_tkeep),
        .m_axis_bramio_41_tstrb(m_axis_bramio_41_tstrb),
        .m_axis_bramio_41_tdata(m_axis_bramio_41_tdata),
        .m_axis_bramio_41_tready(m_axis_bramio_41_tready),
        .m_axis_bramio_42_aclk(m_axis_bramio_42_aclk),
        .m_axis_bramio_42_aresetn(m_axis_bramio_42_aresetn),
        .m_axis_bramio_42_tlast(m_axis_bramio_42_tlast),
        .m_axis_bramio_42_tvalid(m_axis_bramio_42_tvalid),
        .m_axis_bramio_42_tkeep(m_axis_bramio_42_tkeep),
        .m_axis_bramio_42_tstrb(m_axis_bramio_42_tstrb),
        .m_axis_bramio_42_tdata(m_axis_bramio_42_tdata),
        .m_axis_bramio_42_tready(m_axis_bramio_42_tready),
        .m_axis_bramio_43_aclk(m_axis_bramio_43_aclk),
        .m_axis_bramio_43_aresetn(m_axis_bramio_43_aresetn),
        .m_axis_bramio_43_tlast(m_axis_bramio_43_tlast),
        .m_axis_bramio_43_tvalid(m_axis_bramio_43_tvalid),
        .m_axis_bramio_43_tkeep(m_axis_bramio_43_tkeep),
        .m_axis_bramio_43_tstrb(m_axis_bramio_43_tstrb),
        .m_axis_bramio_43_tdata(m_axis_bramio_43_tdata),
        .m_axis_bramio_43_tready(m_axis_bramio_43_tready),
        .m_axis_bramio_44_aclk(m_axis_bramio_44_aclk),
        .m_axis_bramio_44_aresetn(m_axis_bramio_44_aresetn),
        .m_axis_bramio_44_tlast(m_axis_bramio_44_tlast),
        .m_axis_bramio_44_tvalid(m_axis_bramio_44_tvalid),
        .m_axis_bramio_44_tkeep(m_axis_bramio_44_tkeep),
        .m_axis_bramio_44_tstrb(m_axis_bramio_44_tstrb),
        .m_axis_bramio_44_tdata(m_axis_bramio_44_tdata),
        .m_axis_bramio_44_tready(m_axis_bramio_44_tready),
        .m_axis_bramio_45_aclk(m_axis_bramio_45_aclk),
        .m_axis_bramio_45_aresetn(m_axis_bramio_45_aresetn),
        .m_axis_bramio_45_tlast(m_axis_bramio_45_tlast),
        .m_axis_bramio_45_tvalid(m_axis_bramio_45_tvalid),
        .m_axis_bramio_45_tkeep(m_axis_bramio_45_tkeep),
        .m_axis_bramio_45_tstrb(m_axis_bramio_45_tstrb),
        .m_axis_bramio_45_tdata(m_axis_bramio_45_tdata),
        .m_axis_bramio_45_tready(m_axis_bramio_45_tready),
        .m_axis_bramio_46_aclk(m_axis_bramio_46_aclk),
        .m_axis_bramio_46_aresetn(m_axis_bramio_46_aresetn),
        .m_axis_bramio_46_tlast(m_axis_bramio_46_tlast),
        .m_axis_bramio_46_tvalid(m_axis_bramio_46_tvalid),
        .m_axis_bramio_46_tkeep(m_axis_bramio_46_tkeep),
        .m_axis_bramio_46_tstrb(m_axis_bramio_46_tstrb),
        .m_axis_bramio_46_tdata(m_axis_bramio_46_tdata),
        .m_axis_bramio_46_tready(m_axis_bramio_46_tready),
        .m_axis_bramio_47_aclk(m_axis_bramio_47_aclk),
        .m_axis_bramio_47_aresetn(m_axis_bramio_47_aresetn),
        .m_axis_bramio_47_tlast(m_axis_bramio_47_tlast),
        .m_axis_bramio_47_tvalid(m_axis_bramio_47_tvalid),
        .m_axis_bramio_47_tkeep(m_axis_bramio_47_tkeep),
        .m_axis_bramio_47_tstrb(m_axis_bramio_47_tstrb),
        .m_axis_bramio_47_tdata(m_axis_bramio_47_tdata),
        .m_axis_bramio_47_tready(m_axis_bramio_47_tready),
        .m_axis_bramio_48_aclk(m_axis_bramio_48_aclk),
        .m_axis_bramio_48_aresetn(m_axis_bramio_48_aresetn),
        .m_axis_bramio_48_tlast(m_axis_bramio_48_tlast),
        .m_axis_bramio_48_tvalid(m_axis_bramio_48_tvalid),
        .m_axis_bramio_48_tkeep(m_axis_bramio_48_tkeep),
        .m_axis_bramio_48_tstrb(m_axis_bramio_48_tstrb),
        .m_axis_bramio_48_tdata(m_axis_bramio_48_tdata),
        .m_axis_bramio_48_tready(m_axis_bramio_48_tready),
        .m_axis_bramio_49_aclk(m_axis_bramio_49_aclk),
        .m_axis_bramio_49_aresetn(m_axis_bramio_49_aresetn),
        .m_axis_bramio_49_tlast(m_axis_bramio_49_tlast),
        .m_axis_bramio_49_tvalid(m_axis_bramio_49_tvalid),
        .m_axis_bramio_49_tkeep(m_axis_bramio_49_tkeep),
        .m_axis_bramio_49_tstrb(m_axis_bramio_49_tstrb),
        .m_axis_bramio_49_tdata(m_axis_bramio_49_tdata),
        .m_axis_bramio_49_tready(m_axis_bramio_49_tready),
        .m_axis_bramio_50_aclk(m_axis_bramio_50_aclk),
        .m_axis_bramio_50_aresetn(m_axis_bramio_50_aresetn),
        .m_axis_bramio_50_tlast(m_axis_bramio_50_tlast),
        .m_axis_bramio_50_tvalid(m_axis_bramio_50_tvalid),
        .m_axis_bramio_50_tkeep(m_axis_bramio_50_tkeep),
        .m_axis_bramio_50_tstrb(m_axis_bramio_50_tstrb),
        .m_axis_bramio_50_tdata(m_axis_bramio_50_tdata),
        .m_axis_bramio_50_tready(m_axis_bramio_50_tready),
        .m_axis_bramio_51_aclk(m_axis_bramio_51_aclk),
        .m_axis_bramio_51_aresetn(m_axis_bramio_51_aresetn),
        .m_axis_bramio_51_tlast(m_axis_bramio_51_tlast),
        .m_axis_bramio_51_tvalid(m_axis_bramio_51_tvalid),
        .m_axis_bramio_51_tkeep(m_axis_bramio_51_tkeep),
        .m_axis_bramio_51_tstrb(m_axis_bramio_51_tstrb),
        .m_axis_bramio_51_tdata(m_axis_bramio_51_tdata),
        .m_axis_bramio_51_tready(m_axis_bramio_51_tready),
        .m_axis_bramio_52_aclk(m_axis_bramio_52_aclk),
        .m_axis_bramio_52_aresetn(m_axis_bramio_52_aresetn),
        .m_axis_bramio_52_tlast(m_axis_bramio_52_tlast),
        .m_axis_bramio_52_tvalid(m_axis_bramio_52_tvalid),
        .m_axis_bramio_52_tkeep(m_axis_bramio_52_tkeep),
        .m_axis_bramio_52_tstrb(m_axis_bramio_52_tstrb),
        .m_axis_bramio_52_tdata(m_axis_bramio_52_tdata),
        .m_axis_bramio_52_tready(m_axis_bramio_52_tready),
        .m_axis_bramio_53_aclk(m_axis_bramio_53_aclk),
        .m_axis_bramio_53_aresetn(m_axis_bramio_53_aresetn),
        .m_axis_bramio_53_tlast(m_axis_bramio_53_tlast),
        .m_axis_bramio_53_tvalid(m_axis_bramio_53_tvalid),
        .m_axis_bramio_53_tkeep(m_axis_bramio_53_tkeep),
        .m_axis_bramio_53_tstrb(m_axis_bramio_53_tstrb),
        .m_axis_bramio_53_tdata(m_axis_bramio_53_tdata),
        .m_axis_bramio_53_tready(m_axis_bramio_53_tready),
        .m_axis_bramio_54_aclk(m_axis_bramio_54_aclk),
        .m_axis_bramio_54_aresetn(m_axis_bramio_54_aresetn),
        .m_axis_bramio_54_tlast(m_axis_bramio_54_tlast),
        .m_axis_bramio_54_tvalid(m_axis_bramio_54_tvalid),
        .m_axis_bramio_54_tkeep(m_axis_bramio_54_tkeep),
        .m_axis_bramio_54_tstrb(m_axis_bramio_54_tstrb),
        .m_axis_bramio_54_tdata(m_axis_bramio_54_tdata),
        .m_axis_bramio_54_tready(m_axis_bramio_54_tready),
        .m_axis_bramio_55_aclk(m_axis_bramio_55_aclk),
        .m_axis_bramio_55_aresetn(m_axis_bramio_55_aresetn),
        .m_axis_bramio_55_tlast(m_axis_bramio_55_tlast),
        .m_axis_bramio_55_tvalid(m_axis_bramio_55_tvalid),
        .m_axis_bramio_55_tkeep(m_axis_bramio_55_tkeep),
        .m_axis_bramio_55_tstrb(m_axis_bramio_55_tstrb),
        .m_axis_bramio_55_tdata(m_axis_bramio_55_tdata),
        .m_axis_bramio_55_tready(m_axis_bramio_55_tready),
        .m_axis_bramio_56_aclk(m_axis_bramio_56_aclk),
        .m_axis_bramio_56_aresetn(m_axis_bramio_56_aresetn),
        .m_axis_bramio_56_tlast(m_axis_bramio_56_tlast),
        .m_axis_bramio_56_tvalid(m_axis_bramio_56_tvalid),
        .m_axis_bramio_56_tkeep(m_axis_bramio_56_tkeep),
        .m_axis_bramio_56_tstrb(m_axis_bramio_56_tstrb),
        .m_axis_bramio_56_tdata(m_axis_bramio_56_tdata),
        .m_axis_bramio_56_tready(m_axis_bramio_56_tready),
        .m_axis_bramio_57_aclk(m_axis_bramio_57_aclk),
        .m_axis_bramio_57_aresetn(m_axis_bramio_57_aresetn),
        .m_axis_bramio_57_tlast(m_axis_bramio_57_tlast),
        .m_axis_bramio_57_tvalid(m_axis_bramio_57_tvalid),
        .m_axis_bramio_57_tkeep(m_axis_bramio_57_tkeep),
        .m_axis_bramio_57_tstrb(m_axis_bramio_57_tstrb),
        .m_axis_bramio_57_tdata(m_axis_bramio_57_tdata),
        .m_axis_bramio_57_tready(m_axis_bramio_57_tready),
        .m_axis_bramio_58_aclk(m_axis_bramio_58_aclk),
        .m_axis_bramio_58_aresetn(m_axis_bramio_58_aresetn),
        .m_axis_bramio_58_tlast(m_axis_bramio_58_tlast),
        .m_axis_bramio_58_tvalid(m_axis_bramio_58_tvalid),
        .m_axis_bramio_58_tkeep(m_axis_bramio_58_tkeep),
        .m_axis_bramio_58_tstrb(m_axis_bramio_58_tstrb),
        .m_axis_bramio_58_tdata(m_axis_bramio_58_tdata),
        .m_axis_bramio_58_tready(m_axis_bramio_58_tready),
        .m_axis_bramio_59_aclk(m_axis_bramio_59_aclk),
        .m_axis_bramio_59_aresetn(m_axis_bramio_59_aresetn),
        .m_axis_bramio_59_tlast(m_axis_bramio_59_tlast),
        .m_axis_bramio_59_tvalid(m_axis_bramio_59_tvalid),
        .m_axis_bramio_59_tkeep(m_axis_bramio_59_tkeep),
        .m_axis_bramio_59_tstrb(m_axis_bramio_59_tstrb),
        .m_axis_bramio_59_tdata(m_axis_bramio_59_tdata),
        .m_axis_bramio_59_tready(m_axis_bramio_59_tready),
        .m_axis_bramio_60_aclk(m_axis_bramio_60_aclk),
        .m_axis_bramio_60_aresetn(m_axis_bramio_60_aresetn),
        .m_axis_bramio_60_tlast(m_axis_bramio_60_tlast),
        .m_axis_bramio_60_tvalid(m_axis_bramio_60_tvalid),
        .m_axis_bramio_60_tkeep(m_axis_bramio_60_tkeep),
        .m_axis_bramio_60_tstrb(m_axis_bramio_60_tstrb),
        .m_axis_bramio_60_tdata(m_axis_bramio_60_tdata),
        .m_axis_bramio_60_tready(m_axis_bramio_60_tready),
        .m_axis_bramio_61_aclk(m_axis_bramio_61_aclk),
        .m_axis_bramio_61_aresetn(m_axis_bramio_61_aresetn),
        .m_axis_bramio_61_tlast(m_axis_bramio_61_tlast),
        .m_axis_bramio_61_tvalid(m_axis_bramio_61_tvalid),
        .m_axis_bramio_61_tkeep(m_axis_bramio_61_tkeep),
        .m_axis_bramio_61_tstrb(m_axis_bramio_61_tstrb),
        .m_axis_bramio_61_tdata(m_axis_bramio_61_tdata),
        .m_axis_bramio_61_tready(m_axis_bramio_61_tready),
        .m_axis_bramio_62_aclk(m_axis_bramio_62_aclk),
        .m_axis_bramio_62_aresetn(m_axis_bramio_62_aresetn),
        .m_axis_bramio_62_tlast(m_axis_bramio_62_tlast),
        .m_axis_bramio_62_tvalid(m_axis_bramio_62_tvalid),
        .m_axis_bramio_62_tkeep(m_axis_bramio_62_tkeep),
        .m_axis_bramio_62_tstrb(m_axis_bramio_62_tstrb),
        .m_axis_bramio_62_tdata(m_axis_bramio_62_tdata),
        .m_axis_bramio_62_tready(m_axis_bramio_62_tready),
        .m_axis_bramio_63_aclk(m_axis_bramio_63_aclk),
        .m_axis_bramio_63_aresetn(m_axis_bramio_63_aresetn),
        .m_axis_bramio_63_tlast(m_axis_bramio_63_tlast),
        .m_axis_bramio_63_tvalid(m_axis_bramio_63_tvalid),
        .m_axis_bramio_63_tkeep(m_axis_bramio_63_tkeep),
        .m_axis_bramio_63_tstrb(m_axis_bramio_63_tstrb),
        .m_axis_bramio_63_tdata(m_axis_bramio_63_tdata),
        .m_axis_bramio_63_tready(m_axis_bramio_63_tready),
        .m_axis_bramio_64_aclk(m_axis_bramio_64_aclk),
        .m_axis_bramio_64_aresetn(m_axis_bramio_64_aresetn),
        .m_axis_bramio_64_tlast(m_axis_bramio_64_tlast),
        .m_axis_bramio_64_tvalid(m_axis_bramio_64_tvalid),
        .m_axis_bramio_64_tkeep(m_axis_bramio_64_tkeep),
        .m_axis_bramio_64_tstrb(m_axis_bramio_64_tstrb),
        .m_axis_bramio_64_tdata(m_axis_bramio_64_tdata),
        .m_axis_bramio_64_tready(m_axis_bramio_64_tready),
        .m_axis_bramio_65_aclk(m_axis_bramio_65_aclk),
        .m_axis_bramio_65_aresetn(m_axis_bramio_65_aresetn),
        .m_axis_bramio_65_tlast(m_axis_bramio_65_tlast),
        .m_axis_bramio_65_tvalid(m_axis_bramio_65_tvalid),
        .m_axis_bramio_65_tkeep(m_axis_bramio_65_tkeep),
        .m_axis_bramio_65_tstrb(m_axis_bramio_65_tstrb),
        .m_axis_bramio_65_tdata(m_axis_bramio_65_tdata),
        .m_axis_bramio_65_tready(m_axis_bramio_65_tready),
        .m_axis_bramio_66_aclk(m_axis_bramio_66_aclk),
        .m_axis_bramio_66_aresetn(m_axis_bramio_66_aresetn),
        .m_axis_bramio_66_tlast(m_axis_bramio_66_tlast),
        .m_axis_bramio_66_tvalid(m_axis_bramio_66_tvalid),
        .m_axis_bramio_66_tkeep(m_axis_bramio_66_tkeep),
        .m_axis_bramio_66_tstrb(m_axis_bramio_66_tstrb),
        .m_axis_bramio_66_tdata(m_axis_bramio_66_tdata),
        .m_axis_bramio_66_tready(m_axis_bramio_66_tready),
        .m_axis_bramio_67_aclk(m_axis_bramio_67_aclk),
        .m_axis_bramio_67_aresetn(m_axis_bramio_67_aresetn),
        .m_axis_bramio_67_tlast(m_axis_bramio_67_tlast),
        .m_axis_bramio_67_tvalid(m_axis_bramio_67_tvalid),
        .m_axis_bramio_67_tkeep(m_axis_bramio_67_tkeep),
        .m_axis_bramio_67_tstrb(m_axis_bramio_67_tstrb),
        .m_axis_bramio_67_tdata(m_axis_bramio_67_tdata),
        .m_axis_bramio_67_tready(m_axis_bramio_67_tready),
        .m_axis_bramio_68_aclk(m_axis_bramio_68_aclk),
        .m_axis_bramio_68_aresetn(m_axis_bramio_68_aresetn),
        .m_axis_bramio_68_tlast(m_axis_bramio_68_tlast),
        .m_axis_bramio_68_tvalid(m_axis_bramio_68_tvalid),
        .m_axis_bramio_68_tkeep(m_axis_bramio_68_tkeep),
        .m_axis_bramio_68_tstrb(m_axis_bramio_68_tstrb),
        .m_axis_bramio_68_tdata(m_axis_bramio_68_tdata),
        .m_axis_bramio_68_tready(m_axis_bramio_68_tready),
        .m_axis_bramio_69_aclk(m_axis_bramio_69_aclk),
        .m_axis_bramio_69_aresetn(m_axis_bramio_69_aresetn),
        .m_axis_bramio_69_tlast(m_axis_bramio_69_tlast),
        .m_axis_bramio_69_tvalid(m_axis_bramio_69_tvalid),
        .m_axis_bramio_69_tkeep(m_axis_bramio_69_tkeep),
        .m_axis_bramio_69_tstrb(m_axis_bramio_69_tstrb),
        .m_axis_bramio_69_tdata(m_axis_bramio_69_tdata),
        .m_axis_bramio_69_tready(m_axis_bramio_69_tready),
        .m_axis_bramio_70_aclk(m_axis_bramio_70_aclk),
        .m_axis_bramio_70_aresetn(m_axis_bramio_70_aresetn),
        .m_axis_bramio_70_tlast(m_axis_bramio_70_tlast),
        .m_axis_bramio_70_tvalid(m_axis_bramio_70_tvalid),
        .m_axis_bramio_70_tkeep(m_axis_bramio_70_tkeep),
        .m_axis_bramio_70_tstrb(m_axis_bramio_70_tstrb),
        .m_axis_bramio_70_tdata(m_axis_bramio_70_tdata),
        .m_axis_bramio_70_tready(m_axis_bramio_70_tready),
        .m_axis_bramio_71_aclk(m_axis_bramio_71_aclk),
        .m_axis_bramio_71_aresetn(m_axis_bramio_71_aresetn),
        .m_axis_bramio_71_tlast(m_axis_bramio_71_tlast),
        .m_axis_bramio_71_tvalid(m_axis_bramio_71_tvalid),
        .m_axis_bramio_71_tkeep(m_axis_bramio_71_tkeep),
        .m_axis_bramio_71_tstrb(m_axis_bramio_71_tstrb),
        .m_axis_bramio_71_tdata(m_axis_bramio_71_tdata),
        .m_axis_bramio_71_tready(m_axis_bramio_71_tready),
        .m_axis_bramio_72_aclk(m_axis_bramio_72_aclk),
        .m_axis_bramio_72_aresetn(m_axis_bramio_72_aresetn),
        .m_axis_bramio_72_tlast(m_axis_bramio_72_tlast),
        .m_axis_bramio_72_tvalid(m_axis_bramio_72_tvalid),
        .m_axis_bramio_72_tkeep(m_axis_bramio_72_tkeep),
        .m_axis_bramio_72_tstrb(m_axis_bramio_72_tstrb),
        .m_axis_bramio_72_tdata(m_axis_bramio_72_tdata),
        .m_axis_bramio_72_tready(m_axis_bramio_72_tready),
        .m_axis_bramio_73_aclk(m_axis_bramio_73_aclk),
        .m_axis_bramio_73_aresetn(m_axis_bramio_73_aresetn),
        .m_axis_bramio_73_tlast(m_axis_bramio_73_tlast),
        .m_axis_bramio_73_tvalid(m_axis_bramio_73_tvalid),
        .m_axis_bramio_73_tkeep(m_axis_bramio_73_tkeep),
        .m_axis_bramio_73_tstrb(m_axis_bramio_73_tstrb),
        .m_axis_bramio_73_tdata(m_axis_bramio_73_tdata),
        .m_axis_bramio_73_tready(m_axis_bramio_73_tready),
        .m_axis_bramio_74_aclk(m_axis_bramio_74_aclk),
        .m_axis_bramio_74_aresetn(m_axis_bramio_74_aresetn),
        .m_axis_bramio_74_tlast(m_axis_bramio_74_tlast),
        .m_axis_bramio_74_tvalid(m_axis_bramio_74_tvalid),
        .m_axis_bramio_74_tkeep(m_axis_bramio_74_tkeep),
        .m_axis_bramio_74_tstrb(m_axis_bramio_74_tstrb),
        .m_axis_bramio_74_tdata(m_axis_bramio_74_tdata),
        .m_axis_bramio_74_tready(m_axis_bramio_74_tready),
        .m_axis_bramio_75_aclk(m_axis_bramio_75_aclk),
        .m_axis_bramio_75_aresetn(m_axis_bramio_75_aresetn),
        .m_axis_bramio_75_tlast(m_axis_bramio_75_tlast),
        .m_axis_bramio_75_tvalid(m_axis_bramio_75_tvalid),
        .m_axis_bramio_75_tkeep(m_axis_bramio_75_tkeep),
        .m_axis_bramio_75_tstrb(m_axis_bramio_75_tstrb),
        .m_axis_bramio_75_tdata(m_axis_bramio_75_tdata),
        .m_axis_bramio_75_tready(m_axis_bramio_75_tready),
        .m_axis_bramio_76_aclk(m_axis_bramio_76_aclk),
        .m_axis_bramio_76_aresetn(m_axis_bramio_76_aresetn),
        .m_axis_bramio_76_tlast(m_axis_bramio_76_tlast),
        .m_axis_bramio_76_tvalid(m_axis_bramio_76_tvalid),
        .m_axis_bramio_76_tkeep(m_axis_bramio_76_tkeep),
        .m_axis_bramio_76_tstrb(m_axis_bramio_76_tstrb),
        .m_axis_bramio_76_tdata(m_axis_bramio_76_tdata),
        .m_axis_bramio_76_tready(m_axis_bramio_76_tready),
        .m_axis_bramio_77_aclk(m_axis_bramio_77_aclk),
        .m_axis_bramio_77_aresetn(m_axis_bramio_77_aresetn),
        .m_axis_bramio_77_tlast(m_axis_bramio_77_tlast),
        .m_axis_bramio_77_tvalid(m_axis_bramio_77_tvalid),
        .m_axis_bramio_77_tkeep(m_axis_bramio_77_tkeep),
        .m_axis_bramio_77_tstrb(m_axis_bramio_77_tstrb),
        .m_axis_bramio_77_tdata(m_axis_bramio_77_tdata),
        .m_axis_bramio_77_tready(m_axis_bramio_77_tready),
        .m_axis_bramio_78_aclk(m_axis_bramio_78_aclk),
        .m_axis_bramio_78_aresetn(m_axis_bramio_78_aresetn),
        .m_axis_bramio_78_tlast(m_axis_bramio_78_tlast),
        .m_axis_bramio_78_tvalid(m_axis_bramio_78_tvalid),
        .m_axis_bramio_78_tkeep(m_axis_bramio_78_tkeep),
        .m_axis_bramio_78_tstrb(m_axis_bramio_78_tstrb),
        .m_axis_bramio_78_tdata(m_axis_bramio_78_tdata),
        .m_axis_bramio_78_tready(m_axis_bramio_78_tready),
        .m_axis_bramio_79_aclk(m_axis_bramio_79_aclk),
        .m_axis_bramio_79_aresetn(m_axis_bramio_79_aresetn),
        .m_axis_bramio_79_tlast(m_axis_bramio_79_tlast),
        .m_axis_bramio_79_tvalid(m_axis_bramio_79_tvalid),
        .m_axis_bramio_79_tkeep(m_axis_bramio_79_tkeep),
        .m_axis_bramio_79_tstrb(m_axis_bramio_79_tstrb),
        .m_axis_bramio_79_tdata(m_axis_bramio_79_tdata),
        .m_axis_bramio_79_tready(m_axis_bramio_79_tready),
        .m_axis_bramio_80_aclk(m_axis_bramio_80_aclk),
        .m_axis_bramio_80_aresetn(m_axis_bramio_80_aresetn),
        .m_axis_bramio_80_tlast(m_axis_bramio_80_tlast),
        .m_axis_bramio_80_tvalid(m_axis_bramio_80_tvalid),
        .m_axis_bramio_80_tkeep(m_axis_bramio_80_tkeep),
        .m_axis_bramio_80_tstrb(m_axis_bramio_80_tstrb),
        .m_axis_bramio_80_tdata(m_axis_bramio_80_tdata),
        .m_axis_bramio_80_tready(m_axis_bramio_80_tready),
        .m_axis_bramio_81_aclk(m_axis_bramio_81_aclk),
        .m_axis_bramio_81_aresetn(m_axis_bramio_81_aresetn),
        .m_axis_bramio_81_tlast(m_axis_bramio_81_tlast),
        .m_axis_bramio_81_tvalid(m_axis_bramio_81_tvalid),
        .m_axis_bramio_81_tkeep(m_axis_bramio_81_tkeep),
        .m_axis_bramio_81_tstrb(m_axis_bramio_81_tstrb),
        .m_axis_bramio_81_tdata(m_axis_bramio_81_tdata),
        .m_axis_bramio_81_tready(m_axis_bramio_81_tready),
        .m_axis_bramio_82_aclk(m_axis_bramio_82_aclk),
        .m_axis_bramio_82_aresetn(m_axis_bramio_82_aresetn),
        .m_axis_bramio_82_tlast(m_axis_bramio_82_tlast),
        .m_axis_bramio_82_tvalid(m_axis_bramio_82_tvalid),
        .m_axis_bramio_82_tkeep(m_axis_bramio_82_tkeep),
        .m_axis_bramio_82_tstrb(m_axis_bramio_82_tstrb),
        .m_axis_bramio_82_tdata(m_axis_bramio_82_tdata),
        .m_axis_bramio_82_tready(m_axis_bramio_82_tready),
        .m_axis_bramio_83_aclk(m_axis_bramio_83_aclk),
        .m_axis_bramio_83_aresetn(m_axis_bramio_83_aresetn),
        .m_axis_bramio_83_tlast(m_axis_bramio_83_tlast),
        .m_axis_bramio_83_tvalid(m_axis_bramio_83_tvalid),
        .m_axis_bramio_83_tkeep(m_axis_bramio_83_tkeep),
        .m_axis_bramio_83_tstrb(m_axis_bramio_83_tstrb),
        .m_axis_bramio_83_tdata(m_axis_bramio_83_tdata),
        .m_axis_bramio_83_tready(m_axis_bramio_83_tready),
        .m_axis_bramio_84_aclk(m_axis_bramio_84_aclk),
        .m_axis_bramio_84_aresetn(m_axis_bramio_84_aresetn),
        .m_axis_bramio_84_tlast(m_axis_bramio_84_tlast),
        .m_axis_bramio_84_tvalid(m_axis_bramio_84_tvalid),
        .m_axis_bramio_84_tkeep(m_axis_bramio_84_tkeep),
        .m_axis_bramio_84_tstrb(m_axis_bramio_84_tstrb),
        .m_axis_bramio_84_tdata(m_axis_bramio_84_tdata),
        .m_axis_bramio_84_tready(m_axis_bramio_84_tready),
        .m_axis_bramio_85_aclk(m_axis_bramio_85_aclk),
        .m_axis_bramio_85_aresetn(m_axis_bramio_85_aresetn),
        .m_axis_bramio_85_tlast(m_axis_bramio_85_tlast),
        .m_axis_bramio_85_tvalid(m_axis_bramio_85_tvalid),
        .m_axis_bramio_85_tkeep(m_axis_bramio_85_tkeep),
        .m_axis_bramio_85_tstrb(m_axis_bramio_85_tstrb),
        .m_axis_bramio_85_tdata(m_axis_bramio_85_tdata),
        .m_axis_bramio_85_tready(m_axis_bramio_85_tready),
        .m_axis_bramio_86_aclk(m_axis_bramio_86_aclk),
        .m_axis_bramio_86_aresetn(m_axis_bramio_86_aresetn),
        .m_axis_bramio_86_tlast(m_axis_bramio_86_tlast),
        .m_axis_bramio_86_tvalid(m_axis_bramio_86_tvalid),
        .m_axis_bramio_86_tkeep(m_axis_bramio_86_tkeep),
        .m_axis_bramio_86_tstrb(m_axis_bramio_86_tstrb),
        .m_axis_bramio_86_tdata(m_axis_bramio_86_tdata),
        .m_axis_bramio_86_tready(m_axis_bramio_86_tready),
        .m_axis_bramio_87_aclk(m_axis_bramio_87_aclk),
        .m_axis_bramio_87_aresetn(m_axis_bramio_87_aresetn),
        .m_axis_bramio_87_tlast(m_axis_bramio_87_tlast),
        .m_axis_bramio_87_tvalid(m_axis_bramio_87_tvalid),
        .m_axis_bramio_87_tkeep(m_axis_bramio_87_tkeep),
        .m_axis_bramio_87_tstrb(m_axis_bramio_87_tstrb),
        .m_axis_bramio_87_tdata(m_axis_bramio_87_tdata),
        .m_axis_bramio_87_tready(m_axis_bramio_87_tready),
        .m_axis_bramio_88_aclk(m_axis_bramio_88_aclk),
        .m_axis_bramio_88_aresetn(m_axis_bramio_88_aresetn),
        .m_axis_bramio_88_tlast(m_axis_bramio_88_tlast),
        .m_axis_bramio_88_tvalid(m_axis_bramio_88_tvalid),
        .m_axis_bramio_88_tkeep(m_axis_bramio_88_tkeep),
        .m_axis_bramio_88_tstrb(m_axis_bramio_88_tstrb),
        .m_axis_bramio_88_tdata(m_axis_bramio_88_tdata),
        .m_axis_bramio_88_tready(m_axis_bramio_88_tready),
        .m_axis_bramio_89_aclk(m_axis_bramio_89_aclk),
        .m_axis_bramio_89_aresetn(m_axis_bramio_89_aresetn),
        .m_axis_bramio_89_tlast(m_axis_bramio_89_tlast),
        .m_axis_bramio_89_tvalid(m_axis_bramio_89_tvalid),
        .m_axis_bramio_89_tkeep(m_axis_bramio_89_tkeep),
        .m_axis_bramio_89_tstrb(m_axis_bramio_89_tstrb),
        .m_axis_bramio_89_tdata(m_axis_bramio_89_tdata),
        .m_axis_bramio_89_tready(m_axis_bramio_89_tready),
        .m_axis_bramio_90_aclk(m_axis_bramio_90_aclk),
        .m_axis_bramio_90_aresetn(m_axis_bramio_90_aresetn),
        .m_axis_bramio_90_tlast(m_axis_bramio_90_tlast),
        .m_axis_bramio_90_tvalid(m_axis_bramio_90_tvalid),
        .m_axis_bramio_90_tkeep(m_axis_bramio_90_tkeep),
        .m_axis_bramio_90_tstrb(m_axis_bramio_90_tstrb),
        .m_axis_bramio_90_tdata(m_axis_bramio_90_tdata),
        .m_axis_bramio_90_tready(m_axis_bramio_90_tready),
        .m_axis_bramio_91_aclk(m_axis_bramio_91_aclk),
        .m_axis_bramio_91_aresetn(m_axis_bramio_91_aresetn),
        .m_axis_bramio_91_tlast(m_axis_bramio_91_tlast),
        .m_axis_bramio_91_tvalid(m_axis_bramio_91_tvalid),
        .m_axis_bramio_91_tkeep(m_axis_bramio_91_tkeep),
        .m_axis_bramio_91_tstrb(m_axis_bramio_91_tstrb),
        .m_axis_bramio_91_tdata(m_axis_bramio_91_tdata),
        .m_axis_bramio_91_tready(m_axis_bramio_91_tready),
        .m_axis_bramio_92_aclk(m_axis_bramio_92_aclk),
        .m_axis_bramio_92_aresetn(m_axis_bramio_92_aresetn),
        .m_axis_bramio_92_tlast(m_axis_bramio_92_tlast),
        .m_axis_bramio_92_tvalid(m_axis_bramio_92_tvalid),
        .m_axis_bramio_92_tkeep(m_axis_bramio_92_tkeep),
        .m_axis_bramio_92_tstrb(m_axis_bramio_92_tstrb),
        .m_axis_bramio_92_tdata(m_axis_bramio_92_tdata),
        .m_axis_bramio_92_tready(m_axis_bramio_92_tready),
        .m_axis_bramio_93_aclk(m_axis_bramio_93_aclk),
        .m_axis_bramio_93_aresetn(m_axis_bramio_93_aresetn),
        .m_axis_bramio_93_tlast(m_axis_bramio_93_tlast),
        .m_axis_bramio_93_tvalid(m_axis_bramio_93_tvalid),
        .m_axis_bramio_93_tkeep(m_axis_bramio_93_tkeep),
        .m_axis_bramio_93_tstrb(m_axis_bramio_93_tstrb),
        .m_axis_bramio_93_tdata(m_axis_bramio_93_tdata),
        .m_axis_bramio_93_tready(m_axis_bramio_93_tready),
        .m_axis_bramio_94_aclk(m_axis_bramio_94_aclk),
        .m_axis_bramio_94_aresetn(m_axis_bramio_94_aresetn),
        .m_axis_bramio_94_tlast(m_axis_bramio_94_tlast),
        .m_axis_bramio_94_tvalid(m_axis_bramio_94_tvalid),
        .m_axis_bramio_94_tkeep(m_axis_bramio_94_tkeep),
        .m_axis_bramio_94_tstrb(m_axis_bramio_94_tstrb),
        .m_axis_bramio_94_tdata(m_axis_bramio_94_tdata),
        .m_axis_bramio_94_tready(m_axis_bramio_94_tready),
        .m_axis_bramio_95_aclk(m_axis_bramio_95_aclk),
        .m_axis_bramio_95_aresetn(m_axis_bramio_95_aresetn),
        .m_axis_bramio_95_tlast(m_axis_bramio_95_tlast),
        .m_axis_bramio_95_tvalid(m_axis_bramio_95_tvalid),
        .m_axis_bramio_95_tkeep(m_axis_bramio_95_tkeep),
        .m_axis_bramio_95_tstrb(m_axis_bramio_95_tstrb),
        .m_axis_bramio_95_tdata(m_axis_bramio_95_tdata),
        .m_axis_bramio_95_tready(m_axis_bramio_95_tready),
        .m_axis_bramio_96_aclk(m_axis_bramio_96_aclk),
        .m_axis_bramio_96_aresetn(m_axis_bramio_96_aresetn),
        .m_axis_bramio_96_tlast(m_axis_bramio_96_tlast),
        .m_axis_bramio_96_tvalid(m_axis_bramio_96_tvalid),
        .m_axis_bramio_96_tkeep(m_axis_bramio_96_tkeep),
        .m_axis_bramio_96_tstrb(m_axis_bramio_96_tstrb),
        .m_axis_bramio_96_tdata(m_axis_bramio_96_tdata),
        .m_axis_bramio_96_tready(m_axis_bramio_96_tready),
        .m_axis_bramio_97_aclk(m_axis_bramio_97_aclk),
        .m_axis_bramio_97_aresetn(m_axis_bramio_97_aresetn),
        .m_axis_bramio_97_tlast(m_axis_bramio_97_tlast),
        .m_axis_bramio_97_tvalid(m_axis_bramio_97_tvalid),
        .m_axis_bramio_97_tkeep(m_axis_bramio_97_tkeep),
        .m_axis_bramio_97_tstrb(m_axis_bramio_97_tstrb),
        .m_axis_bramio_97_tdata(m_axis_bramio_97_tdata),
        .m_axis_bramio_97_tready(m_axis_bramio_97_tready),
        .m_axis_bramio_98_aclk(m_axis_bramio_98_aclk),
        .m_axis_bramio_98_aresetn(m_axis_bramio_98_aresetn),
        .m_axis_bramio_98_tlast(m_axis_bramio_98_tlast),
        .m_axis_bramio_98_tvalid(m_axis_bramio_98_tvalid),
        .m_axis_bramio_98_tkeep(m_axis_bramio_98_tkeep),
        .m_axis_bramio_98_tstrb(m_axis_bramio_98_tstrb),
        .m_axis_bramio_98_tdata(m_axis_bramio_98_tdata),
        .m_axis_bramio_98_tready(m_axis_bramio_98_tready),
        .m_axis_bramio_99_aclk(m_axis_bramio_99_aclk),
        .m_axis_bramio_99_aresetn(m_axis_bramio_99_aresetn),
        .m_axis_bramio_99_tlast(m_axis_bramio_99_tlast),
        .m_axis_bramio_99_tvalid(m_axis_bramio_99_tvalid),
        .m_axis_bramio_99_tkeep(m_axis_bramio_99_tkeep),
        .m_axis_bramio_99_tstrb(m_axis_bramio_99_tstrb),
        .m_axis_bramio_99_tdata(m_axis_bramio_99_tdata),
        .m_axis_bramio_99_tready(m_axis_bramio_99_tready),
        .m_axis_bramio_100_aclk(m_axis_bramio_100_aclk),
        .m_axis_bramio_100_aresetn(m_axis_bramio_100_aresetn),
        .m_axis_bramio_100_tlast(m_axis_bramio_100_tlast),
        .m_axis_bramio_100_tvalid(m_axis_bramio_100_tvalid),
        .m_axis_bramio_100_tkeep(m_axis_bramio_100_tkeep),
        .m_axis_bramio_100_tstrb(m_axis_bramio_100_tstrb),
        .m_axis_bramio_100_tdata(m_axis_bramio_100_tdata),
        .m_axis_bramio_100_tready(m_axis_bramio_100_tready),
        .m_axis_bramio_101_aclk(m_axis_bramio_101_aclk),
        .m_axis_bramio_101_aresetn(m_axis_bramio_101_aresetn),
        .m_axis_bramio_101_tlast(m_axis_bramio_101_tlast),
        .m_axis_bramio_101_tvalid(m_axis_bramio_101_tvalid),
        .m_axis_bramio_101_tkeep(m_axis_bramio_101_tkeep),
        .m_axis_bramio_101_tstrb(m_axis_bramio_101_tstrb),
        .m_axis_bramio_101_tdata(m_axis_bramio_101_tdata),
        .m_axis_bramio_101_tready(m_axis_bramio_101_tready),
        .m_axis_bramio_102_aclk(m_axis_bramio_102_aclk),
        .m_axis_bramio_102_aresetn(m_axis_bramio_102_aresetn),
        .m_axis_bramio_102_tlast(m_axis_bramio_102_tlast),
        .m_axis_bramio_102_tvalid(m_axis_bramio_102_tvalid),
        .m_axis_bramio_102_tkeep(m_axis_bramio_102_tkeep),
        .m_axis_bramio_102_tstrb(m_axis_bramio_102_tstrb),
        .m_axis_bramio_102_tdata(m_axis_bramio_102_tdata),
        .m_axis_bramio_102_tready(m_axis_bramio_102_tready),
        .m_axis_bramio_103_aclk(m_axis_bramio_103_aclk),
        .m_axis_bramio_103_aresetn(m_axis_bramio_103_aresetn),
        .m_axis_bramio_103_tlast(m_axis_bramio_103_tlast),
        .m_axis_bramio_103_tvalid(m_axis_bramio_103_tvalid),
        .m_axis_bramio_103_tkeep(m_axis_bramio_103_tkeep),
        .m_axis_bramio_103_tstrb(m_axis_bramio_103_tstrb),
        .m_axis_bramio_103_tdata(m_axis_bramio_103_tdata),
        .m_axis_bramio_103_tready(m_axis_bramio_103_tready),
        .m_axis_bramio_104_aclk(m_axis_bramio_104_aclk),
        .m_axis_bramio_104_aresetn(m_axis_bramio_104_aresetn),
        .m_axis_bramio_104_tlast(m_axis_bramio_104_tlast),
        .m_axis_bramio_104_tvalid(m_axis_bramio_104_tvalid),
        .m_axis_bramio_104_tkeep(m_axis_bramio_104_tkeep),
        .m_axis_bramio_104_tstrb(m_axis_bramio_104_tstrb),
        .m_axis_bramio_104_tdata(m_axis_bramio_104_tdata),
        .m_axis_bramio_104_tready(m_axis_bramio_104_tready),
        .m_axis_bramio_105_aclk(m_axis_bramio_105_aclk),
        .m_axis_bramio_105_aresetn(m_axis_bramio_105_aresetn),
        .m_axis_bramio_105_tlast(m_axis_bramio_105_tlast),
        .m_axis_bramio_105_tvalid(m_axis_bramio_105_tvalid),
        .m_axis_bramio_105_tkeep(m_axis_bramio_105_tkeep),
        .m_axis_bramio_105_tstrb(m_axis_bramio_105_tstrb),
        .m_axis_bramio_105_tdata(m_axis_bramio_105_tdata),
        .m_axis_bramio_105_tready(m_axis_bramio_105_tready),
        .m_axis_bramio_106_aclk(m_axis_bramio_106_aclk),
        .m_axis_bramio_106_aresetn(m_axis_bramio_106_aresetn),
        .m_axis_bramio_106_tlast(m_axis_bramio_106_tlast),
        .m_axis_bramio_106_tvalid(m_axis_bramio_106_tvalid),
        .m_axis_bramio_106_tkeep(m_axis_bramio_106_tkeep),
        .m_axis_bramio_106_tstrb(m_axis_bramio_106_tstrb),
        .m_axis_bramio_106_tdata(m_axis_bramio_106_tdata),
        .m_axis_bramio_106_tready(m_axis_bramio_106_tready),
        .m_axis_bramio_107_aclk(m_axis_bramio_107_aclk),
        .m_axis_bramio_107_aresetn(m_axis_bramio_107_aresetn),
        .m_axis_bramio_107_tlast(m_axis_bramio_107_tlast),
        .m_axis_bramio_107_tvalid(m_axis_bramio_107_tvalid),
        .m_axis_bramio_107_tkeep(m_axis_bramio_107_tkeep),
        .m_axis_bramio_107_tstrb(m_axis_bramio_107_tstrb),
        .m_axis_bramio_107_tdata(m_axis_bramio_107_tdata),
        .m_axis_bramio_107_tready(m_axis_bramio_107_tready),
        .m_axis_bramio_108_aclk(m_axis_bramio_108_aclk),
        .m_axis_bramio_108_aresetn(m_axis_bramio_108_aresetn),
        .m_axis_bramio_108_tlast(m_axis_bramio_108_tlast),
        .m_axis_bramio_108_tvalid(m_axis_bramio_108_tvalid),
        .m_axis_bramio_108_tkeep(m_axis_bramio_108_tkeep),
        .m_axis_bramio_108_tstrb(m_axis_bramio_108_tstrb),
        .m_axis_bramio_108_tdata(m_axis_bramio_108_tdata),
        .m_axis_bramio_108_tready(m_axis_bramio_108_tready),
        .m_axis_bramio_109_aclk(m_axis_bramio_109_aclk),
        .m_axis_bramio_109_aresetn(m_axis_bramio_109_aresetn),
        .m_axis_bramio_109_tlast(m_axis_bramio_109_tlast),
        .m_axis_bramio_109_tvalid(m_axis_bramio_109_tvalid),
        .m_axis_bramio_109_tkeep(m_axis_bramio_109_tkeep),
        .m_axis_bramio_109_tstrb(m_axis_bramio_109_tstrb),
        .m_axis_bramio_109_tdata(m_axis_bramio_109_tdata),
        .m_axis_bramio_109_tready(m_axis_bramio_109_tready),
        .m_axis_bramio_110_aclk(m_axis_bramio_110_aclk),
        .m_axis_bramio_110_aresetn(m_axis_bramio_110_aresetn),
        .m_axis_bramio_110_tlast(m_axis_bramio_110_tlast),
        .m_axis_bramio_110_tvalid(m_axis_bramio_110_tvalid),
        .m_axis_bramio_110_tkeep(m_axis_bramio_110_tkeep),
        .m_axis_bramio_110_tstrb(m_axis_bramio_110_tstrb),
        .m_axis_bramio_110_tdata(m_axis_bramio_110_tdata),
        .m_axis_bramio_110_tready(m_axis_bramio_110_tready),
        .m_axis_bramio_111_aclk(m_axis_bramio_111_aclk),
        .m_axis_bramio_111_aresetn(m_axis_bramio_111_aresetn),
        .m_axis_bramio_111_tlast(m_axis_bramio_111_tlast),
        .m_axis_bramio_111_tvalid(m_axis_bramio_111_tvalid),
        .m_axis_bramio_111_tkeep(m_axis_bramio_111_tkeep),
        .m_axis_bramio_111_tstrb(m_axis_bramio_111_tstrb),
        .m_axis_bramio_111_tdata(m_axis_bramio_111_tdata),
        .m_axis_bramio_111_tready(m_axis_bramio_111_tready),
        .m_axis_bramio_112_aclk(m_axis_bramio_112_aclk),
        .m_axis_bramio_112_aresetn(m_axis_bramio_112_aresetn),
        .m_axis_bramio_112_tlast(m_axis_bramio_112_tlast),
        .m_axis_bramio_112_tvalid(m_axis_bramio_112_tvalid),
        .m_axis_bramio_112_tkeep(m_axis_bramio_112_tkeep),
        .m_axis_bramio_112_tstrb(m_axis_bramio_112_tstrb),
        .m_axis_bramio_112_tdata(m_axis_bramio_112_tdata),
        .m_axis_bramio_112_tready(m_axis_bramio_112_tready),
        .m_axis_bramio_113_aclk(m_axis_bramio_113_aclk),
        .m_axis_bramio_113_aresetn(m_axis_bramio_113_aresetn),
        .m_axis_bramio_113_tlast(m_axis_bramio_113_tlast),
        .m_axis_bramio_113_tvalid(m_axis_bramio_113_tvalid),
        .m_axis_bramio_113_tkeep(m_axis_bramio_113_tkeep),
        .m_axis_bramio_113_tstrb(m_axis_bramio_113_tstrb),
        .m_axis_bramio_113_tdata(m_axis_bramio_113_tdata),
        .m_axis_bramio_113_tready(m_axis_bramio_113_tready),
        .m_axis_bramio_114_aclk(m_axis_bramio_114_aclk),
        .m_axis_bramio_114_aresetn(m_axis_bramio_114_aresetn),
        .m_axis_bramio_114_tlast(m_axis_bramio_114_tlast),
        .m_axis_bramio_114_tvalid(m_axis_bramio_114_tvalid),
        .m_axis_bramio_114_tkeep(m_axis_bramio_114_tkeep),
        .m_axis_bramio_114_tstrb(m_axis_bramio_114_tstrb),
        .m_axis_bramio_114_tdata(m_axis_bramio_114_tdata),
        .m_axis_bramio_114_tready(m_axis_bramio_114_tready),
        .m_axis_bramio_115_aclk(m_axis_bramio_115_aclk),
        .m_axis_bramio_115_aresetn(m_axis_bramio_115_aresetn),
        .m_axis_bramio_115_tlast(m_axis_bramio_115_tlast),
        .m_axis_bramio_115_tvalid(m_axis_bramio_115_tvalid),
        .m_axis_bramio_115_tkeep(m_axis_bramio_115_tkeep),
        .m_axis_bramio_115_tstrb(m_axis_bramio_115_tstrb),
        .m_axis_bramio_115_tdata(m_axis_bramio_115_tdata),
        .m_axis_bramio_115_tready(m_axis_bramio_115_tready),
        .m_axis_bramio_116_aclk(m_axis_bramio_116_aclk),
        .m_axis_bramio_116_aresetn(m_axis_bramio_116_aresetn),
        .m_axis_bramio_116_tlast(m_axis_bramio_116_tlast),
        .m_axis_bramio_116_tvalid(m_axis_bramio_116_tvalid),
        .m_axis_bramio_116_tkeep(m_axis_bramio_116_tkeep),
        .m_axis_bramio_116_tstrb(m_axis_bramio_116_tstrb),
        .m_axis_bramio_116_tdata(m_axis_bramio_116_tdata),
        .m_axis_bramio_116_tready(m_axis_bramio_116_tready),
        .m_axis_bramio_117_aclk(m_axis_bramio_117_aclk),
        .m_axis_bramio_117_aresetn(m_axis_bramio_117_aresetn),
        .m_axis_bramio_117_tlast(m_axis_bramio_117_tlast),
        .m_axis_bramio_117_tvalid(m_axis_bramio_117_tvalid),
        .m_axis_bramio_117_tkeep(m_axis_bramio_117_tkeep),
        .m_axis_bramio_117_tstrb(m_axis_bramio_117_tstrb),
        .m_axis_bramio_117_tdata(m_axis_bramio_117_tdata),
        .m_axis_bramio_117_tready(m_axis_bramio_117_tready),
        .m_axis_bramio_118_aclk(m_axis_bramio_118_aclk),
        .m_axis_bramio_118_aresetn(m_axis_bramio_118_aresetn),
        .m_axis_bramio_118_tlast(m_axis_bramio_118_tlast),
        .m_axis_bramio_118_tvalid(m_axis_bramio_118_tvalid),
        .m_axis_bramio_118_tkeep(m_axis_bramio_118_tkeep),
        .m_axis_bramio_118_tstrb(m_axis_bramio_118_tstrb),
        .m_axis_bramio_118_tdata(m_axis_bramio_118_tdata),
        .m_axis_bramio_118_tready(m_axis_bramio_118_tready),
        .m_axis_bramio_119_aclk(m_axis_bramio_119_aclk),
        .m_axis_bramio_119_aresetn(m_axis_bramio_119_aresetn),
        .m_axis_bramio_119_tlast(m_axis_bramio_119_tlast),
        .m_axis_bramio_119_tvalid(m_axis_bramio_119_tvalid),
        .m_axis_bramio_119_tkeep(m_axis_bramio_119_tkeep),
        .m_axis_bramio_119_tstrb(m_axis_bramio_119_tstrb),
        .m_axis_bramio_119_tdata(m_axis_bramio_119_tdata),
        .m_axis_bramio_119_tready(m_axis_bramio_119_tready),
        .m_axis_bramio_120_aclk(m_axis_bramio_120_aclk),
        .m_axis_bramio_120_aresetn(m_axis_bramio_120_aresetn),
        .m_axis_bramio_120_tlast(m_axis_bramio_120_tlast),
        .m_axis_bramio_120_tvalid(m_axis_bramio_120_tvalid),
        .m_axis_bramio_120_tkeep(m_axis_bramio_120_tkeep),
        .m_axis_bramio_120_tstrb(m_axis_bramio_120_tstrb),
        .m_axis_bramio_120_tdata(m_axis_bramio_120_tdata),
        .m_axis_bramio_120_tready(m_axis_bramio_120_tready),
        .m_axis_bramio_121_aclk(m_axis_bramio_121_aclk),
        .m_axis_bramio_121_aresetn(m_axis_bramio_121_aresetn),
        .m_axis_bramio_121_tlast(m_axis_bramio_121_tlast),
        .m_axis_bramio_121_tvalid(m_axis_bramio_121_tvalid),
        .m_axis_bramio_121_tkeep(m_axis_bramio_121_tkeep),
        .m_axis_bramio_121_tstrb(m_axis_bramio_121_tstrb),
        .m_axis_bramio_121_tdata(m_axis_bramio_121_tdata),
        .m_axis_bramio_121_tready(m_axis_bramio_121_tready),
        .m_axis_bramio_122_aclk(m_axis_bramio_122_aclk),
        .m_axis_bramio_122_aresetn(m_axis_bramio_122_aresetn),
        .m_axis_bramio_122_tlast(m_axis_bramio_122_tlast),
        .m_axis_bramio_122_tvalid(m_axis_bramio_122_tvalid),
        .m_axis_bramio_122_tkeep(m_axis_bramio_122_tkeep),
        .m_axis_bramio_122_tstrb(m_axis_bramio_122_tstrb),
        .m_axis_bramio_122_tdata(m_axis_bramio_122_tdata),
        .m_axis_bramio_122_tready(m_axis_bramio_122_tready),
        .m_axis_bramio_123_aclk(m_axis_bramio_123_aclk),
        .m_axis_bramio_123_aresetn(m_axis_bramio_123_aresetn),
        .m_axis_bramio_123_tlast(m_axis_bramio_123_tlast),
        .m_axis_bramio_123_tvalid(m_axis_bramio_123_tvalid),
        .m_axis_bramio_123_tkeep(m_axis_bramio_123_tkeep),
        .m_axis_bramio_123_tstrb(m_axis_bramio_123_tstrb),
        .m_axis_bramio_123_tdata(m_axis_bramio_123_tdata),
        .m_axis_bramio_123_tready(m_axis_bramio_123_tready),
        .m_axis_bramio_124_aclk(m_axis_bramio_124_aclk),
        .m_axis_bramio_124_aresetn(m_axis_bramio_124_aresetn),
        .m_axis_bramio_124_tlast(m_axis_bramio_124_tlast),
        .m_axis_bramio_124_tvalid(m_axis_bramio_124_tvalid),
        .m_axis_bramio_124_tkeep(m_axis_bramio_124_tkeep),
        .m_axis_bramio_124_tstrb(m_axis_bramio_124_tstrb),
        .m_axis_bramio_124_tdata(m_axis_bramio_124_tdata),
        .m_axis_bramio_124_tready(m_axis_bramio_124_tready),
        .m_axis_bramio_125_aclk(m_axis_bramio_125_aclk),
        .m_axis_bramio_125_aresetn(m_axis_bramio_125_aresetn),
        .m_axis_bramio_125_tlast(m_axis_bramio_125_tlast),
        .m_axis_bramio_125_tvalid(m_axis_bramio_125_tvalid),
        .m_axis_bramio_125_tkeep(m_axis_bramio_125_tkeep),
        .m_axis_bramio_125_tstrb(m_axis_bramio_125_tstrb),
        .m_axis_bramio_125_tdata(m_axis_bramio_125_tdata),
        .m_axis_bramio_125_tready(m_axis_bramio_125_tready),
        .m_axis_bramio_126_aclk(m_axis_bramio_126_aclk),
        .m_axis_bramio_126_aresetn(m_axis_bramio_126_aresetn),
        .m_axis_bramio_126_tlast(m_axis_bramio_126_tlast),
        .m_axis_bramio_126_tvalid(m_axis_bramio_126_tvalid),
        .m_axis_bramio_126_tkeep(m_axis_bramio_126_tkeep),
        .m_axis_bramio_126_tstrb(m_axis_bramio_126_tstrb),
        .m_axis_bramio_126_tdata(m_axis_bramio_126_tdata),
        .m_axis_bramio_126_tready(m_axis_bramio_126_tready),
        .m_axis_bramio_127_aclk(m_axis_bramio_127_aclk),
        .m_axis_bramio_127_aresetn(m_axis_bramio_127_aresetn),
        .m_axis_bramio_127_tlast(m_axis_bramio_127_tlast),
        .m_axis_bramio_127_tvalid(m_axis_bramio_127_tvalid),
        .m_axis_bramio_127_tkeep(m_axis_bramio_127_tkeep),
        .m_axis_bramio_127_tstrb(m_axis_bramio_127_tstrb),
        .m_axis_bramio_127_tdata(m_axis_bramio_127_tdata),
        .m_axis_bramio_127_tready(m_axis_bramio_127_tready)
    );
    
    out_bram_args #(
        .C_QUEUE_DEPTH(C_QUEUE_DEPTH),
        .C_NUM_OUTPUT_BRAMs(C_NUM_OUTPUT_BRAMs),
        .M_AXIS_BRAM_0_WIDTH(M_AXIS_BRAM_0_WIDTH),
        .M_AXIS_BRAM_1_WIDTH(M_AXIS_BRAM_1_WIDTH),
        .M_AXIS_BRAM_2_WIDTH(M_AXIS_BRAM_2_WIDTH),
        .M_AXIS_BRAM_3_WIDTH(M_AXIS_BRAM_3_WIDTH),
        .M_AXIS_BRAM_4_WIDTH(M_AXIS_BRAM_4_WIDTH),
        .M_AXIS_BRAM_5_WIDTH(M_AXIS_BRAM_5_WIDTH),
        .M_AXIS_BRAM_6_WIDTH(M_AXIS_BRAM_6_WIDTH),
        .M_AXIS_BRAM_7_WIDTH(M_AXIS_BRAM_7_WIDTH),
        .M_AXIS_BRAM_8_WIDTH(M_AXIS_BRAM_8_WIDTH),
        .M_AXIS_BRAM_9_WIDTH(M_AXIS_BRAM_9_WIDTH),
        .M_AXIS_BRAM_10_WIDTH(M_AXIS_BRAM_10_WIDTH),
        .M_AXIS_BRAM_11_WIDTH(M_AXIS_BRAM_11_WIDTH),
        .M_AXIS_BRAM_12_WIDTH(M_AXIS_BRAM_12_WIDTH),
        .M_AXIS_BRAM_13_WIDTH(M_AXIS_BRAM_13_WIDTH),
        .M_AXIS_BRAM_14_WIDTH(M_AXIS_BRAM_14_WIDTH),
        .M_AXIS_BRAM_15_WIDTH(M_AXIS_BRAM_15_WIDTH),
        .M_AXIS_BRAM_16_WIDTH(M_AXIS_BRAM_16_WIDTH),
        .M_AXIS_BRAM_17_WIDTH(M_AXIS_BRAM_17_WIDTH),
        .M_AXIS_BRAM_18_WIDTH(M_AXIS_BRAM_18_WIDTH),
        .M_AXIS_BRAM_19_WIDTH(M_AXIS_BRAM_19_WIDTH),
        .M_AXIS_BRAM_20_WIDTH(M_AXIS_BRAM_20_WIDTH),
        .M_AXIS_BRAM_21_WIDTH(M_AXIS_BRAM_21_WIDTH),
        .M_AXIS_BRAM_22_WIDTH(M_AXIS_BRAM_22_WIDTH),
        .M_AXIS_BRAM_23_WIDTH(M_AXIS_BRAM_23_WIDTH),
        .M_AXIS_BRAM_24_WIDTH(M_AXIS_BRAM_24_WIDTH),
        .M_AXIS_BRAM_25_WIDTH(M_AXIS_BRAM_25_WIDTH),
        .M_AXIS_BRAM_26_WIDTH(M_AXIS_BRAM_26_WIDTH),
        .M_AXIS_BRAM_27_WIDTH(M_AXIS_BRAM_27_WIDTH),
        .M_AXIS_BRAM_28_WIDTH(M_AXIS_BRAM_28_WIDTH),
        .M_AXIS_BRAM_29_WIDTH(M_AXIS_BRAM_29_WIDTH),
        .M_AXIS_BRAM_30_WIDTH(M_AXIS_BRAM_30_WIDTH),
        .M_AXIS_BRAM_31_WIDTH(M_AXIS_BRAM_31_WIDTH),
        .M_AXIS_BRAM_32_WIDTH(M_AXIS_BRAM_32_WIDTH),
        .M_AXIS_BRAM_33_WIDTH(M_AXIS_BRAM_33_WIDTH),
        .M_AXIS_BRAM_34_WIDTH(M_AXIS_BRAM_34_WIDTH),
        .M_AXIS_BRAM_35_WIDTH(M_AXIS_BRAM_35_WIDTH),
        .M_AXIS_BRAM_36_WIDTH(M_AXIS_BRAM_36_WIDTH),
        .M_AXIS_BRAM_37_WIDTH(M_AXIS_BRAM_37_WIDTH),
        .M_AXIS_BRAM_38_WIDTH(M_AXIS_BRAM_38_WIDTH),
        .M_AXIS_BRAM_39_WIDTH(M_AXIS_BRAM_39_WIDTH),
        .M_AXIS_BRAM_40_WIDTH(M_AXIS_BRAM_40_WIDTH),
        .M_AXIS_BRAM_41_WIDTH(M_AXIS_BRAM_41_WIDTH),
        .M_AXIS_BRAM_42_WIDTH(M_AXIS_BRAM_42_WIDTH),
        .M_AXIS_BRAM_43_WIDTH(M_AXIS_BRAM_43_WIDTH),
        .M_AXIS_BRAM_44_WIDTH(M_AXIS_BRAM_44_WIDTH),
        .M_AXIS_BRAM_45_WIDTH(M_AXIS_BRAM_45_WIDTH),
        .M_AXIS_BRAM_46_WIDTH(M_AXIS_BRAM_46_WIDTH),
        .M_AXIS_BRAM_47_WIDTH(M_AXIS_BRAM_47_WIDTH),
        .M_AXIS_BRAM_48_WIDTH(M_AXIS_BRAM_48_WIDTH),
        .M_AXIS_BRAM_49_WIDTH(M_AXIS_BRAM_49_WIDTH),
        .M_AXIS_BRAM_50_WIDTH(M_AXIS_BRAM_50_WIDTH),
        .M_AXIS_BRAM_51_WIDTH(M_AXIS_BRAM_51_WIDTH),
        .M_AXIS_BRAM_52_WIDTH(M_AXIS_BRAM_52_WIDTH),
        .M_AXIS_BRAM_53_WIDTH(M_AXIS_BRAM_53_WIDTH),
        .M_AXIS_BRAM_54_WIDTH(M_AXIS_BRAM_54_WIDTH),
        .M_AXIS_BRAM_55_WIDTH(M_AXIS_BRAM_55_WIDTH),
        .M_AXIS_BRAM_56_WIDTH(M_AXIS_BRAM_56_WIDTH),
        .M_AXIS_BRAM_57_WIDTH(M_AXIS_BRAM_57_WIDTH),
        .M_AXIS_BRAM_58_WIDTH(M_AXIS_BRAM_58_WIDTH),
        .M_AXIS_BRAM_59_WIDTH(M_AXIS_BRAM_59_WIDTH),
        .M_AXIS_BRAM_60_WIDTH(M_AXIS_BRAM_60_WIDTH),
        .M_AXIS_BRAM_61_WIDTH(M_AXIS_BRAM_61_WIDTH),
        .M_AXIS_BRAM_62_WIDTH(M_AXIS_BRAM_62_WIDTH),
        .M_AXIS_BRAM_63_WIDTH(M_AXIS_BRAM_63_WIDTH),
        .M_AXIS_BRAM_64_WIDTH(M_AXIS_BRAM_64_WIDTH),
        .M_AXIS_BRAM_65_WIDTH(M_AXIS_BRAM_65_WIDTH),
        .M_AXIS_BRAM_66_WIDTH(M_AXIS_BRAM_66_WIDTH),
        .M_AXIS_BRAM_67_WIDTH(M_AXIS_BRAM_67_WIDTH),
        .M_AXIS_BRAM_68_WIDTH(M_AXIS_BRAM_68_WIDTH),
        .M_AXIS_BRAM_69_WIDTH(M_AXIS_BRAM_69_WIDTH),
        .M_AXIS_BRAM_70_WIDTH(M_AXIS_BRAM_70_WIDTH),
        .M_AXIS_BRAM_71_WIDTH(M_AXIS_BRAM_71_WIDTH),
        .M_AXIS_BRAM_72_WIDTH(M_AXIS_BRAM_72_WIDTH),
        .M_AXIS_BRAM_73_WIDTH(M_AXIS_BRAM_73_WIDTH),
        .M_AXIS_BRAM_74_WIDTH(M_AXIS_BRAM_74_WIDTH),
        .M_AXIS_BRAM_75_WIDTH(M_AXIS_BRAM_75_WIDTH),
        .M_AXIS_BRAM_76_WIDTH(M_AXIS_BRAM_76_WIDTH),
        .M_AXIS_BRAM_77_WIDTH(M_AXIS_BRAM_77_WIDTH),
        .M_AXIS_BRAM_78_WIDTH(M_AXIS_BRAM_78_WIDTH),
        .M_AXIS_BRAM_79_WIDTH(M_AXIS_BRAM_79_WIDTH),
        .M_AXIS_BRAM_80_WIDTH(M_AXIS_BRAM_80_WIDTH),
        .M_AXIS_BRAM_81_WIDTH(M_AXIS_BRAM_81_WIDTH),
        .M_AXIS_BRAM_82_WIDTH(M_AXIS_BRAM_82_WIDTH),
        .M_AXIS_BRAM_83_WIDTH(M_AXIS_BRAM_83_WIDTH),
        .M_AXIS_BRAM_84_WIDTH(M_AXIS_BRAM_84_WIDTH),
        .M_AXIS_BRAM_85_WIDTH(M_AXIS_BRAM_85_WIDTH),
        .M_AXIS_BRAM_86_WIDTH(M_AXIS_BRAM_86_WIDTH),
        .M_AXIS_BRAM_87_WIDTH(M_AXIS_BRAM_87_WIDTH),
        .M_AXIS_BRAM_88_WIDTH(M_AXIS_BRAM_88_WIDTH),
        .M_AXIS_BRAM_89_WIDTH(M_AXIS_BRAM_89_WIDTH),
        .M_AXIS_BRAM_90_WIDTH(M_AXIS_BRAM_90_WIDTH),
        .M_AXIS_BRAM_91_WIDTH(M_AXIS_BRAM_91_WIDTH),
        .M_AXIS_BRAM_92_WIDTH(M_AXIS_BRAM_92_WIDTH),
        .M_AXIS_BRAM_93_WIDTH(M_AXIS_BRAM_93_WIDTH),
        .M_AXIS_BRAM_94_WIDTH(M_AXIS_BRAM_94_WIDTH),
        .M_AXIS_BRAM_95_WIDTH(M_AXIS_BRAM_95_WIDTH),
        .M_AXIS_BRAM_96_WIDTH(M_AXIS_BRAM_96_WIDTH),
        .M_AXIS_BRAM_97_WIDTH(M_AXIS_BRAM_97_WIDTH),
        .M_AXIS_BRAM_98_WIDTH(M_AXIS_BRAM_98_WIDTH),
        .M_AXIS_BRAM_99_WIDTH(M_AXIS_BRAM_99_WIDTH),
        .M_AXIS_BRAM_100_WIDTH(M_AXIS_BRAM_100_WIDTH),
        .M_AXIS_BRAM_101_WIDTH(M_AXIS_BRAM_101_WIDTH),
        .M_AXIS_BRAM_102_WIDTH(M_AXIS_BRAM_102_WIDTH),
        .M_AXIS_BRAM_103_WIDTH(M_AXIS_BRAM_103_WIDTH),
        .M_AXIS_BRAM_104_WIDTH(M_AXIS_BRAM_104_WIDTH),
        .M_AXIS_BRAM_105_WIDTH(M_AXIS_BRAM_105_WIDTH),
        .M_AXIS_BRAM_106_WIDTH(M_AXIS_BRAM_106_WIDTH),
        .M_AXIS_BRAM_107_WIDTH(M_AXIS_BRAM_107_WIDTH),
        .M_AXIS_BRAM_108_WIDTH(M_AXIS_BRAM_108_WIDTH),
        .M_AXIS_BRAM_109_WIDTH(M_AXIS_BRAM_109_WIDTH),
        .M_AXIS_BRAM_110_WIDTH(M_AXIS_BRAM_110_WIDTH),
        .M_AXIS_BRAM_111_WIDTH(M_AXIS_BRAM_111_WIDTH),
        .M_AXIS_BRAM_112_WIDTH(M_AXIS_BRAM_112_WIDTH),
        .M_AXIS_BRAM_113_WIDTH(M_AXIS_BRAM_113_WIDTH),
        .M_AXIS_BRAM_114_WIDTH(M_AXIS_BRAM_114_WIDTH),
        .M_AXIS_BRAM_115_WIDTH(M_AXIS_BRAM_115_WIDTH),
        .M_AXIS_BRAM_116_WIDTH(M_AXIS_BRAM_116_WIDTH),
        .M_AXIS_BRAM_117_WIDTH(M_AXIS_BRAM_117_WIDTH),
        .M_AXIS_BRAM_118_WIDTH(M_AXIS_BRAM_118_WIDTH),
        .M_AXIS_BRAM_119_WIDTH(M_AXIS_BRAM_119_WIDTH),
        .M_AXIS_BRAM_120_WIDTH(M_AXIS_BRAM_120_WIDTH),
        .M_AXIS_BRAM_121_WIDTH(M_AXIS_BRAM_121_WIDTH),
        .M_AXIS_BRAM_122_WIDTH(M_AXIS_BRAM_122_WIDTH),
        .M_AXIS_BRAM_123_WIDTH(M_AXIS_BRAM_123_WIDTH),
        .M_AXIS_BRAM_124_WIDTH(M_AXIS_BRAM_124_WIDTH),
        .M_AXIS_BRAM_125_WIDTH(M_AXIS_BRAM_125_WIDTH),
        .M_AXIS_BRAM_126_WIDTH(M_AXIS_BRAM_126_WIDTH),
        .M_AXIS_BRAM_127_WIDTH(M_AXIS_BRAM_127_WIDTH),
        .M_AXIS_BRAM_0_DEPTH(M_AXIS_BRAM_0_DEPTH),
        .M_AXIS_BRAM_1_DEPTH(M_AXIS_BRAM_1_DEPTH),
        .M_AXIS_BRAM_2_DEPTH(M_AXIS_BRAM_2_DEPTH),
        .M_AXIS_BRAM_3_DEPTH(M_AXIS_BRAM_3_DEPTH),
        .M_AXIS_BRAM_4_DEPTH(M_AXIS_BRAM_4_DEPTH),
        .M_AXIS_BRAM_5_DEPTH(M_AXIS_BRAM_5_DEPTH),
        .M_AXIS_BRAM_6_DEPTH(M_AXIS_BRAM_6_DEPTH),
        .M_AXIS_BRAM_7_DEPTH(M_AXIS_BRAM_7_DEPTH),
        .M_AXIS_BRAM_8_DEPTH(M_AXIS_BRAM_8_DEPTH),
        .M_AXIS_BRAM_9_DEPTH(M_AXIS_BRAM_9_DEPTH),
        .M_AXIS_BRAM_10_DEPTH(M_AXIS_BRAM_10_DEPTH),
        .M_AXIS_BRAM_11_DEPTH(M_AXIS_BRAM_11_DEPTH),
        .M_AXIS_BRAM_12_DEPTH(M_AXIS_BRAM_12_DEPTH),
        .M_AXIS_BRAM_13_DEPTH(M_AXIS_BRAM_13_DEPTH),
        .M_AXIS_BRAM_14_DEPTH(M_AXIS_BRAM_14_DEPTH),
        .M_AXIS_BRAM_15_DEPTH(M_AXIS_BRAM_15_DEPTH),
        .M_AXIS_BRAM_16_DEPTH(M_AXIS_BRAM_16_DEPTH),
        .M_AXIS_BRAM_17_DEPTH(M_AXIS_BRAM_17_DEPTH),
        .M_AXIS_BRAM_18_DEPTH(M_AXIS_BRAM_18_DEPTH),
        .M_AXIS_BRAM_19_DEPTH(M_AXIS_BRAM_19_DEPTH),
        .M_AXIS_BRAM_20_DEPTH(M_AXIS_BRAM_20_DEPTH),
        .M_AXIS_BRAM_21_DEPTH(M_AXIS_BRAM_21_DEPTH),
        .M_AXIS_BRAM_22_DEPTH(M_AXIS_BRAM_22_DEPTH),
        .M_AXIS_BRAM_23_DEPTH(M_AXIS_BRAM_23_DEPTH),
        .M_AXIS_BRAM_24_DEPTH(M_AXIS_BRAM_24_DEPTH),
        .M_AXIS_BRAM_25_DEPTH(M_AXIS_BRAM_25_DEPTH),
        .M_AXIS_BRAM_26_DEPTH(M_AXIS_BRAM_26_DEPTH),
        .M_AXIS_BRAM_27_DEPTH(M_AXIS_BRAM_27_DEPTH),
        .M_AXIS_BRAM_28_DEPTH(M_AXIS_BRAM_28_DEPTH),
        .M_AXIS_BRAM_29_DEPTH(M_AXIS_BRAM_29_DEPTH),
        .M_AXIS_BRAM_30_DEPTH(M_AXIS_BRAM_30_DEPTH),
        .M_AXIS_BRAM_31_DEPTH(M_AXIS_BRAM_31_DEPTH),
        .M_AXIS_BRAM_32_DEPTH(M_AXIS_BRAM_32_DEPTH),
        .M_AXIS_BRAM_33_DEPTH(M_AXIS_BRAM_33_DEPTH),
        .M_AXIS_BRAM_34_DEPTH(M_AXIS_BRAM_34_DEPTH),
        .M_AXIS_BRAM_35_DEPTH(M_AXIS_BRAM_35_DEPTH),
        .M_AXIS_BRAM_36_DEPTH(M_AXIS_BRAM_36_DEPTH),
        .M_AXIS_BRAM_37_DEPTH(M_AXIS_BRAM_37_DEPTH),
        .M_AXIS_BRAM_38_DEPTH(M_AXIS_BRAM_38_DEPTH),
        .M_AXIS_BRAM_39_DEPTH(M_AXIS_BRAM_39_DEPTH),
        .M_AXIS_BRAM_40_DEPTH(M_AXIS_BRAM_40_DEPTH),
        .M_AXIS_BRAM_41_DEPTH(M_AXIS_BRAM_41_DEPTH),
        .M_AXIS_BRAM_42_DEPTH(M_AXIS_BRAM_42_DEPTH),
        .M_AXIS_BRAM_43_DEPTH(M_AXIS_BRAM_43_DEPTH),
        .M_AXIS_BRAM_44_DEPTH(M_AXIS_BRAM_44_DEPTH),
        .M_AXIS_BRAM_45_DEPTH(M_AXIS_BRAM_45_DEPTH),
        .M_AXIS_BRAM_46_DEPTH(M_AXIS_BRAM_46_DEPTH),
        .M_AXIS_BRAM_47_DEPTH(M_AXIS_BRAM_47_DEPTH),
        .M_AXIS_BRAM_48_DEPTH(M_AXIS_BRAM_48_DEPTH),
        .M_AXIS_BRAM_49_DEPTH(M_AXIS_BRAM_49_DEPTH),
        .M_AXIS_BRAM_50_DEPTH(M_AXIS_BRAM_50_DEPTH),
        .M_AXIS_BRAM_51_DEPTH(M_AXIS_BRAM_51_DEPTH),
        .M_AXIS_BRAM_52_DEPTH(M_AXIS_BRAM_52_DEPTH),
        .M_AXIS_BRAM_53_DEPTH(M_AXIS_BRAM_53_DEPTH),
        .M_AXIS_BRAM_54_DEPTH(M_AXIS_BRAM_54_DEPTH),
        .M_AXIS_BRAM_55_DEPTH(M_AXIS_BRAM_55_DEPTH),
        .M_AXIS_BRAM_56_DEPTH(M_AXIS_BRAM_56_DEPTH),
        .M_AXIS_BRAM_57_DEPTH(M_AXIS_BRAM_57_DEPTH),
        .M_AXIS_BRAM_58_DEPTH(M_AXIS_BRAM_58_DEPTH),
        .M_AXIS_BRAM_59_DEPTH(M_AXIS_BRAM_59_DEPTH),
        .M_AXIS_BRAM_60_DEPTH(M_AXIS_BRAM_60_DEPTH),
        .M_AXIS_BRAM_61_DEPTH(M_AXIS_BRAM_61_DEPTH),
        .M_AXIS_BRAM_62_DEPTH(M_AXIS_BRAM_62_DEPTH),
        .M_AXIS_BRAM_63_DEPTH(M_AXIS_BRAM_63_DEPTH),
        .M_AXIS_BRAM_64_DEPTH(M_AXIS_BRAM_64_DEPTH),
        .M_AXIS_BRAM_65_DEPTH(M_AXIS_BRAM_65_DEPTH),
        .M_AXIS_BRAM_66_DEPTH(M_AXIS_BRAM_66_DEPTH),
        .M_AXIS_BRAM_67_DEPTH(M_AXIS_BRAM_67_DEPTH),
        .M_AXIS_BRAM_68_DEPTH(M_AXIS_BRAM_68_DEPTH),
        .M_AXIS_BRAM_69_DEPTH(M_AXIS_BRAM_69_DEPTH),
        .M_AXIS_BRAM_70_DEPTH(M_AXIS_BRAM_70_DEPTH),
        .M_AXIS_BRAM_71_DEPTH(M_AXIS_BRAM_71_DEPTH),
        .M_AXIS_BRAM_72_DEPTH(M_AXIS_BRAM_72_DEPTH),
        .M_AXIS_BRAM_73_DEPTH(M_AXIS_BRAM_73_DEPTH),
        .M_AXIS_BRAM_74_DEPTH(M_AXIS_BRAM_74_DEPTH),
        .M_AXIS_BRAM_75_DEPTH(M_AXIS_BRAM_75_DEPTH),
        .M_AXIS_BRAM_76_DEPTH(M_AXIS_BRAM_76_DEPTH),
        .M_AXIS_BRAM_77_DEPTH(M_AXIS_BRAM_77_DEPTH),
        .M_AXIS_BRAM_78_DEPTH(M_AXIS_BRAM_78_DEPTH),
        .M_AXIS_BRAM_79_DEPTH(M_AXIS_BRAM_79_DEPTH),
        .M_AXIS_BRAM_80_DEPTH(M_AXIS_BRAM_80_DEPTH),
        .M_AXIS_BRAM_81_DEPTH(M_AXIS_BRAM_81_DEPTH),
        .M_AXIS_BRAM_82_DEPTH(M_AXIS_BRAM_82_DEPTH),
        .M_AXIS_BRAM_83_DEPTH(M_AXIS_BRAM_83_DEPTH),
        .M_AXIS_BRAM_84_DEPTH(M_AXIS_BRAM_84_DEPTH),
        .M_AXIS_BRAM_85_DEPTH(M_AXIS_BRAM_85_DEPTH),
        .M_AXIS_BRAM_86_DEPTH(M_AXIS_BRAM_86_DEPTH),
        .M_AXIS_BRAM_87_DEPTH(M_AXIS_BRAM_87_DEPTH),
        .M_AXIS_BRAM_88_DEPTH(M_AXIS_BRAM_88_DEPTH),
        .M_AXIS_BRAM_89_DEPTH(M_AXIS_BRAM_89_DEPTH),
        .M_AXIS_BRAM_90_DEPTH(M_AXIS_BRAM_90_DEPTH),
        .M_AXIS_BRAM_91_DEPTH(M_AXIS_BRAM_91_DEPTH),
        .M_AXIS_BRAM_92_DEPTH(M_AXIS_BRAM_92_DEPTH),
        .M_AXIS_BRAM_93_DEPTH(M_AXIS_BRAM_93_DEPTH),
        .M_AXIS_BRAM_94_DEPTH(M_AXIS_BRAM_94_DEPTH),
        .M_AXIS_BRAM_95_DEPTH(M_AXIS_BRAM_95_DEPTH),
        .M_AXIS_BRAM_96_DEPTH(M_AXIS_BRAM_96_DEPTH),
        .M_AXIS_BRAM_97_DEPTH(M_AXIS_BRAM_97_DEPTH),
        .M_AXIS_BRAM_98_DEPTH(M_AXIS_BRAM_98_DEPTH),
        .M_AXIS_BRAM_99_DEPTH(M_AXIS_BRAM_99_DEPTH),
        .M_AXIS_BRAM_100_DEPTH(M_AXIS_BRAM_100_DEPTH),
        .M_AXIS_BRAM_101_DEPTH(M_AXIS_BRAM_101_DEPTH),
        .M_AXIS_BRAM_102_DEPTH(M_AXIS_BRAM_102_DEPTH),
        .M_AXIS_BRAM_103_DEPTH(M_AXIS_BRAM_103_DEPTH),
        .M_AXIS_BRAM_104_DEPTH(M_AXIS_BRAM_104_DEPTH),
        .M_AXIS_BRAM_105_DEPTH(M_AXIS_BRAM_105_DEPTH),
        .M_AXIS_BRAM_106_DEPTH(M_AXIS_BRAM_106_DEPTH),
        .M_AXIS_BRAM_107_DEPTH(M_AXIS_BRAM_107_DEPTH),
        .M_AXIS_BRAM_108_DEPTH(M_AXIS_BRAM_108_DEPTH),
        .M_AXIS_BRAM_109_DEPTH(M_AXIS_BRAM_109_DEPTH),
        .M_AXIS_BRAM_110_DEPTH(M_AXIS_BRAM_110_DEPTH),
        .M_AXIS_BRAM_111_DEPTH(M_AXIS_BRAM_111_DEPTH),
        .M_AXIS_BRAM_112_DEPTH(M_AXIS_BRAM_112_DEPTH),
        .M_AXIS_BRAM_113_DEPTH(M_AXIS_BRAM_113_DEPTH),
        .M_AXIS_BRAM_114_DEPTH(M_AXIS_BRAM_114_DEPTH),
        .M_AXIS_BRAM_115_DEPTH(M_AXIS_BRAM_115_DEPTH),
        .M_AXIS_BRAM_116_DEPTH(M_AXIS_BRAM_116_DEPTH),
        .M_AXIS_BRAM_117_DEPTH(M_AXIS_BRAM_117_DEPTH),
        .M_AXIS_BRAM_118_DEPTH(M_AXIS_BRAM_118_DEPTH),
        .M_AXIS_BRAM_119_DEPTH(M_AXIS_BRAM_119_DEPTH),
        .M_AXIS_BRAM_120_DEPTH(M_AXIS_BRAM_120_DEPTH),
        .M_AXIS_BRAM_121_DEPTH(M_AXIS_BRAM_121_DEPTH),
        .M_AXIS_BRAM_122_DEPTH(M_AXIS_BRAM_122_DEPTH),
        .M_AXIS_BRAM_123_DEPTH(M_AXIS_BRAM_123_DEPTH),
        .M_AXIS_BRAM_124_DEPTH(M_AXIS_BRAM_124_DEPTH),
        .M_AXIS_BRAM_125_DEPTH(M_AXIS_BRAM_125_DEPTH),
        .M_AXIS_BRAM_126_DEPTH(M_AXIS_BRAM_126_DEPTH),
        .M_AXIS_BRAM_127_DEPTH(M_AXIS_BRAM_127_DEPTH),
        .M_AXIS_BRAM_0_DMWIDTH(M_AXIS_BRAM_0_DMWIDTH),
        .M_AXIS_BRAM_1_DMWIDTH(M_AXIS_BRAM_1_DMWIDTH),
        .M_AXIS_BRAM_2_DMWIDTH(M_AXIS_BRAM_2_DMWIDTH),
        .M_AXIS_BRAM_3_DMWIDTH(M_AXIS_BRAM_3_DMWIDTH),
        .M_AXIS_BRAM_4_DMWIDTH(M_AXIS_BRAM_4_DMWIDTH),
        .M_AXIS_BRAM_5_DMWIDTH(M_AXIS_BRAM_5_DMWIDTH),
        .M_AXIS_BRAM_6_DMWIDTH(M_AXIS_BRAM_6_DMWIDTH),
        .M_AXIS_BRAM_7_DMWIDTH(M_AXIS_BRAM_7_DMWIDTH),
        .M_AXIS_BRAM_8_DMWIDTH(M_AXIS_BRAM_8_DMWIDTH),
        .M_AXIS_BRAM_9_DMWIDTH(M_AXIS_BRAM_9_DMWIDTH),
        .M_AXIS_BRAM_10_DMWIDTH(M_AXIS_BRAM_10_DMWIDTH),
        .M_AXIS_BRAM_11_DMWIDTH(M_AXIS_BRAM_11_DMWIDTH),
        .M_AXIS_BRAM_12_DMWIDTH(M_AXIS_BRAM_12_DMWIDTH),
        .M_AXIS_BRAM_13_DMWIDTH(M_AXIS_BRAM_13_DMWIDTH),
        .M_AXIS_BRAM_14_DMWIDTH(M_AXIS_BRAM_14_DMWIDTH),
        .M_AXIS_BRAM_15_DMWIDTH(M_AXIS_BRAM_15_DMWIDTH),
        .M_AXIS_BRAM_16_DMWIDTH(M_AXIS_BRAM_16_DMWIDTH),
        .M_AXIS_BRAM_17_DMWIDTH(M_AXIS_BRAM_17_DMWIDTH),
        .M_AXIS_BRAM_18_DMWIDTH(M_AXIS_BRAM_18_DMWIDTH),
        .M_AXIS_BRAM_19_DMWIDTH(M_AXIS_BRAM_19_DMWIDTH),
        .M_AXIS_BRAM_20_DMWIDTH(M_AXIS_BRAM_20_DMWIDTH),
        .M_AXIS_BRAM_21_DMWIDTH(M_AXIS_BRAM_21_DMWIDTH),
        .M_AXIS_BRAM_22_DMWIDTH(M_AXIS_BRAM_22_DMWIDTH),
        .M_AXIS_BRAM_23_DMWIDTH(M_AXIS_BRAM_23_DMWIDTH),
        .M_AXIS_BRAM_24_DMWIDTH(M_AXIS_BRAM_24_DMWIDTH),
        .M_AXIS_BRAM_25_DMWIDTH(M_AXIS_BRAM_25_DMWIDTH),
        .M_AXIS_BRAM_26_DMWIDTH(M_AXIS_BRAM_26_DMWIDTH),
        .M_AXIS_BRAM_27_DMWIDTH(M_AXIS_BRAM_27_DMWIDTH),
        .M_AXIS_BRAM_28_DMWIDTH(M_AXIS_BRAM_28_DMWIDTH),
        .M_AXIS_BRAM_29_DMWIDTH(M_AXIS_BRAM_29_DMWIDTH),
        .M_AXIS_BRAM_30_DMWIDTH(M_AXIS_BRAM_30_DMWIDTH),
        .M_AXIS_BRAM_31_DMWIDTH(M_AXIS_BRAM_31_DMWIDTH),
        .M_AXIS_BRAM_32_DMWIDTH(M_AXIS_BRAM_32_DMWIDTH),
        .M_AXIS_BRAM_33_DMWIDTH(M_AXIS_BRAM_33_DMWIDTH),
        .M_AXIS_BRAM_34_DMWIDTH(M_AXIS_BRAM_34_DMWIDTH),
        .M_AXIS_BRAM_35_DMWIDTH(M_AXIS_BRAM_35_DMWIDTH),
        .M_AXIS_BRAM_36_DMWIDTH(M_AXIS_BRAM_36_DMWIDTH),
        .M_AXIS_BRAM_37_DMWIDTH(M_AXIS_BRAM_37_DMWIDTH),
        .M_AXIS_BRAM_38_DMWIDTH(M_AXIS_BRAM_38_DMWIDTH),
        .M_AXIS_BRAM_39_DMWIDTH(M_AXIS_BRAM_39_DMWIDTH),
        .M_AXIS_BRAM_40_DMWIDTH(M_AXIS_BRAM_40_DMWIDTH),
        .M_AXIS_BRAM_41_DMWIDTH(M_AXIS_BRAM_41_DMWIDTH),
        .M_AXIS_BRAM_42_DMWIDTH(M_AXIS_BRAM_42_DMWIDTH),
        .M_AXIS_BRAM_43_DMWIDTH(M_AXIS_BRAM_43_DMWIDTH),
        .M_AXIS_BRAM_44_DMWIDTH(M_AXIS_BRAM_44_DMWIDTH),
        .M_AXIS_BRAM_45_DMWIDTH(M_AXIS_BRAM_45_DMWIDTH),
        .M_AXIS_BRAM_46_DMWIDTH(M_AXIS_BRAM_46_DMWIDTH),
        .M_AXIS_BRAM_47_DMWIDTH(M_AXIS_BRAM_47_DMWIDTH),
        .M_AXIS_BRAM_48_DMWIDTH(M_AXIS_BRAM_48_DMWIDTH),
        .M_AXIS_BRAM_49_DMWIDTH(M_AXIS_BRAM_49_DMWIDTH),
        .M_AXIS_BRAM_50_DMWIDTH(M_AXIS_BRAM_50_DMWIDTH),
        .M_AXIS_BRAM_51_DMWIDTH(M_AXIS_BRAM_51_DMWIDTH),
        .M_AXIS_BRAM_52_DMWIDTH(M_AXIS_BRAM_52_DMWIDTH),
        .M_AXIS_BRAM_53_DMWIDTH(M_AXIS_BRAM_53_DMWIDTH),
        .M_AXIS_BRAM_54_DMWIDTH(M_AXIS_BRAM_54_DMWIDTH),
        .M_AXIS_BRAM_55_DMWIDTH(M_AXIS_BRAM_55_DMWIDTH),
        .M_AXIS_BRAM_56_DMWIDTH(M_AXIS_BRAM_56_DMWIDTH),
        .M_AXIS_BRAM_57_DMWIDTH(M_AXIS_BRAM_57_DMWIDTH),
        .M_AXIS_BRAM_58_DMWIDTH(M_AXIS_BRAM_58_DMWIDTH),
        .M_AXIS_BRAM_59_DMWIDTH(M_AXIS_BRAM_59_DMWIDTH),
        .M_AXIS_BRAM_60_DMWIDTH(M_AXIS_BRAM_60_DMWIDTH),
        .M_AXIS_BRAM_61_DMWIDTH(M_AXIS_BRAM_61_DMWIDTH),
        .M_AXIS_BRAM_62_DMWIDTH(M_AXIS_BRAM_62_DMWIDTH),
        .M_AXIS_BRAM_63_DMWIDTH(M_AXIS_BRAM_63_DMWIDTH),
        .M_AXIS_BRAM_64_DMWIDTH(M_AXIS_BRAM_64_DMWIDTH),
        .M_AXIS_BRAM_65_DMWIDTH(M_AXIS_BRAM_65_DMWIDTH),
        .M_AXIS_BRAM_66_DMWIDTH(M_AXIS_BRAM_66_DMWIDTH),
        .M_AXIS_BRAM_67_DMWIDTH(M_AXIS_BRAM_67_DMWIDTH),
        .M_AXIS_BRAM_68_DMWIDTH(M_AXIS_BRAM_68_DMWIDTH),
        .M_AXIS_BRAM_69_DMWIDTH(M_AXIS_BRAM_69_DMWIDTH),
        .M_AXIS_BRAM_70_DMWIDTH(M_AXIS_BRAM_70_DMWIDTH),
        .M_AXIS_BRAM_71_DMWIDTH(M_AXIS_BRAM_71_DMWIDTH),
        .M_AXIS_BRAM_72_DMWIDTH(M_AXIS_BRAM_72_DMWIDTH),
        .M_AXIS_BRAM_73_DMWIDTH(M_AXIS_BRAM_73_DMWIDTH),
        .M_AXIS_BRAM_74_DMWIDTH(M_AXIS_BRAM_74_DMWIDTH),
        .M_AXIS_BRAM_75_DMWIDTH(M_AXIS_BRAM_75_DMWIDTH),
        .M_AXIS_BRAM_76_DMWIDTH(M_AXIS_BRAM_76_DMWIDTH),
        .M_AXIS_BRAM_77_DMWIDTH(M_AXIS_BRAM_77_DMWIDTH),
        .M_AXIS_BRAM_78_DMWIDTH(M_AXIS_BRAM_78_DMWIDTH),
        .M_AXIS_BRAM_79_DMWIDTH(M_AXIS_BRAM_79_DMWIDTH),
        .M_AXIS_BRAM_80_DMWIDTH(M_AXIS_BRAM_80_DMWIDTH),
        .M_AXIS_BRAM_81_DMWIDTH(M_AXIS_BRAM_81_DMWIDTH),
        .M_AXIS_BRAM_82_DMWIDTH(M_AXIS_BRAM_82_DMWIDTH),
        .M_AXIS_BRAM_83_DMWIDTH(M_AXIS_BRAM_83_DMWIDTH),
        .M_AXIS_BRAM_84_DMWIDTH(M_AXIS_BRAM_84_DMWIDTH),
        .M_AXIS_BRAM_85_DMWIDTH(M_AXIS_BRAM_85_DMWIDTH),
        .M_AXIS_BRAM_86_DMWIDTH(M_AXIS_BRAM_86_DMWIDTH),
        .M_AXIS_BRAM_87_DMWIDTH(M_AXIS_BRAM_87_DMWIDTH),
        .M_AXIS_BRAM_88_DMWIDTH(M_AXIS_BRAM_88_DMWIDTH),
        .M_AXIS_BRAM_89_DMWIDTH(M_AXIS_BRAM_89_DMWIDTH),
        .M_AXIS_BRAM_90_DMWIDTH(M_AXIS_BRAM_90_DMWIDTH),
        .M_AXIS_BRAM_91_DMWIDTH(M_AXIS_BRAM_91_DMWIDTH),
        .M_AXIS_BRAM_92_DMWIDTH(M_AXIS_BRAM_92_DMWIDTH),
        .M_AXIS_BRAM_93_DMWIDTH(M_AXIS_BRAM_93_DMWIDTH),
        .M_AXIS_BRAM_94_DMWIDTH(M_AXIS_BRAM_94_DMWIDTH),
        .M_AXIS_BRAM_95_DMWIDTH(M_AXIS_BRAM_95_DMWIDTH),
        .M_AXIS_BRAM_96_DMWIDTH(M_AXIS_BRAM_96_DMWIDTH),
        .M_AXIS_BRAM_97_DMWIDTH(M_AXIS_BRAM_97_DMWIDTH),
        .M_AXIS_BRAM_98_DMWIDTH(M_AXIS_BRAM_98_DMWIDTH),
        .M_AXIS_BRAM_99_DMWIDTH(M_AXIS_BRAM_99_DMWIDTH),
        .M_AXIS_BRAM_100_DMWIDTH(M_AXIS_BRAM_100_DMWIDTH),
        .M_AXIS_BRAM_101_DMWIDTH(M_AXIS_BRAM_101_DMWIDTH),
        .M_AXIS_BRAM_102_DMWIDTH(M_AXIS_BRAM_102_DMWIDTH),
        .M_AXIS_BRAM_103_DMWIDTH(M_AXIS_BRAM_103_DMWIDTH),
        .M_AXIS_BRAM_104_DMWIDTH(M_AXIS_BRAM_104_DMWIDTH),
        .M_AXIS_BRAM_105_DMWIDTH(M_AXIS_BRAM_105_DMWIDTH),
        .M_AXIS_BRAM_106_DMWIDTH(M_AXIS_BRAM_106_DMWIDTH),
        .M_AXIS_BRAM_107_DMWIDTH(M_AXIS_BRAM_107_DMWIDTH),
        .M_AXIS_BRAM_108_DMWIDTH(M_AXIS_BRAM_108_DMWIDTH),
        .M_AXIS_BRAM_109_DMWIDTH(M_AXIS_BRAM_109_DMWIDTH),
        .M_AXIS_BRAM_110_DMWIDTH(M_AXIS_BRAM_110_DMWIDTH),
        .M_AXIS_BRAM_111_DMWIDTH(M_AXIS_BRAM_111_DMWIDTH),
        .M_AXIS_BRAM_112_DMWIDTH(M_AXIS_BRAM_112_DMWIDTH),
        .M_AXIS_BRAM_113_DMWIDTH(M_AXIS_BRAM_113_DMWIDTH),
        .M_AXIS_BRAM_114_DMWIDTH(M_AXIS_BRAM_114_DMWIDTH),
        .M_AXIS_BRAM_115_DMWIDTH(M_AXIS_BRAM_115_DMWIDTH),
        .M_AXIS_BRAM_116_DMWIDTH(M_AXIS_BRAM_116_DMWIDTH),
        .M_AXIS_BRAM_117_DMWIDTH(M_AXIS_BRAM_117_DMWIDTH),
        .M_AXIS_BRAM_118_DMWIDTH(M_AXIS_BRAM_118_DMWIDTH),
        .M_AXIS_BRAM_119_DMWIDTH(M_AXIS_BRAM_119_DMWIDTH),
        .M_AXIS_BRAM_120_DMWIDTH(M_AXIS_BRAM_120_DMWIDTH),
        .M_AXIS_BRAM_121_DMWIDTH(M_AXIS_BRAM_121_DMWIDTH),
        .M_AXIS_BRAM_122_DMWIDTH(M_AXIS_BRAM_122_DMWIDTH),
        .M_AXIS_BRAM_123_DMWIDTH(M_AXIS_BRAM_123_DMWIDTH),
        .M_AXIS_BRAM_124_DMWIDTH(M_AXIS_BRAM_124_DMWIDTH),
        .M_AXIS_BRAM_125_DMWIDTH(M_AXIS_BRAM_125_DMWIDTH),
        .M_AXIS_BRAM_126_DMWIDTH(M_AXIS_BRAM_126_DMWIDTH),
        .M_AXIS_BRAM_127_DMWIDTH(M_AXIS_BRAM_127_DMWIDTH),
        .M_AXIS_BRAM_0_IS_ASYNC(M_AXIS_BRAM_0_IS_ASYNC),
        .M_AXIS_BRAM_1_IS_ASYNC(M_AXIS_BRAM_1_IS_ASYNC),
        .M_AXIS_BRAM_2_IS_ASYNC(M_AXIS_BRAM_2_IS_ASYNC),
        .M_AXIS_BRAM_3_IS_ASYNC(M_AXIS_BRAM_3_IS_ASYNC),
        .M_AXIS_BRAM_4_IS_ASYNC(M_AXIS_BRAM_4_IS_ASYNC),
        .M_AXIS_BRAM_5_IS_ASYNC(M_AXIS_BRAM_5_IS_ASYNC),
        .M_AXIS_BRAM_6_IS_ASYNC(M_AXIS_BRAM_6_IS_ASYNC),
        .M_AXIS_BRAM_7_IS_ASYNC(M_AXIS_BRAM_7_IS_ASYNC),
        .M_AXIS_BRAM_8_IS_ASYNC(M_AXIS_BRAM_8_IS_ASYNC),
        .M_AXIS_BRAM_9_IS_ASYNC(M_AXIS_BRAM_9_IS_ASYNC),
        .M_AXIS_BRAM_10_IS_ASYNC(M_AXIS_BRAM_10_IS_ASYNC),
        .M_AXIS_BRAM_11_IS_ASYNC(M_AXIS_BRAM_11_IS_ASYNC),
        .M_AXIS_BRAM_12_IS_ASYNC(M_AXIS_BRAM_12_IS_ASYNC),
        .M_AXIS_BRAM_13_IS_ASYNC(M_AXIS_BRAM_13_IS_ASYNC),
        .M_AXIS_BRAM_14_IS_ASYNC(M_AXIS_BRAM_14_IS_ASYNC),
        .M_AXIS_BRAM_15_IS_ASYNC(M_AXIS_BRAM_15_IS_ASYNC),
        .M_AXIS_BRAM_16_IS_ASYNC(M_AXIS_BRAM_16_IS_ASYNC),
        .M_AXIS_BRAM_17_IS_ASYNC(M_AXIS_BRAM_17_IS_ASYNC),
        .M_AXIS_BRAM_18_IS_ASYNC(M_AXIS_BRAM_18_IS_ASYNC),
        .M_AXIS_BRAM_19_IS_ASYNC(M_AXIS_BRAM_19_IS_ASYNC),
        .M_AXIS_BRAM_20_IS_ASYNC(M_AXIS_BRAM_20_IS_ASYNC),
        .M_AXIS_BRAM_21_IS_ASYNC(M_AXIS_BRAM_21_IS_ASYNC),
        .M_AXIS_BRAM_22_IS_ASYNC(M_AXIS_BRAM_22_IS_ASYNC),
        .M_AXIS_BRAM_23_IS_ASYNC(M_AXIS_BRAM_23_IS_ASYNC),
        .M_AXIS_BRAM_24_IS_ASYNC(M_AXIS_BRAM_24_IS_ASYNC),
        .M_AXIS_BRAM_25_IS_ASYNC(M_AXIS_BRAM_25_IS_ASYNC),
        .M_AXIS_BRAM_26_IS_ASYNC(M_AXIS_BRAM_26_IS_ASYNC),
        .M_AXIS_BRAM_27_IS_ASYNC(M_AXIS_BRAM_27_IS_ASYNC),
        .M_AXIS_BRAM_28_IS_ASYNC(M_AXIS_BRAM_28_IS_ASYNC),
        .M_AXIS_BRAM_29_IS_ASYNC(M_AXIS_BRAM_29_IS_ASYNC),
        .M_AXIS_BRAM_30_IS_ASYNC(M_AXIS_BRAM_30_IS_ASYNC),
        .M_AXIS_BRAM_31_IS_ASYNC(M_AXIS_BRAM_31_IS_ASYNC),
        .M_AXIS_BRAM_32_IS_ASYNC(M_AXIS_BRAM_32_IS_ASYNC),
        .M_AXIS_BRAM_33_IS_ASYNC(M_AXIS_BRAM_33_IS_ASYNC),
        .M_AXIS_BRAM_34_IS_ASYNC(M_AXIS_BRAM_34_IS_ASYNC),
        .M_AXIS_BRAM_35_IS_ASYNC(M_AXIS_BRAM_35_IS_ASYNC),
        .M_AXIS_BRAM_36_IS_ASYNC(M_AXIS_BRAM_36_IS_ASYNC),
        .M_AXIS_BRAM_37_IS_ASYNC(M_AXIS_BRAM_37_IS_ASYNC),
        .M_AXIS_BRAM_38_IS_ASYNC(M_AXIS_BRAM_38_IS_ASYNC),
        .M_AXIS_BRAM_39_IS_ASYNC(M_AXIS_BRAM_39_IS_ASYNC),
        .M_AXIS_BRAM_40_IS_ASYNC(M_AXIS_BRAM_40_IS_ASYNC),
        .M_AXIS_BRAM_41_IS_ASYNC(M_AXIS_BRAM_41_IS_ASYNC),
        .M_AXIS_BRAM_42_IS_ASYNC(M_AXIS_BRAM_42_IS_ASYNC),
        .M_AXIS_BRAM_43_IS_ASYNC(M_AXIS_BRAM_43_IS_ASYNC),
        .M_AXIS_BRAM_44_IS_ASYNC(M_AXIS_BRAM_44_IS_ASYNC),
        .M_AXIS_BRAM_45_IS_ASYNC(M_AXIS_BRAM_45_IS_ASYNC),
        .M_AXIS_BRAM_46_IS_ASYNC(M_AXIS_BRAM_46_IS_ASYNC),
        .M_AXIS_BRAM_47_IS_ASYNC(M_AXIS_BRAM_47_IS_ASYNC),
        .M_AXIS_BRAM_48_IS_ASYNC(M_AXIS_BRAM_48_IS_ASYNC),
        .M_AXIS_BRAM_49_IS_ASYNC(M_AXIS_BRAM_49_IS_ASYNC),
        .M_AXIS_BRAM_50_IS_ASYNC(M_AXIS_BRAM_50_IS_ASYNC),
        .M_AXIS_BRAM_51_IS_ASYNC(M_AXIS_BRAM_51_IS_ASYNC),
        .M_AXIS_BRAM_52_IS_ASYNC(M_AXIS_BRAM_52_IS_ASYNC),
        .M_AXIS_BRAM_53_IS_ASYNC(M_AXIS_BRAM_53_IS_ASYNC),
        .M_AXIS_BRAM_54_IS_ASYNC(M_AXIS_BRAM_54_IS_ASYNC),
        .M_AXIS_BRAM_55_IS_ASYNC(M_AXIS_BRAM_55_IS_ASYNC),
        .M_AXIS_BRAM_56_IS_ASYNC(M_AXIS_BRAM_56_IS_ASYNC),
        .M_AXIS_BRAM_57_IS_ASYNC(M_AXIS_BRAM_57_IS_ASYNC),
        .M_AXIS_BRAM_58_IS_ASYNC(M_AXIS_BRAM_58_IS_ASYNC),
        .M_AXIS_BRAM_59_IS_ASYNC(M_AXIS_BRAM_59_IS_ASYNC),
        .M_AXIS_BRAM_60_IS_ASYNC(M_AXIS_BRAM_60_IS_ASYNC),
        .M_AXIS_BRAM_61_IS_ASYNC(M_AXIS_BRAM_61_IS_ASYNC),
        .M_AXIS_BRAM_62_IS_ASYNC(M_AXIS_BRAM_62_IS_ASYNC),
        .M_AXIS_BRAM_63_IS_ASYNC(M_AXIS_BRAM_63_IS_ASYNC),
        .M_AXIS_BRAM_64_IS_ASYNC(M_AXIS_BRAM_64_IS_ASYNC),
        .M_AXIS_BRAM_65_IS_ASYNC(M_AXIS_BRAM_65_IS_ASYNC),
        .M_AXIS_BRAM_66_IS_ASYNC(M_AXIS_BRAM_66_IS_ASYNC),
        .M_AXIS_BRAM_67_IS_ASYNC(M_AXIS_BRAM_67_IS_ASYNC),
        .M_AXIS_BRAM_68_IS_ASYNC(M_AXIS_BRAM_68_IS_ASYNC),
        .M_AXIS_BRAM_69_IS_ASYNC(M_AXIS_BRAM_69_IS_ASYNC),
        .M_AXIS_BRAM_70_IS_ASYNC(M_AXIS_BRAM_70_IS_ASYNC),
        .M_AXIS_BRAM_71_IS_ASYNC(M_AXIS_BRAM_71_IS_ASYNC),
        .M_AXIS_BRAM_72_IS_ASYNC(M_AXIS_BRAM_72_IS_ASYNC),
        .M_AXIS_BRAM_73_IS_ASYNC(M_AXIS_BRAM_73_IS_ASYNC),
        .M_AXIS_BRAM_74_IS_ASYNC(M_AXIS_BRAM_74_IS_ASYNC),
        .M_AXIS_BRAM_75_IS_ASYNC(M_AXIS_BRAM_75_IS_ASYNC),
        .M_AXIS_BRAM_76_IS_ASYNC(M_AXIS_BRAM_76_IS_ASYNC),
        .M_AXIS_BRAM_77_IS_ASYNC(M_AXIS_BRAM_77_IS_ASYNC),
        .M_AXIS_BRAM_78_IS_ASYNC(M_AXIS_BRAM_78_IS_ASYNC),
        .M_AXIS_BRAM_79_IS_ASYNC(M_AXIS_BRAM_79_IS_ASYNC),
        .M_AXIS_BRAM_80_IS_ASYNC(M_AXIS_BRAM_80_IS_ASYNC),
        .M_AXIS_BRAM_81_IS_ASYNC(M_AXIS_BRAM_81_IS_ASYNC),
        .M_AXIS_BRAM_82_IS_ASYNC(M_AXIS_BRAM_82_IS_ASYNC),
        .M_AXIS_BRAM_83_IS_ASYNC(M_AXIS_BRAM_83_IS_ASYNC),
        .M_AXIS_BRAM_84_IS_ASYNC(M_AXIS_BRAM_84_IS_ASYNC),
        .M_AXIS_BRAM_85_IS_ASYNC(M_AXIS_BRAM_85_IS_ASYNC),
        .M_AXIS_BRAM_86_IS_ASYNC(M_AXIS_BRAM_86_IS_ASYNC),
        .M_AXIS_BRAM_87_IS_ASYNC(M_AXIS_BRAM_87_IS_ASYNC),
        .M_AXIS_BRAM_88_IS_ASYNC(M_AXIS_BRAM_88_IS_ASYNC),
        .M_AXIS_BRAM_89_IS_ASYNC(M_AXIS_BRAM_89_IS_ASYNC),
        .M_AXIS_BRAM_90_IS_ASYNC(M_AXIS_BRAM_90_IS_ASYNC),
        .M_AXIS_BRAM_91_IS_ASYNC(M_AXIS_BRAM_91_IS_ASYNC),
        .M_AXIS_BRAM_92_IS_ASYNC(M_AXIS_BRAM_92_IS_ASYNC),
        .M_AXIS_BRAM_93_IS_ASYNC(M_AXIS_BRAM_93_IS_ASYNC),
        .M_AXIS_BRAM_94_IS_ASYNC(M_AXIS_BRAM_94_IS_ASYNC),
        .M_AXIS_BRAM_95_IS_ASYNC(M_AXIS_BRAM_95_IS_ASYNC),
        .M_AXIS_BRAM_96_IS_ASYNC(M_AXIS_BRAM_96_IS_ASYNC),
        .M_AXIS_BRAM_97_IS_ASYNC(M_AXIS_BRAM_97_IS_ASYNC),
        .M_AXIS_BRAM_98_IS_ASYNC(M_AXIS_BRAM_98_IS_ASYNC),
        .M_AXIS_BRAM_99_IS_ASYNC(M_AXIS_BRAM_99_IS_ASYNC),
        .M_AXIS_BRAM_100_IS_ASYNC(M_AXIS_BRAM_100_IS_ASYNC),
        .M_AXIS_BRAM_101_IS_ASYNC(M_AXIS_BRAM_101_IS_ASYNC),
        .M_AXIS_BRAM_102_IS_ASYNC(M_AXIS_BRAM_102_IS_ASYNC),
        .M_AXIS_BRAM_103_IS_ASYNC(M_AXIS_BRAM_103_IS_ASYNC),
        .M_AXIS_BRAM_104_IS_ASYNC(M_AXIS_BRAM_104_IS_ASYNC),
        .M_AXIS_BRAM_105_IS_ASYNC(M_AXIS_BRAM_105_IS_ASYNC),
        .M_AXIS_BRAM_106_IS_ASYNC(M_AXIS_BRAM_106_IS_ASYNC),
        .M_AXIS_BRAM_107_IS_ASYNC(M_AXIS_BRAM_107_IS_ASYNC),
        .M_AXIS_BRAM_108_IS_ASYNC(M_AXIS_BRAM_108_IS_ASYNC),
        .M_AXIS_BRAM_109_IS_ASYNC(M_AXIS_BRAM_109_IS_ASYNC),
        .M_AXIS_BRAM_110_IS_ASYNC(M_AXIS_BRAM_110_IS_ASYNC),
        .M_AXIS_BRAM_111_IS_ASYNC(M_AXIS_BRAM_111_IS_ASYNC),
        .M_AXIS_BRAM_112_IS_ASYNC(M_AXIS_BRAM_112_IS_ASYNC),
        .M_AXIS_BRAM_113_IS_ASYNC(M_AXIS_BRAM_113_IS_ASYNC),
        .M_AXIS_BRAM_114_IS_ASYNC(M_AXIS_BRAM_114_IS_ASYNC),
        .M_AXIS_BRAM_115_IS_ASYNC(M_AXIS_BRAM_115_IS_ASYNC),
        .M_AXIS_BRAM_116_IS_ASYNC(M_AXIS_BRAM_116_IS_ASYNC),
        .M_AXIS_BRAM_117_IS_ASYNC(M_AXIS_BRAM_117_IS_ASYNC),
        .M_AXIS_BRAM_118_IS_ASYNC(M_AXIS_BRAM_118_IS_ASYNC),
        .M_AXIS_BRAM_119_IS_ASYNC(M_AXIS_BRAM_119_IS_ASYNC),
        .M_AXIS_BRAM_120_IS_ASYNC(M_AXIS_BRAM_120_IS_ASYNC),
        .M_AXIS_BRAM_121_IS_ASYNC(M_AXIS_BRAM_121_IS_ASYNC),
        .M_AXIS_BRAM_122_IS_ASYNC(M_AXIS_BRAM_122_IS_ASYNC),
        .M_AXIS_BRAM_123_IS_ASYNC(M_AXIS_BRAM_123_IS_ASYNC),
        .M_AXIS_BRAM_124_IS_ASYNC(M_AXIS_BRAM_124_IS_ASYNC),
        .M_AXIS_BRAM_125_IS_ASYNC(M_AXIS_BRAM_125_IS_ASYNC),
        .M_AXIS_BRAM_126_IS_ASYNC(M_AXIS_BRAM_126_IS_ASYNC),
        .M_AXIS_BRAM_127_IS_ASYNC(M_AXIS_BRAM_127_IS_ASYNC),
        .M_AXIS_BRAM_0_PORTS(M_AXIS_BRAM_0_PORTS),
        .M_AXIS_BRAM_1_PORTS(M_AXIS_BRAM_1_PORTS),
        .M_AXIS_BRAM_2_PORTS(M_AXIS_BRAM_2_PORTS),
        .M_AXIS_BRAM_3_PORTS(M_AXIS_BRAM_3_PORTS),
        .M_AXIS_BRAM_4_PORTS(M_AXIS_BRAM_4_PORTS),
        .M_AXIS_BRAM_5_PORTS(M_AXIS_BRAM_5_PORTS),
        .M_AXIS_BRAM_6_PORTS(M_AXIS_BRAM_6_PORTS),
        .M_AXIS_BRAM_7_PORTS(M_AXIS_BRAM_7_PORTS),
        .M_AXIS_BRAM_8_PORTS(M_AXIS_BRAM_8_PORTS),
        .M_AXIS_BRAM_9_PORTS(M_AXIS_BRAM_9_PORTS),
        .M_AXIS_BRAM_10_PORTS(M_AXIS_BRAM_10_PORTS),
        .M_AXIS_BRAM_11_PORTS(M_AXIS_BRAM_11_PORTS),
        .M_AXIS_BRAM_12_PORTS(M_AXIS_BRAM_12_PORTS),
        .M_AXIS_BRAM_13_PORTS(M_AXIS_BRAM_13_PORTS),
        .M_AXIS_BRAM_14_PORTS(M_AXIS_BRAM_14_PORTS),
        .M_AXIS_BRAM_15_PORTS(M_AXIS_BRAM_15_PORTS),
        .M_AXIS_BRAM_16_PORTS(M_AXIS_BRAM_16_PORTS),
        .M_AXIS_BRAM_17_PORTS(M_AXIS_BRAM_17_PORTS),
        .M_AXIS_BRAM_18_PORTS(M_AXIS_BRAM_18_PORTS),
        .M_AXIS_BRAM_19_PORTS(M_AXIS_BRAM_19_PORTS),
        .M_AXIS_BRAM_20_PORTS(M_AXIS_BRAM_20_PORTS),
        .M_AXIS_BRAM_21_PORTS(M_AXIS_BRAM_21_PORTS),
        .M_AXIS_BRAM_22_PORTS(M_AXIS_BRAM_22_PORTS),
        .M_AXIS_BRAM_23_PORTS(M_AXIS_BRAM_23_PORTS),
        .M_AXIS_BRAM_24_PORTS(M_AXIS_BRAM_24_PORTS),
        .M_AXIS_BRAM_25_PORTS(M_AXIS_BRAM_25_PORTS),
        .M_AXIS_BRAM_26_PORTS(M_AXIS_BRAM_26_PORTS),
        .M_AXIS_BRAM_27_PORTS(M_AXIS_BRAM_27_PORTS),
        .M_AXIS_BRAM_28_PORTS(M_AXIS_BRAM_28_PORTS),
        .M_AXIS_BRAM_29_PORTS(M_AXIS_BRAM_29_PORTS),
        .M_AXIS_BRAM_30_PORTS(M_AXIS_BRAM_30_PORTS),
        .M_AXIS_BRAM_31_PORTS(M_AXIS_BRAM_31_PORTS),
        .M_AXIS_BRAM_32_PORTS(M_AXIS_BRAM_32_PORTS),
        .M_AXIS_BRAM_33_PORTS(M_AXIS_BRAM_33_PORTS),
        .M_AXIS_BRAM_34_PORTS(M_AXIS_BRAM_34_PORTS),
        .M_AXIS_BRAM_35_PORTS(M_AXIS_BRAM_35_PORTS),
        .M_AXIS_BRAM_36_PORTS(M_AXIS_BRAM_36_PORTS),
        .M_AXIS_BRAM_37_PORTS(M_AXIS_BRAM_37_PORTS),
        .M_AXIS_BRAM_38_PORTS(M_AXIS_BRAM_38_PORTS),
        .M_AXIS_BRAM_39_PORTS(M_AXIS_BRAM_39_PORTS),
        .M_AXIS_BRAM_40_PORTS(M_AXIS_BRAM_40_PORTS),
        .M_AXIS_BRAM_41_PORTS(M_AXIS_BRAM_41_PORTS),
        .M_AXIS_BRAM_42_PORTS(M_AXIS_BRAM_42_PORTS),
        .M_AXIS_BRAM_43_PORTS(M_AXIS_BRAM_43_PORTS),
        .M_AXIS_BRAM_44_PORTS(M_AXIS_BRAM_44_PORTS),
        .M_AXIS_BRAM_45_PORTS(M_AXIS_BRAM_45_PORTS),
        .M_AXIS_BRAM_46_PORTS(M_AXIS_BRAM_46_PORTS),
        .M_AXIS_BRAM_47_PORTS(M_AXIS_BRAM_47_PORTS),
        .M_AXIS_BRAM_48_PORTS(M_AXIS_BRAM_48_PORTS),
        .M_AXIS_BRAM_49_PORTS(M_AXIS_BRAM_49_PORTS),
        .M_AXIS_BRAM_50_PORTS(M_AXIS_BRAM_50_PORTS),
        .M_AXIS_BRAM_51_PORTS(M_AXIS_BRAM_51_PORTS),
        .M_AXIS_BRAM_52_PORTS(M_AXIS_BRAM_52_PORTS),
        .M_AXIS_BRAM_53_PORTS(M_AXIS_BRAM_53_PORTS),
        .M_AXIS_BRAM_54_PORTS(M_AXIS_BRAM_54_PORTS),
        .M_AXIS_BRAM_55_PORTS(M_AXIS_BRAM_55_PORTS),
        .M_AXIS_BRAM_56_PORTS(M_AXIS_BRAM_56_PORTS),
        .M_AXIS_BRAM_57_PORTS(M_AXIS_BRAM_57_PORTS),
        .M_AXIS_BRAM_58_PORTS(M_AXIS_BRAM_58_PORTS),
        .M_AXIS_BRAM_59_PORTS(M_AXIS_BRAM_59_PORTS),
        .M_AXIS_BRAM_60_PORTS(M_AXIS_BRAM_60_PORTS),
        .M_AXIS_BRAM_61_PORTS(M_AXIS_BRAM_61_PORTS),
        .M_AXIS_BRAM_62_PORTS(M_AXIS_BRAM_62_PORTS),
        .M_AXIS_BRAM_63_PORTS(M_AXIS_BRAM_63_PORTS),
        .M_AXIS_BRAM_64_PORTS(M_AXIS_BRAM_64_PORTS),
        .M_AXIS_BRAM_65_PORTS(M_AXIS_BRAM_65_PORTS),
        .M_AXIS_BRAM_66_PORTS(M_AXIS_BRAM_66_PORTS),
        .M_AXIS_BRAM_67_PORTS(M_AXIS_BRAM_67_PORTS),
        .M_AXIS_BRAM_68_PORTS(M_AXIS_BRAM_68_PORTS),
        .M_AXIS_BRAM_69_PORTS(M_AXIS_BRAM_69_PORTS),
        .M_AXIS_BRAM_70_PORTS(M_AXIS_BRAM_70_PORTS),
        .M_AXIS_BRAM_71_PORTS(M_AXIS_BRAM_71_PORTS),
        .M_AXIS_BRAM_72_PORTS(M_AXIS_BRAM_72_PORTS),
        .M_AXIS_BRAM_73_PORTS(M_AXIS_BRAM_73_PORTS),
        .M_AXIS_BRAM_74_PORTS(M_AXIS_BRAM_74_PORTS),
        .M_AXIS_BRAM_75_PORTS(M_AXIS_BRAM_75_PORTS),
        .M_AXIS_BRAM_76_PORTS(M_AXIS_BRAM_76_PORTS),
        .M_AXIS_BRAM_77_PORTS(M_AXIS_BRAM_77_PORTS),
        .M_AXIS_BRAM_78_PORTS(M_AXIS_BRAM_78_PORTS),
        .M_AXIS_BRAM_79_PORTS(M_AXIS_BRAM_79_PORTS),
        .M_AXIS_BRAM_80_PORTS(M_AXIS_BRAM_80_PORTS),
        .M_AXIS_BRAM_81_PORTS(M_AXIS_BRAM_81_PORTS),
        .M_AXIS_BRAM_82_PORTS(M_AXIS_BRAM_82_PORTS),
        .M_AXIS_BRAM_83_PORTS(M_AXIS_BRAM_83_PORTS),
        .M_AXIS_BRAM_84_PORTS(M_AXIS_BRAM_84_PORTS),
        .M_AXIS_BRAM_85_PORTS(M_AXIS_BRAM_85_PORTS),
        .M_AXIS_BRAM_86_PORTS(M_AXIS_BRAM_86_PORTS),
        .M_AXIS_BRAM_87_PORTS(M_AXIS_BRAM_87_PORTS),
        .M_AXIS_BRAM_88_PORTS(M_AXIS_BRAM_88_PORTS),
        .M_AXIS_BRAM_89_PORTS(M_AXIS_BRAM_89_PORTS),
        .M_AXIS_BRAM_90_PORTS(M_AXIS_BRAM_90_PORTS),
        .M_AXIS_BRAM_91_PORTS(M_AXIS_BRAM_91_PORTS),
        .M_AXIS_BRAM_92_PORTS(M_AXIS_BRAM_92_PORTS),
        .M_AXIS_BRAM_93_PORTS(M_AXIS_BRAM_93_PORTS),
        .M_AXIS_BRAM_94_PORTS(M_AXIS_BRAM_94_PORTS),
        .M_AXIS_BRAM_95_PORTS(M_AXIS_BRAM_95_PORTS),
        .M_AXIS_BRAM_96_PORTS(M_AXIS_BRAM_96_PORTS),
        .M_AXIS_BRAM_97_PORTS(M_AXIS_BRAM_97_PORTS),
        .M_AXIS_BRAM_98_PORTS(M_AXIS_BRAM_98_PORTS),
        .M_AXIS_BRAM_99_PORTS(M_AXIS_BRAM_99_PORTS),
        .M_AXIS_BRAM_100_PORTS(M_AXIS_BRAM_100_PORTS),
        .M_AXIS_BRAM_101_PORTS(M_AXIS_BRAM_101_PORTS),
        .M_AXIS_BRAM_102_PORTS(M_AXIS_BRAM_102_PORTS),
        .M_AXIS_BRAM_103_PORTS(M_AXIS_BRAM_103_PORTS),
        .M_AXIS_BRAM_104_PORTS(M_AXIS_BRAM_104_PORTS),
        .M_AXIS_BRAM_105_PORTS(M_AXIS_BRAM_105_PORTS),
        .M_AXIS_BRAM_106_PORTS(M_AXIS_BRAM_106_PORTS),
        .M_AXIS_BRAM_107_PORTS(M_AXIS_BRAM_107_PORTS),
        .M_AXIS_BRAM_108_PORTS(M_AXIS_BRAM_108_PORTS),
        .M_AXIS_BRAM_109_PORTS(M_AXIS_BRAM_109_PORTS),
        .M_AXIS_BRAM_110_PORTS(M_AXIS_BRAM_110_PORTS),
        .M_AXIS_BRAM_111_PORTS(M_AXIS_BRAM_111_PORTS),
        .M_AXIS_BRAM_112_PORTS(M_AXIS_BRAM_112_PORTS),
        .M_AXIS_BRAM_113_PORTS(M_AXIS_BRAM_113_PORTS),
        .M_AXIS_BRAM_114_PORTS(M_AXIS_BRAM_114_PORTS),
        .M_AXIS_BRAM_115_PORTS(M_AXIS_BRAM_115_PORTS),
        .M_AXIS_BRAM_116_PORTS(M_AXIS_BRAM_116_PORTS),
        .M_AXIS_BRAM_117_PORTS(M_AXIS_BRAM_117_PORTS),
        .M_AXIS_BRAM_118_PORTS(M_AXIS_BRAM_118_PORTS),
        .M_AXIS_BRAM_119_PORTS(M_AXIS_BRAM_119_PORTS),
        .M_AXIS_BRAM_120_PORTS(M_AXIS_BRAM_120_PORTS),
        .M_AXIS_BRAM_121_PORTS(M_AXIS_BRAM_121_PORTS),
        .M_AXIS_BRAM_122_PORTS(M_AXIS_BRAM_122_PORTS),
        .M_AXIS_BRAM_123_PORTS(M_AXIS_BRAM_123_PORTS),
        .M_AXIS_BRAM_124_PORTS(M_AXIS_BRAM_124_PORTS),
        .M_AXIS_BRAM_125_PORTS(M_AXIS_BRAM_125_PORTS),
        .M_AXIS_BRAM_126_PORTS(M_AXIS_BRAM_126_PORTS),
        .M_AXIS_BRAM_127_PORTS(M_AXIS_BRAM_127_PORTS),
        .M_AXIS_BRAM_0_MB_DEPTH(M_AXIS_BRAM_0_MB_DEPTH),
        .M_AXIS_BRAM_1_MB_DEPTH(M_AXIS_BRAM_1_MB_DEPTH),
        .M_AXIS_BRAM_2_MB_DEPTH(M_AXIS_BRAM_2_MB_DEPTH),
        .M_AXIS_BRAM_3_MB_DEPTH(M_AXIS_BRAM_3_MB_DEPTH),
        .M_AXIS_BRAM_4_MB_DEPTH(M_AXIS_BRAM_4_MB_DEPTH),
        .M_AXIS_BRAM_5_MB_DEPTH(M_AXIS_BRAM_5_MB_DEPTH),
        .M_AXIS_BRAM_6_MB_DEPTH(M_AXIS_BRAM_6_MB_DEPTH),
        .M_AXIS_BRAM_7_MB_DEPTH(M_AXIS_BRAM_7_MB_DEPTH),
        .M_AXIS_BRAM_8_MB_DEPTH(M_AXIS_BRAM_8_MB_DEPTH),
        .M_AXIS_BRAM_9_MB_DEPTH(M_AXIS_BRAM_9_MB_DEPTH),
        .M_AXIS_BRAM_10_MB_DEPTH(M_AXIS_BRAM_10_MB_DEPTH),
        .M_AXIS_BRAM_11_MB_DEPTH(M_AXIS_BRAM_11_MB_DEPTH),
        .M_AXIS_BRAM_12_MB_DEPTH(M_AXIS_BRAM_12_MB_DEPTH),
        .M_AXIS_BRAM_13_MB_DEPTH(M_AXIS_BRAM_13_MB_DEPTH),
        .M_AXIS_BRAM_14_MB_DEPTH(M_AXIS_BRAM_14_MB_DEPTH),
        .M_AXIS_BRAM_15_MB_DEPTH(M_AXIS_BRAM_15_MB_DEPTH),
        .M_AXIS_BRAM_16_MB_DEPTH(M_AXIS_BRAM_16_MB_DEPTH),
        .M_AXIS_BRAM_17_MB_DEPTH(M_AXIS_BRAM_17_MB_DEPTH),
        .M_AXIS_BRAM_18_MB_DEPTH(M_AXIS_BRAM_18_MB_DEPTH),
        .M_AXIS_BRAM_19_MB_DEPTH(M_AXIS_BRAM_19_MB_DEPTH),
        .M_AXIS_BRAM_20_MB_DEPTH(M_AXIS_BRAM_20_MB_DEPTH),
        .M_AXIS_BRAM_21_MB_DEPTH(M_AXIS_BRAM_21_MB_DEPTH),
        .M_AXIS_BRAM_22_MB_DEPTH(M_AXIS_BRAM_22_MB_DEPTH),
        .M_AXIS_BRAM_23_MB_DEPTH(M_AXIS_BRAM_23_MB_DEPTH),
        .M_AXIS_BRAM_24_MB_DEPTH(M_AXIS_BRAM_24_MB_DEPTH),
        .M_AXIS_BRAM_25_MB_DEPTH(M_AXIS_BRAM_25_MB_DEPTH),
        .M_AXIS_BRAM_26_MB_DEPTH(M_AXIS_BRAM_26_MB_DEPTH),
        .M_AXIS_BRAM_27_MB_DEPTH(M_AXIS_BRAM_27_MB_DEPTH),
        .M_AXIS_BRAM_28_MB_DEPTH(M_AXIS_BRAM_28_MB_DEPTH),
        .M_AXIS_BRAM_29_MB_DEPTH(M_AXIS_BRAM_29_MB_DEPTH),
        .M_AXIS_BRAM_30_MB_DEPTH(M_AXIS_BRAM_30_MB_DEPTH),
        .M_AXIS_BRAM_31_MB_DEPTH(M_AXIS_BRAM_31_MB_DEPTH),
        .M_AXIS_BRAM_32_MB_DEPTH(M_AXIS_BRAM_32_MB_DEPTH),
        .M_AXIS_BRAM_33_MB_DEPTH(M_AXIS_BRAM_33_MB_DEPTH),
        .M_AXIS_BRAM_34_MB_DEPTH(M_AXIS_BRAM_34_MB_DEPTH),
        .M_AXIS_BRAM_35_MB_DEPTH(M_AXIS_BRAM_35_MB_DEPTH),
        .M_AXIS_BRAM_36_MB_DEPTH(M_AXIS_BRAM_36_MB_DEPTH),
        .M_AXIS_BRAM_37_MB_DEPTH(M_AXIS_BRAM_37_MB_DEPTH),
        .M_AXIS_BRAM_38_MB_DEPTH(M_AXIS_BRAM_38_MB_DEPTH),
        .M_AXIS_BRAM_39_MB_DEPTH(M_AXIS_BRAM_39_MB_DEPTH),
        .M_AXIS_BRAM_40_MB_DEPTH(M_AXIS_BRAM_40_MB_DEPTH),
        .M_AXIS_BRAM_41_MB_DEPTH(M_AXIS_BRAM_41_MB_DEPTH),
        .M_AXIS_BRAM_42_MB_DEPTH(M_AXIS_BRAM_42_MB_DEPTH),
        .M_AXIS_BRAM_43_MB_DEPTH(M_AXIS_BRAM_43_MB_DEPTH),
        .M_AXIS_BRAM_44_MB_DEPTH(M_AXIS_BRAM_44_MB_DEPTH),
        .M_AXIS_BRAM_45_MB_DEPTH(M_AXIS_BRAM_45_MB_DEPTH),
        .M_AXIS_BRAM_46_MB_DEPTH(M_AXIS_BRAM_46_MB_DEPTH),
        .M_AXIS_BRAM_47_MB_DEPTH(M_AXIS_BRAM_47_MB_DEPTH),
        .M_AXIS_BRAM_48_MB_DEPTH(M_AXIS_BRAM_48_MB_DEPTH),
        .M_AXIS_BRAM_49_MB_DEPTH(M_AXIS_BRAM_49_MB_DEPTH),
        .M_AXIS_BRAM_50_MB_DEPTH(M_AXIS_BRAM_50_MB_DEPTH),
        .M_AXIS_BRAM_51_MB_DEPTH(M_AXIS_BRAM_51_MB_DEPTH),
        .M_AXIS_BRAM_52_MB_DEPTH(M_AXIS_BRAM_52_MB_DEPTH),
        .M_AXIS_BRAM_53_MB_DEPTH(M_AXIS_BRAM_53_MB_DEPTH),
        .M_AXIS_BRAM_54_MB_DEPTH(M_AXIS_BRAM_54_MB_DEPTH),
        .M_AXIS_BRAM_55_MB_DEPTH(M_AXIS_BRAM_55_MB_DEPTH),
        .M_AXIS_BRAM_56_MB_DEPTH(M_AXIS_BRAM_56_MB_DEPTH),
        .M_AXIS_BRAM_57_MB_DEPTH(M_AXIS_BRAM_57_MB_DEPTH),
        .M_AXIS_BRAM_58_MB_DEPTH(M_AXIS_BRAM_58_MB_DEPTH),
        .M_AXIS_BRAM_59_MB_DEPTH(M_AXIS_BRAM_59_MB_DEPTH),
        .M_AXIS_BRAM_60_MB_DEPTH(M_AXIS_BRAM_60_MB_DEPTH),
        .M_AXIS_BRAM_61_MB_DEPTH(M_AXIS_BRAM_61_MB_DEPTH),
        .M_AXIS_BRAM_62_MB_DEPTH(M_AXIS_BRAM_62_MB_DEPTH),
        .M_AXIS_BRAM_63_MB_DEPTH(M_AXIS_BRAM_63_MB_DEPTH),
        .M_AXIS_BRAM_64_MB_DEPTH(M_AXIS_BRAM_64_MB_DEPTH),
        .M_AXIS_BRAM_65_MB_DEPTH(M_AXIS_BRAM_65_MB_DEPTH),
        .M_AXIS_BRAM_66_MB_DEPTH(M_AXIS_BRAM_66_MB_DEPTH),
        .M_AXIS_BRAM_67_MB_DEPTH(M_AXIS_BRAM_67_MB_DEPTH),
        .M_AXIS_BRAM_68_MB_DEPTH(M_AXIS_BRAM_68_MB_DEPTH),
        .M_AXIS_BRAM_69_MB_DEPTH(M_AXIS_BRAM_69_MB_DEPTH),
        .M_AXIS_BRAM_70_MB_DEPTH(M_AXIS_BRAM_70_MB_DEPTH),
        .M_AXIS_BRAM_71_MB_DEPTH(M_AXIS_BRAM_71_MB_DEPTH),
        .M_AXIS_BRAM_72_MB_DEPTH(M_AXIS_BRAM_72_MB_DEPTH),
        .M_AXIS_BRAM_73_MB_DEPTH(M_AXIS_BRAM_73_MB_DEPTH),
        .M_AXIS_BRAM_74_MB_DEPTH(M_AXIS_BRAM_74_MB_DEPTH),
        .M_AXIS_BRAM_75_MB_DEPTH(M_AXIS_BRAM_75_MB_DEPTH),
        .M_AXIS_BRAM_76_MB_DEPTH(M_AXIS_BRAM_76_MB_DEPTH),
        .M_AXIS_BRAM_77_MB_DEPTH(M_AXIS_BRAM_77_MB_DEPTH),
        .M_AXIS_BRAM_78_MB_DEPTH(M_AXIS_BRAM_78_MB_DEPTH),
        .M_AXIS_BRAM_79_MB_DEPTH(M_AXIS_BRAM_79_MB_DEPTH),
        .M_AXIS_BRAM_80_MB_DEPTH(M_AXIS_BRAM_80_MB_DEPTH),
        .M_AXIS_BRAM_81_MB_DEPTH(M_AXIS_BRAM_81_MB_DEPTH),
        .M_AXIS_BRAM_82_MB_DEPTH(M_AXIS_BRAM_82_MB_DEPTH),
        .M_AXIS_BRAM_83_MB_DEPTH(M_AXIS_BRAM_83_MB_DEPTH),
        .M_AXIS_BRAM_84_MB_DEPTH(M_AXIS_BRAM_84_MB_DEPTH),
        .M_AXIS_BRAM_85_MB_DEPTH(M_AXIS_BRAM_85_MB_DEPTH),
        .M_AXIS_BRAM_86_MB_DEPTH(M_AXIS_BRAM_86_MB_DEPTH),
        .M_AXIS_BRAM_87_MB_DEPTH(M_AXIS_BRAM_87_MB_DEPTH),
        .M_AXIS_BRAM_88_MB_DEPTH(M_AXIS_BRAM_88_MB_DEPTH),
        .M_AXIS_BRAM_89_MB_DEPTH(M_AXIS_BRAM_89_MB_DEPTH),
        .M_AXIS_BRAM_90_MB_DEPTH(M_AXIS_BRAM_90_MB_DEPTH),
        .M_AXIS_BRAM_91_MB_DEPTH(M_AXIS_BRAM_91_MB_DEPTH),
        .M_AXIS_BRAM_92_MB_DEPTH(M_AXIS_BRAM_92_MB_DEPTH),
        .M_AXIS_BRAM_93_MB_DEPTH(M_AXIS_BRAM_93_MB_DEPTH),
        .M_AXIS_BRAM_94_MB_DEPTH(M_AXIS_BRAM_94_MB_DEPTH),
        .M_AXIS_BRAM_95_MB_DEPTH(M_AXIS_BRAM_95_MB_DEPTH),
        .M_AXIS_BRAM_96_MB_DEPTH(M_AXIS_BRAM_96_MB_DEPTH),
        .M_AXIS_BRAM_97_MB_DEPTH(M_AXIS_BRAM_97_MB_DEPTH),
        .M_AXIS_BRAM_98_MB_DEPTH(M_AXIS_BRAM_98_MB_DEPTH),
        .M_AXIS_BRAM_99_MB_DEPTH(M_AXIS_BRAM_99_MB_DEPTH),
        .M_AXIS_BRAM_100_MB_DEPTH(M_AXIS_BRAM_100_MB_DEPTH),
        .M_AXIS_BRAM_101_MB_DEPTH(M_AXIS_BRAM_101_MB_DEPTH),
        .M_AXIS_BRAM_102_MB_DEPTH(M_AXIS_BRAM_102_MB_DEPTH),
        .M_AXIS_BRAM_103_MB_DEPTH(M_AXIS_BRAM_103_MB_DEPTH),
        .M_AXIS_BRAM_104_MB_DEPTH(M_AXIS_BRAM_104_MB_DEPTH),
        .M_AXIS_BRAM_105_MB_DEPTH(M_AXIS_BRAM_105_MB_DEPTH),
        .M_AXIS_BRAM_106_MB_DEPTH(M_AXIS_BRAM_106_MB_DEPTH),
        .M_AXIS_BRAM_107_MB_DEPTH(M_AXIS_BRAM_107_MB_DEPTH),
        .M_AXIS_BRAM_108_MB_DEPTH(M_AXIS_BRAM_108_MB_DEPTH),
        .M_AXIS_BRAM_109_MB_DEPTH(M_AXIS_BRAM_109_MB_DEPTH),
        .M_AXIS_BRAM_110_MB_DEPTH(M_AXIS_BRAM_110_MB_DEPTH),
        .M_AXIS_BRAM_111_MB_DEPTH(M_AXIS_BRAM_111_MB_DEPTH),
        .M_AXIS_BRAM_112_MB_DEPTH(M_AXIS_BRAM_112_MB_DEPTH),
        .M_AXIS_BRAM_113_MB_DEPTH(M_AXIS_BRAM_113_MB_DEPTH),
        .M_AXIS_BRAM_114_MB_DEPTH(M_AXIS_BRAM_114_MB_DEPTH),
        .M_AXIS_BRAM_115_MB_DEPTH(M_AXIS_BRAM_115_MB_DEPTH),
        .M_AXIS_BRAM_116_MB_DEPTH(M_AXIS_BRAM_116_MB_DEPTH),
        .M_AXIS_BRAM_117_MB_DEPTH(M_AXIS_BRAM_117_MB_DEPTH),
        .M_AXIS_BRAM_118_MB_DEPTH(M_AXIS_BRAM_118_MB_DEPTH),
        .M_AXIS_BRAM_119_MB_DEPTH(M_AXIS_BRAM_119_MB_DEPTH),
        .M_AXIS_BRAM_120_MB_DEPTH(M_AXIS_BRAM_120_MB_DEPTH),
        .M_AXIS_BRAM_121_MB_DEPTH(M_AXIS_BRAM_121_MB_DEPTH),
        .M_AXIS_BRAM_122_MB_DEPTH(M_AXIS_BRAM_122_MB_DEPTH),
        .M_AXIS_BRAM_123_MB_DEPTH(M_AXIS_BRAM_123_MB_DEPTH),
        .M_AXIS_BRAM_124_MB_DEPTH(M_AXIS_BRAM_124_MB_DEPTH),
        .M_AXIS_BRAM_125_MB_DEPTH(M_AXIS_BRAM_125_MB_DEPTH),
        .M_AXIS_BRAM_126_MB_DEPTH(M_AXIS_BRAM_126_MB_DEPTH),
        .M_AXIS_BRAM_127_MB_DEPTH(M_AXIS_BRAM_127_MB_DEPTH),
        .M_AXIS_BRAM_0_ADDR_WIDTH(M_AXIS_BRAM_0_ADDR_WIDTH),
        .M_AXIS_BRAM_1_ADDR_WIDTH(M_AXIS_BRAM_1_ADDR_WIDTH),
        .M_AXIS_BRAM_2_ADDR_WIDTH(M_AXIS_BRAM_2_ADDR_WIDTH),
        .M_AXIS_BRAM_3_ADDR_WIDTH(M_AXIS_BRAM_3_ADDR_WIDTH),
        .M_AXIS_BRAM_4_ADDR_WIDTH(M_AXIS_BRAM_4_ADDR_WIDTH),
        .M_AXIS_BRAM_5_ADDR_WIDTH(M_AXIS_BRAM_5_ADDR_WIDTH),
        .M_AXIS_BRAM_6_ADDR_WIDTH(M_AXIS_BRAM_6_ADDR_WIDTH),
        .M_AXIS_BRAM_7_ADDR_WIDTH(M_AXIS_BRAM_7_ADDR_WIDTH),
        .M_AXIS_BRAM_8_ADDR_WIDTH(M_AXIS_BRAM_8_ADDR_WIDTH),
        .M_AXIS_BRAM_9_ADDR_WIDTH(M_AXIS_BRAM_9_ADDR_WIDTH),
        .M_AXIS_BRAM_10_ADDR_WIDTH(M_AXIS_BRAM_10_ADDR_WIDTH),
        .M_AXIS_BRAM_11_ADDR_WIDTH(M_AXIS_BRAM_11_ADDR_WIDTH),
        .M_AXIS_BRAM_12_ADDR_WIDTH(M_AXIS_BRAM_12_ADDR_WIDTH),
        .M_AXIS_BRAM_13_ADDR_WIDTH(M_AXIS_BRAM_13_ADDR_WIDTH),
        .M_AXIS_BRAM_14_ADDR_WIDTH(M_AXIS_BRAM_14_ADDR_WIDTH),
        .M_AXIS_BRAM_15_ADDR_WIDTH(M_AXIS_BRAM_15_ADDR_WIDTH),
        .M_AXIS_BRAM_16_ADDR_WIDTH(M_AXIS_BRAM_16_ADDR_WIDTH),
        .M_AXIS_BRAM_17_ADDR_WIDTH(M_AXIS_BRAM_17_ADDR_WIDTH),
        .M_AXIS_BRAM_18_ADDR_WIDTH(M_AXIS_BRAM_18_ADDR_WIDTH),
        .M_AXIS_BRAM_19_ADDR_WIDTH(M_AXIS_BRAM_19_ADDR_WIDTH),
        .M_AXIS_BRAM_20_ADDR_WIDTH(M_AXIS_BRAM_20_ADDR_WIDTH),
        .M_AXIS_BRAM_21_ADDR_WIDTH(M_AXIS_BRAM_21_ADDR_WIDTH),
        .M_AXIS_BRAM_22_ADDR_WIDTH(M_AXIS_BRAM_22_ADDR_WIDTH),
        .M_AXIS_BRAM_23_ADDR_WIDTH(M_AXIS_BRAM_23_ADDR_WIDTH),
        .M_AXIS_BRAM_24_ADDR_WIDTH(M_AXIS_BRAM_24_ADDR_WIDTH),
        .M_AXIS_BRAM_25_ADDR_WIDTH(M_AXIS_BRAM_25_ADDR_WIDTH),
        .M_AXIS_BRAM_26_ADDR_WIDTH(M_AXIS_BRAM_26_ADDR_WIDTH),
        .M_AXIS_BRAM_27_ADDR_WIDTH(M_AXIS_BRAM_27_ADDR_WIDTH),
        .M_AXIS_BRAM_28_ADDR_WIDTH(M_AXIS_BRAM_28_ADDR_WIDTH),
        .M_AXIS_BRAM_29_ADDR_WIDTH(M_AXIS_BRAM_29_ADDR_WIDTH),
        .M_AXIS_BRAM_30_ADDR_WIDTH(M_AXIS_BRAM_30_ADDR_WIDTH),
        .M_AXIS_BRAM_31_ADDR_WIDTH(M_AXIS_BRAM_31_ADDR_WIDTH),
        .M_AXIS_BRAM_32_ADDR_WIDTH(M_AXIS_BRAM_32_ADDR_WIDTH),
        .M_AXIS_BRAM_33_ADDR_WIDTH(M_AXIS_BRAM_33_ADDR_WIDTH),
        .M_AXIS_BRAM_34_ADDR_WIDTH(M_AXIS_BRAM_34_ADDR_WIDTH),
        .M_AXIS_BRAM_35_ADDR_WIDTH(M_AXIS_BRAM_35_ADDR_WIDTH),
        .M_AXIS_BRAM_36_ADDR_WIDTH(M_AXIS_BRAM_36_ADDR_WIDTH),
        .M_AXIS_BRAM_37_ADDR_WIDTH(M_AXIS_BRAM_37_ADDR_WIDTH),
        .M_AXIS_BRAM_38_ADDR_WIDTH(M_AXIS_BRAM_38_ADDR_WIDTH),
        .M_AXIS_BRAM_39_ADDR_WIDTH(M_AXIS_BRAM_39_ADDR_WIDTH),
        .M_AXIS_BRAM_40_ADDR_WIDTH(M_AXIS_BRAM_40_ADDR_WIDTH),
        .M_AXIS_BRAM_41_ADDR_WIDTH(M_AXIS_BRAM_41_ADDR_WIDTH),
        .M_AXIS_BRAM_42_ADDR_WIDTH(M_AXIS_BRAM_42_ADDR_WIDTH),
        .M_AXIS_BRAM_43_ADDR_WIDTH(M_AXIS_BRAM_43_ADDR_WIDTH),
        .M_AXIS_BRAM_44_ADDR_WIDTH(M_AXIS_BRAM_44_ADDR_WIDTH),
        .M_AXIS_BRAM_45_ADDR_WIDTH(M_AXIS_BRAM_45_ADDR_WIDTH),
        .M_AXIS_BRAM_46_ADDR_WIDTH(M_AXIS_BRAM_46_ADDR_WIDTH),
        .M_AXIS_BRAM_47_ADDR_WIDTH(M_AXIS_BRAM_47_ADDR_WIDTH),
        .M_AXIS_BRAM_48_ADDR_WIDTH(M_AXIS_BRAM_48_ADDR_WIDTH),
        .M_AXIS_BRAM_49_ADDR_WIDTH(M_AXIS_BRAM_49_ADDR_WIDTH),
        .M_AXIS_BRAM_50_ADDR_WIDTH(M_AXIS_BRAM_50_ADDR_WIDTH),
        .M_AXIS_BRAM_51_ADDR_WIDTH(M_AXIS_BRAM_51_ADDR_WIDTH),
        .M_AXIS_BRAM_52_ADDR_WIDTH(M_AXIS_BRAM_52_ADDR_WIDTH),
        .M_AXIS_BRAM_53_ADDR_WIDTH(M_AXIS_BRAM_53_ADDR_WIDTH),
        .M_AXIS_BRAM_54_ADDR_WIDTH(M_AXIS_BRAM_54_ADDR_WIDTH),
        .M_AXIS_BRAM_55_ADDR_WIDTH(M_AXIS_BRAM_55_ADDR_WIDTH),
        .M_AXIS_BRAM_56_ADDR_WIDTH(M_AXIS_BRAM_56_ADDR_WIDTH),
        .M_AXIS_BRAM_57_ADDR_WIDTH(M_AXIS_BRAM_57_ADDR_WIDTH),
        .M_AXIS_BRAM_58_ADDR_WIDTH(M_AXIS_BRAM_58_ADDR_WIDTH),
        .M_AXIS_BRAM_59_ADDR_WIDTH(M_AXIS_BRAM_59_ADDR_WIDTH),
        .M_AXIS_BRAM_60_ADDR_WIDTH(M_AXIS_BRAM_60_ADDR_WIDTH),
        .M_AXIS_BRAM_61_ADDR_WIDTH(M_AXIS_BRAM_61_ADDR_WIDTH),
        .M_AXIS_BRAM_62_ADDR_WIDTH(M_AXIS_BRAM_62_ADDR_WIDTH),
        .M_AXIS_BRAM_63_ADDR_WIDTH(M_AXIS_BRAM_63_ADDR_WIDTH),
        .M_AXIS_BRAM_64_ADDR_WIDTH(M_AXIS_BRAM_64_ADDR_WIDTH),
        .M_AXIS_BRAM_65_ADDR_WIDTH(M_AXIS_BRAM_65_ADDR_WIDTH),
        .M_AXIS_BRAM_66_ADDR_WIDTH(M_AXIS_BRAM_66_ADDR_WIDTH),
        .M_AXIS_BRAM_67_ADDR_WIDTH(M_AXIS_BRAM_67_ADDR_WIDTH),
        .M_AXIS_BRAM_68_ADDR_WIDTH(M_AXIS_BRAM_68_ADDR_WIDTH),
        .M_AXIS_BRAM_69_ADDR_WIDTH(M_AXIS_BRAM_69_ADDR_WIDTH),
        .M_AXIS_BRAM_70_ADDR_WIDTH(M_AXIS_BRAM_70_ADDR_WIDTH),
        .M_AXIS_BRAM_71_ADDR_WIDTH(M_AXIS_BRAM_71_ADDR_WIDTH),
        .M_AXIS_BRAM_72_ADDR_WIDTH(M_AXIS_BRAM_72_ADDR_WIDTH),
        .M_AXIS_BRAM_73_ADDR_WIDTH(M_AXIS_BRAM_73_ADDR_WIDTH),
        .M_AXIS_BRAM_74_ADDR_WIDTH(M_AXIS_BRAM_74_ADDR_WIDTH),
        .M_AXIS_BRAM_75_ADDR_WIDTH(M_AXIS_BRAM_75_ADDR_WIDTH),
        .M_AXIS_BRAM_76_ADDR_WIDTH(M_AXIS_BRAM_76_ADDR_WIDTH),
        .M_AXIS_BRAM_77_ADDR_WIDTH(M_AXIS_BRAM_77_ADDR_WIDTH),
        .M_AXIS_BRAM_78_ADDR_WIDTH(M_AXIS_BRAM_78_ADDR_WIDTH),
        .M_AXIS_BRAM_79_ADDR_WIDTH(M_AXIS_BRAM_79_ADDR_WIDTH),
        .M_AXIS_BRAM_80_ADDR_WIDTH(M_AXIS_BRAM_80_ADDR_WIDTH),
        .M_AXIS_BRAM_81_ADDR_WIDTH(M_AXIS_BRAM_81_ADDR_WIDTH),
        .M_AXIS_BRAM_82_ADDR_WIDTH(M_AXIS_BRAM_82_ADDR_WIDTH),
        .M_AXIS_BRAM_83_ADDR_WIDTH(M_AXIS_BRAM_83_ADDR_WIDTH),
        .M_AXIS_BRAM_84_ADDR_WIDTH(M_AXIS_BRAM_84_ADDR_WIDTH),
        .M_AXIS_BRAM_85_ADDR_WIDTH(M_AXIS_BRAM_85_ADDR_WIDTH),
        .M_AXIS_BRAM_86_ADDR_WIDTH(M_AXIS_BRAM_86_ADDR_WIDTH),
        .M_AXIS_BRAM_87_ADDR_WIDTH(M_AXIS_BRAM_87_ADDR_WIDTH),
        .M_AXIS_BRAM_88_ADDR_WIDTH(M_AXIS_BRAM_88_ADDR_WIDTH),
        .M_AXIS_BRAM_89_ADDR_WIDTH(M_AXIS_BRAM_89_ADDR_WIDTH),
        .M_AXIS_BRAM_90_ADDR_WIDTH(M_AXIS_BRAM_90_ADDR_WIDTH),
        .M_AXIS_BRAM_91_ADDR_WIDTH(M_AXIS_BRAM_91_ADDR_WIDTH),
        .M_AXIS_BRAM_92_ADDR_WIDTH(M_AXIS_BRAM_92_ADDR_WIDTH),
        .M_AXIS_BRAM_93_ADDR_WIDTH(M_AXIS_BRAM_93_ADDR_WIDTH),
        .M_AXIS_BRAM_94_ADDR_WIDTH(M_AXIS_BRAM_94_ADDR_WIDTH),
        .M_AXIS_BRAM_95_ADDR_WIDTH(M_AXIS_BRAM_95_ADDR_WIDTH),
        .M_AXIS_BRAM_96_ADDR_WIDTH(M_AXIS_BRAM_96_ADDR_WIDTH),
        .M_AXIS_BRAM_97_ADDR_WIDTH(M_AXIS_BRAM_97_ADDR_WIDTH),
        .M_AXIS_BRAM_98_ADDR_WIDTH(M_AXIS_BRAM_98_ADDR_WIDTH),
        .M_AXIS_BRAM_99_ADDR_WIDTH(M_AXIS_BRAM_99_ADDR_WIDTH),
        .M_AXIS_BRAM_100_ADDR_WIDTH(M_AXIS_BRAM_100_ADDR_WIDTH),
        .M_AXIS_BRAM_101_ADDR_WIDTH(M_AXIS_BRAM_101_ADDR_WIDTH),
        .M_AXIS_BRAM_102_ADDR_WIDTH(M_AXIS_BRAM_102_ADDR_WIDTH),
        .M_AXIS_BRAM_103_ADDR_WIDTH(M_AXIS_BRAM_103_ADDR_WIDTH),
        .M_AXIS_BRAM_104_ADDR_WIDTH(M_AXIS_BRAM_104_ADDR_WIDTH),
        .M_AXIS_BRAM_105_ADDR_WIDTH(M_AXIS_BRAM_105_ADDR_WIDTH),
        .M_AXIS_BRAM_106_ADDR_WIDTH(M_AXIS_BRAM_106_ADDR_WIDTH),
        .M_AXIS_BRAM_107_ADDR_WIDTH(M_AXIS_BRAM_107_ADDR_WIDTH),
        .M_AXIS_BRAM_108_ADDR_WIDTH(M_AXIS_BRAM_108_ADDR_WIDTH),
        .M_AXIS_BRAM_109_ADDR_WIDTH(M_AXIS_BRAM_109_ADDR_WIDTH),
        .M_AXIS_BRAM_110_ADDR_WIDTH(M_AXIS_BRAM_110_ADDR_WIDTH),
        .M_AXIS_BRAM_111_ADDR_WIDTH(M_AXIS_BRAM_111_ADDR_WIDTH),
        .M_AXIS_BRAM_112_ADDR_WIDTH(M_AXIS_BRAM_112_ADDR_WIDTH),
        .M_AXIS_BRAM_113_ADDR_WIDTH(M_AXIS_BRAM_113_ADDR_WIDTH),
        .M_AXIS_BRAM_114_ADDR_WIDTH(M_AXIS_BRAM_114_ADDR_WIDTH),
        .M_AXIS_BRAM_115_ADDR_WIDTH(M_AXIS_BRAM_115_ADDR_WIDTH),
        .M_AXIS_BRAM_116_ADDR_WIDTH(M_AXIS_BRAM_116_ADDR_WIDTH),
        .M_AXIS_BRAM_117_ADDR_WIDTH(M_AXIS_BRAM_117_ADDR_WIDTH),
        .M_AXIS_BRAM_118_ADDR_WIDTH(M_AXIS_BRAM_118_ADDR_WIDTH),
        .M_AXIS_BRAM_119_ADDR_WIDTH(M_AXIS_BRAM_119_ADDR_WIDTH),
        .M_AXIS_BRAM_120_ADDR_WIDTH(M_AXIS_BRAM_120_ADDR_WIDTH),
        .M_AXIS_BRAM_121_ADDR_WIDTH(M_AXIS_BRAM_121_ADDR_WIDTH),
        .M_AXIS_BRAM_122_ADDR_WIDTH(M_AXIS_BRAM_122_ADDR_WIDTH),
        .M_AXIS_BRAM_123_ADDR_WIDTH(M_AXIS_BRAM_123_ADDR_WIDTH),
        .M_AXIS_BRAM_124_ADDR_WIDTH(M_AXIS_BRAM_124_ADDR_WIDTH),
        .M_AXIS_BRAM_125_ADDR_WIDTH(M_AXIS_BRAM_125_ADDR_WIDTH),
        .M_AXIS_BRAM_126_ADDR_WIDTH(M_AXIS_BRAM_126_ADDR_WIDTH),
        .M_AXIS_BRAM_127_ADDR_WIDTH(M_AXIS_BRAM_127_ADDR_WIDTH)
    ) out_bram_args_i (
        .acc_clk(acc_aclk),
        .acc_aresetn(acc_aresetn),
        .dm_clk(s_axi_aclk),
        .dm_aresetn(s_axi_aresetn),
        .outbram_allow(outbram_ctrl_allow),
        .acc_start(ap_start_single),
        .acc_done(ap_done),
        .outbram_ready(outbram_ctrl_ready),
        .outbram_canstart(outbram_ctrl_canstart),
        .outbram_depth(outbram_depth),
        .outbram_depth_write(outbram_depth_write),
        .m_axis_bram_0_aclk(m_axis_bram_0_aclk),
        .m_axis_bram_0_aresetn(m_axis_bram_0_aresetn),
        .m_axis_bram_0_tlast(m_axis_bram_0_tlast),
        .m_axis_bram_0_tvalid(m_axis_bram_0_tvalid),
        .m_axis_bram_0_tkeep(m_axis_bram_0_tkeep),
        .m_axis_bram_0_tstrb(m_axis_bram_0_tstrb),
        .m_axis_bram_0_tdata(m_axis_bram_0_tdata),
        .m_axis_bram_0_tready(m_axis_bram_0_tready),
        .ap_bram_0_addr0(ap_bram_oarg_0_addr0),
        .ap_bram_0_din0(ap_bram_oarg_0_din0),
        .ap_bram_0_dout0(ap_bram_oarg_0_dout0),
        .ap_bram_0_we0(ap_bram_oarg_0_we0),
        .ap_bram_0_en0(ap_bram_oarg_0_en0),
        .ap_bram_0_addr1(ap_bram_oarg_0_addr1),
        .ap_bram_0_din1(ap_bram_oarg_0_din1),
        .ap_bram_0_dout1(ap_bram_oarg_0_dout1),
        .ap_bram_0_we1(ap_bram_oarg_0_we1),
        .ap_bram_0_en1(ap_bram_oarg_0_en1),
        .m_axis_bram_1_aclk(m_axis_bram_1_aclk),
        .m_axis_bram_1_aresetn(m_axis_bram_1_aresetn),
        .m_axis_bram_1_tlast(m_axis_bram_1_tlast),
        .m_axis_bram_1_tvalid(m_axis_bram_1_tvalid),
        .m_axis_bram_1_tkeep(m_axis_bram_1_tkeep),
        .m_axis_bram_1_tstrb(m_axis_bram_1_tstrb),
        .m_axis_bram_1_tdata(m_axis_bram_1_tdata),
        .m_axis_bram_1_tready(m_axis_bram_1_tready),
        .ap_bram_1_addr0(ap_bram_oarg_1_addr0),
        .ap_bram_1_din0(ap_bram_oarg_1_din0),
        .ap_bram_1_dout0(ap_bram_oarg_1_dout0),
        .ap_bram_1_we0(ap_bram_oarg_1_we0),
        .ap_bram_1_en0(ap_bram_oarg_1_en0),
        .ap_bram_1_addr1(ap_bram_oarg_1_addr1),
        .ap_bram_1_din1(ap_bram_oarg_1_din1),
        .ap_bram_1_dout1(ap_bram_oarg_1_dout1),
        .ap_bram_1_we1(ap_bram_oarg_1_we1),
        .ap_bram_1_en1(ap_bram_oarg_1_en1),
        .m_axis_bram_2_aclk(m_axis_bram_2_aclk),
        .m_axis_bram_2_aresetn(m_axis_bram_2_aresetn),
        .m_axis_bram_2_tlast(m_axis_bram_2_tlast),
        .m_axis_bram_2_tvalid(m_axis_bram_2_tvalid),
        .m_axis_bram_2_tkeep(m_axis_bram_2_tkeep),
        .m_axis_bram_2_tstrb(m_axis_bram_2_tstrb),
        .m_axis_bram_2_tdata(m_axis_bram_2_tdata),
        .m_axis_bram_2_tready(m_axis_bram_2_tready),
        .ap_bram_2_addr0(ap_bram_oarg_2_addr0),
        .ap_bram_2_din0(ap_bram_oarg_2_din0),
        .ap_bram_2_dout0(ap_bram_oarg_2_dout0),
        .ap_bram_2_we0(ap_bram_oarg_2_we0),
        .ap_bram_2_en0(ap_bram_oarg_2_en0),
        .ap_bram_2_addr1(ap_bram_oarg_2_addr1),
        .ap_bram_2_din1(ap_bram_oarg_2_din1),
        .ap_bram_2_dout1(ap_bram_oarg_2_dout1),
        .ap_bram_2_we1(ap_bram_oarg_2_we1),
        .ap_bram_2_en1(ap_bram_oarg_2_en1),
        .m_axis_bram_3_aclk(m_axis_bram_3_aclk),
        .m_axis_bram_3_aresetn(m_axis_bram_3_aresetn),
        .m_axis_bram_3_tlast(m_axis_bram_3_tlast),
        .m_axis_bram_3_tvalid(m_axis_bram_3_tvalid),
        .m_axis_bram_3_tkeep(m_axis_bram_3_tkeep),
        .m_axis_bram_3_tstrb(m_axis_bram_3_tstrb),
        .m_axis_bram_3_tdata(m_axis_bram_3_tdata),
        .m_axis_bram_3_tready(m_axis_bram_3_tready),
        .ap_bram_3_addr0(ap_bram_oarg_3_addr0),
        .ap_bram_3_din0(ap_bram_oarg_3_din0),
        .ap_bram_3_dout0(ap_bram_oarg_3_dout0),
        .ap_bram_3_we0(ap_bram_oarg_3_we0),
        .ap_bram_3_en0(ap_bram_oarg_3_en0),
        .ap_bram_3_addr1(ap_bram_oarg_3_addr1),
        .ap_bram_3_din1(ap_bram_oarg_3_din1),
        .ap_bram_3_dout1(ap_bram_oarg_3_dout1),
        .ap_bram_3_we1(ap_bram_oarg_3_we1),
        .ap_bram_3_en1(ap_bram_oarg_3_en1),
        .m_axis_bram_4_aclk(m_axis_bram_4_aclk),
        .m_axis_bram_4_aresetn(m_axis_bram_4_aresetn),
        .m_axis_bram_4_tlast(m_axis_bram_4_tlast),
        .m_axis_bram_4_tvalid(m_axis_bram_4_tvalid),
        .m_axis_bram_4_tkeep(m_axis_bram_4_tkeep),
        .m_axis_bram_4_tstrb(m_axis_bram_4_tstrb),
        .m_axis_bram_4_tdata(m_axis_bram_4_tdata),
        .m_axis_bram_4_tready(m_axis_bram_4_tready),
        .ap_bram_4_addr0(ap_bram_oarg_4_addr0),
        .ap_bram_4_din0(ap_bram_oarg_4_din0),
        .ap_bram_4_dout0(ap_bram_oarg_4_dout0),
        .ap_bram_4_we0(ap_bram_oarg_4_we0),
        .ap_bram_4_en0(ap_bram_oarg_4_en0),
        .ap_bram_4_addr1(ap_bram_oarg_4_addr1),
        .ap_bram_4_din1(ap_bram_oarg_4_din1),
        .ap_bram_4_dout1(ap_bram_oarg_4_dout1),
        .ap_bram_4_we1(ap_bram_oarg_4_we1),
        .ap_bram_4_en1(ap_bram_oarg_4_en1),
        .m_axis_bram_5_aclk(m_axis_bram_5_aclk),
        .m_axis_bram_5_aresetn(m_axis_bram_5_aresetn),
        .m_axis_bram_5_tlast(m_axis_bram_5_tlast),
        .m_axis_bram_5_tvalid(m_axis_bram_5_tvalid),
        .m_axis_bram_5_tkeep(m_axis_bram_5_tkeep),
        .m_axis_bram_5_tstrb(m_axis_bram_5_tstrb),
        .m_axis_bram_5_tdata(m_axis_bram_5_tdata),
        .m_axis_bram_5_tready(m_axis_bram_5_tready),
        .ap_bram_5_addr0(ap_bram_oarg_5_addr0),
        .ap_bram_5_din0(ap_bram_oarg_5_din0),
        .ap_bram_5_dout0(ap_bram_oarg_5_dout0),
        .ap_bram_5_we0(ap_bram_oarg_5_we0),
        .ap_bram_5_en0(ap_bram_oarg_5_en0),
        .ap_bram_5_addr1(ap_bram_oarg_5_addr1),
        .ap_bram_5_din1(ap_bram_oarg_5_din1),
        .ap_bram_5_dout1(ap_bram_oarg_5_dout1),
        .ap_bram_5_we1(ap_bram_oarg_5_we1),
        .ap_bram_5_en1(ap_bram_oarg_5_en1),
        .m_axis_bram_6_aclk(m_axis_bram_6_aclk),
        .m_axis_bram_6_aresetn(m_axis_bram_6_aresetn),
        .m_axis_bram_6_tlast(m_axis_bram_6_tlast),
        .m_axis_bram_6_tvalid(m_axis_bram_6_tvalid),
        .m_axis_bram_6_tkeep(m_axis_bram_6_tkeep),
        .m_axis_bram_6_tstrb(m_axis_bram_6_tstrb),
        .m_axis_bram_6_tdata(m_axis_bram_6_tdata),
        .m_axis_bram_6_tready(m_axis_bram_6_tready),
        .ap_bram_6_addr0(ap_bram_oarg_6_addr0),
        .ap_bram_6_din0(ap_bram_oarg_6_din0),
        .ap_bram_6_dout0(ap_bram_oarg_6_dout0),
        .ap_bram_6_we0(ap_bram_oarg_6_we0),
        .ap_bram_6_en0(ap_bram_oarg_6_en0),
        .ap_bram_6_addr1(ap_bram_oarg_6_addr1),
        .ap_bram_6_din1(ap_bram_oarg_6_din1),
        .ap_bram_6_dout1(ap_bram_oarg_6_dout1),
        .ap_bram_6_we1(ap_bram_oarg_6_we1),
        .ap_bram_6_en1(ap_bram_oarg_6_en1),
        .m_axis_bram_7_aclk(m_axis_bram_7_aclk),
        .m_axis_bram_7_aresetn(m_axis_bram_7_aresetn),
        .m_axis_bram_7_tlast(m_axis_bram_7_tlast),
        .m_axis_bram_7_tvalid(m_axis_bram_7_tvalid),
        .m_axis_bram_7_tkeep(m_axis_bram_7_tkeep),
        .m_axis_bram_7_tstrb(m_axis_bram_7_tstrb),
        .m_axis_bram_7_tdata(m_axis_bram_7_tdata),
        .m_axis_bram_7_tready(m_axis_bram_7_tready),
        .ap_bram_7_addr0(ap_bram_oarg_7_addr0),
        .ap_bram_7_din0(ap_bram_oarg_7_din0),
        .ap_bram_7_dout0(ap_bram_oarg_7_dout0),
        .ap_bram_7_we0(ap_bram_oarg_7_we0),
        .ap_bram_7_en0(ap_bram_oarg_7_en0),
        .ap_bram_7_addr1(ap_bram_oarg_7_addr1),
        .ap_bram_7_din1(ap_bram_oarg_7_din1),
        .ap_bram_7_dout1(ap_bram_oarg_7_dout1),
        .ap_bram_7_we1(ap_bram_oarg_7_we1),
        .ap_bram_7_en1(ap_bram_oarg_7_en1),
        .m_axis_bram_8_aclk(m_axis_bram_8_aclk),
        .m_axis_bram_8_aresetn(m_axis_bram_8_aresetn),
        .m_axis_bram_8_tlast(m_axis_bram_8_tlast),
        .m_axis_bram_8_tvalid(m_axis_bram_8_tvalid),
        .m_axis_bram_8_tkeep(m_axis_bram_8_tkeep),
        .m_axis_bram_8_tstrb(m_axis_bram_8_tstrb),
        .m_axis_bram_8_tdata(m_axis_bram_8_tdata),
        .m_axis_bram_8_tready(m_axis_bram_8_tready),
        .ap_bram_8_addr0(ap_bram_oarg_8_addr0),
        .ap_bram_8_din0(ap_bram_oarg_8_din0),
        .ap_bram_8_dout0(ap_bram_oarg_8_dout0),
        .ap_bram_8_we0(ap_bram_oarg_8_we0),
        .ap_bram_8_en0(ap_bram_oarg_8_en0),
        .ap_bram_8_addr1(ap_bram_oarg_8_addr1),
        .ap_bram_8_din1(ap_bram_oarg_8_din1),
        .ap_bram_8_dout1(ap_bram_oarg_8_dout1),
        .ap_bram_8_we1(ap_bram_oarg_8_we1),
        .ap_bram_8_en1(ap_bram_oarg_8_en1),
        .m_axis_bram_9_aclk(m_axis_bram_9_aclk),
        .m_axis_bram_9_aresetn(m_axis_bram_9_aresetn),
        .m_axis_bram_9_tlast(m_axis_bram_9_tlast),
        .m_axis_bram_9_tvalid(m_axis_bram_9_tvalid),
        .m_axis_bram_9_tkeep(m_axis_bram_9_tkeep),
        .m_axis_bram_9_tstrb(m_axis_bram_9_tstrb),
        .m_axis_bram_9_tdata(m_axis_bram_9_tdata),
        .m_axis_bram_9_tready(m_axis_bram_9_tready),
        .ap_bram_9_addr0(ap_bram_oarg_9_addr0),
        .ap_bram_9_din0(ap_bram_oarg_9_din0),
        .ap_bram_9_dout0(ap_bram_oarg_9_dout0),
        .ap_bram_9_we0(ap_bram_oarg_9_we0),
        .ap_bram_9_en0(ap_bram_oarg_9_en0),
        .ap_bram_9_addr1(ap_bram_oarg_9_addr1),
        .ap_bram_9_din1(ap_bram_oarg_9_din1),
        .ap_bram_9_dout1(ap_bram_oarg_9_dout1),
        .ap_bram_9_we1(ap_bram_oarg_9_we1),
        .ap_bram_9_en1(ap_bram_oarg_9_en1),
        .m_axis_bram_10_aclk(m_axis_bram_10_aclk),
        .m_axis_bram_10_aresetn(m_axis_bram_10_aresetn),
        .m_axis_bram_10_tlast(m_axis_bram_10_tlast),
        .m_axis_bram_10_tvalid(m_axis_bram_10_tvalid),
        .m_axis_bram_10_tkeep(m_axis_bram_10_tkeep),
        .m_axis_bram_10_tstrb(m_axis_bram_10_tstrb),
        .m_axis_bram_10_tdata(m_axis_bram_10_tdata),
        .m_axis_bram_10_tready(m_axis_bram_10_tready),
        .ap_bram_10_addr0(ap_bram_oarg_10_addr0),
        .ap_bram_10_din0(ap_bram_oarg_10_din0),
        .ap_bram_10_dout0(ap_bram_oarg_10_dout0),
        .ap_bram_10_we0(ap_bram_oarg_10_we0),
        .ap_bram_10_en0(ap_bram_oarg_10_en0),
        .ap_bram_10_addr1(ap_bram_oarg_10_addr1),
        .ap_bram_10_din1(ap_bram_oarg_10_din1),
        .ap_bram_10_dout1(ap_bram_oarg_10_dout1),
        .ap_bram_10_we1(ap_bram_oarg_10_we1),
        .ap_bram_10_en1(ap_bram_oarg_10_en1),
        .m_axis_bram_11_aclk(m_axis_bram_11_aclk),
        .m_axis_bram_11_aresetn(m_axis_bram_11_aresetn),
        .m_axis_bram_11_tlast(m_axis_bram_11_tlast),
        .m_axis_bram_11_tvalid(m_axis_bram_11_tvalid),
        .m_axis_bram_11_tkeep(m_axis_bram_11_tkeep),
        .m_axis_bram_11_tstrb(m_axis_bram_11_tstrb),
        .m_axis_bram_11_tdata(m_axis_bram_11_tdata),
        .m_axis_bram_11_tready(m_axis_bram_11_tready),
        .ap_bram_11_addr0(ap_bram_oarg_11_addr0),
        .ap_bram_11_din0(ap_bram_oarg_11_din0),
        .ap_bram_11_dout0(ap_bram_oarg_11_dout0),
        .ap_bram_11_we0(ap_bram_oarg_11_we0),
        .ap_bram_11_en0(ap_bram_oarg_11_en0),
        .ap_bram_11_addr1(ap_bram_oarg_11_addr1),
        .ap_bram_11_din1(ap_bram_oarg_11_din1),
        .ap_bram_11_dout1(ap_bram_oarg_11_dout1),
        .ap_bram_11_we1(ap_bram_oarg_11_we1),
        .ap_bram_11_en1(ap_bram_oarg_11_en1),
        .m_axis_bram_12_aclk(m_axis_bram_12_aclk),
        .m_axis_bram_12_aresetn(m_axis_bram_12_aresetn),
        .m_axis_bram_12_tlast(m_axis_bram_12_tlast),
        .m_axis_bram_12_tvalid(m_axis_bram_12_tvalid),
        .m_axis_bram_12_tkeep(m_axis_bram_12_tkeep),
        .m_axis_bram_12_tstrb(m_axis_bram_12_tstrb),
        .m_axis_bram_12_tdata(m_axis_bram_12_tdata),
        .m_axis_bram_12_tready(m_axis_bram_12_tready),
        .ap_bram_12_addr0(ap_bram_oarg_12_addr0),
        .ap_bram_12_din0(ap_bram_oarg_12_din0),
        .ap_bram_12_dout0(ap_bram_oarg_12_dout0),
        .ap_bram_12_we0(ap_bram_oarg_12_we0),
        .ap_bram_12_en0(ap_bram_oarg_12_en0),
        .ap_bram_12_addr1(ap_bram_oarg_12_addr1),
        .ap_bram_12_din1(ap_bram_oarg_12_din1),
        .ap_bram_12_dout1(ap_bram_oarg_12_dout1),
        .ap_bram_12_we1(ap_bram_oarg_12_we1),
        .ap_bram_12_en1(ap_bram_oarg_12_en1),
        .m_axis_bram_13_aclk(m_axis_bram_13_aclk),
        .m_axis_bram_13_aresetn(m_axis_bram_13_aresetn),
        .m_axis_bram_13_tlast(m_axis_bram_13_tlast),
        .m_axis_bram_13_tvalid(m_axis_bram_13_tvalid),
        .m_axis_bram_13_tkeep(m_axis_bram_13_tkeep),
        .m_axis_bram_13_tstrb(m_axis_bram_13_tstrb),
        .m_axis_bram_13_tdata(m_axis_bram_13_tdata),
        .m_axis_bram_13_tready(m_axis_bram_13_tready),
        .ap_bram_13_addr0(ap_bram_oarg_13_addr0),
        .ap_bram_13_din0(ap_bram_oarg_13_din0),
        .ap_bram_13_dout0(ap_bram_oarg_13_dout0),
        .ap_bram_13_we0(ap_bram_oarg_13_we0),
        .ap_bram_13_en0(ap_bram_oarg_13_en0),
        .ap_bram_13_addr1(ap_bram_oarg_13_addr1),
        .ap_bram_13_din1(ap_bram_oarg_13_din1),
        .ap_bram_13_dout1(ap_bram_oarg_13_dout1),
        .ap_bram_13_we1(ap_bram_oarg_13_we1),
        .ap_bram_13_en1(ap_bram_oarg_13_en1),
        .m_axis_bram_14_aclk(m_axis_bram_14_aclk),
        .m_axis_bram_14_aresetn(m_axis_bram_14_aresetn),
        .m_axis_bram_14_tlast(m_axis_bram_14_tlast),
        .m_axis_bram_14_tvalid(m_axis_bram_14_tvalid),
        .m_axis_bram_14_tkeep(m_axis_bram_14_tkeep),
        .m_axis_bram_14_tstrb(m_axis_bram_14_tstrb),
        .m_axis_bram_14_tdata(m_axis_bram_14_tdata),
        .m_axis_bram_14_tready(m_axis_bram_14_tready),
        .ap_bram_14_addr0(ap_bram_oarg_14_addr0),
        .ap_bram_14_din0(ap_bram_oarg_14_din0),
        .ap_bram_14_dout0(ap_bram_oarg_14_dout0),
        .ap_bram_14_we0(ap_bram_oarg_14_we0),
        .ap_bram_14_en0(ap_bram_oarg_14_en0),
        .ap_bram_14_addr1(ap_bram_oarg_14_addr1),
        .ap_bram_14_din1(ap_bram_oarg_14_din1),
        .ap_bram_14_dout1(ap_bram_oarg_14_dout1),
        .ap_bram_14_we1(ap_bram_oarg_14_we1),
        .ap_bram_14_en1(ap_bram_oarg_14_en1),
        .m_axis_bram_15_aclk(m_axis_bram_15_aclk),
        .m_axis_bram_15_aresetn(m_axis_bram_15_aresetn),
        .m_axis_bram_15_tlast(m_axis_bram_15_tlast),
        .m_axis_bram_15_tvalid(m_axis_bram_15_tvalid),
        .m_axis_bram_15_tkeep(m_axis_bram_15_tkeep),
        .m_axis_bram_15_tstrb(m_axis_bram_15_tstrb),
        .m_axis_bram_15_tdata(m_axis_bram_15_tdata),
        .m_axis_bram_15_tready(m_axis_bram_15_tready),
        .ap_bram_15_addr0(ap_bram_oarg_15_addr0),
        .ap_bram_15_din0(ap_bram_oarg_15_din0),
        .ap_bram_15_dout0(ap_bram_oarg_15_dout0),
        .ap_bram_15_we0(ap_bram_oarg_15_we0),
        .ap_bram_15_en0(ap_bram_oarg_15_en0),
        .ap_bram_15_addr1(ap_bram_oarg_15_addr1),
        .ap_bram_15_din1(ap_bram_oarg_15_din1),
        .ap_bram_15_dout1(ap_bram_oarg_15_dout1),
        .ap_bram_15_we1(ap_bram_oarg_15_we1),
        .ap_bram_15_en1(ap_bram_oarg_15_en1),
        .m_axis_bram_16_aclk(m_axis_bram_16_aclk),
        .m_axis_bram_16_aresetn(m_axis_bram_16_aresetn),
        .m_axis_bram_16_tlast(m_axis_bram_16_tlast),
        .m_axis_bram_16_tvalid(m_axis_bram_16_tvalid),
        .m_axis_bram_16_tkeep(m_axis_bram_16_tkeep),
        .m_axis_bram_16_tstrb(m_axis_bram_16_tstrb),
        .m_axis_bram_16_tdata(m_axis_bram_16_tdata),
        .m_axis_bram_16_tready(m_axis_bram_16_tready),
        .ap_bram_16_addr0(ap_bram_oarg_16_addr0),
        .ap_bram_16_din0(ap_bram_oarg_16_din0),
        .ap_bram_16_dout0(ap_bram_oarg_16_dout0),
        .ap_bram_16_we0(ap_bram_oarg_16_we0),
        .ap_bram_16_en0(ap_bram_oarg_16_en0),
        .ap_bram_16_addr1(ap_bram_oarg_16_addr1),
        .ap_bram_16_din1(ap_bram_oarg_16_din1),
        .ap_bram_16_dout1(ap_bram_oarg_16_dout1),
        .ap_bram_16_we1(ap_bram_oarg_16_we1),
        .ap_bram_16_en1(ap_bram_oarg_16_en1),
        .m_axis_bram_17_aclk(m_axis_bram_17_aclk),
        .m_axis_bram_17_aresetn(m_axis_bram_17_aresetn),
        .m_axis_bram_17_tlast(m_axis_bram_17_tlast),
        .m_axis_bram_17_tvalid(m_axis_bram_17_tvalid),
        .m_axis_bram_17_tkeep(m_axis_bram_17_tkeep),
        .m_axis_bram_17_tstrb(m_axis_bram_17_tstrb),
        .m_axis_bram_17_tdata(m_axis_bram_17_tdata),
        .m_axis_bram_17_tready(m_axis_bram_17_tready),
        .ap_bram_17_addr0(ap_bram_oarg_17_addr0),
        .ap_bram_17_din0(ap_bram_oarg_17_din0),
        .ap_bram_17_dout0(ap_bram_oarg_17_dout0),
        .ap_bram_17_we0(ap_bram_oarg_17_we0),
        .ap_bram_17_en0(ap_bram_oarg_17_en0),
        .ap_bram_17_addr1(ap_bram_oarg_17_addr1),
        .ap_bram_17_din1(ap_bram_oarg_17_din1),
        .ap_bram_17_dout1(ap_bram_oarg_17_dout1),
        .ap_bram_17_we1(ap_bram_oarg_17_we1),
        .ap_bram_17_en1(ap_bram_oarg_17_en1),
        .m_axis_bram_18_aclk(m_axis_bram_18_aclk),
        .m_axis_bram_18_aresetn(m_axis_bram_18_aresetn),
        .m_axis_bram_18_tlast(m_axis_bram_18_tlast),
        .m_axis_bram_18_tvalid(m_axis_bram_18_tvalid),
        .m_axis_bram_18_tkeep(m_axis_bram_18_tkeep),
        .m_axis_bram_18_tstrb(m_axis_bram_18_tstrb),
        .m_axis_bram_18_tdata(m_axis_bram_18_tdata),
        .m_axis_bram_18_tready(m_axis_bram_18_tready),
        .ap_bram_18_addr0(ap_bram_oarg_18_addr0),
        .ap_bram_18_din0(ap_bram_oarg_18_din0),
        .ap_bram_18_dout0(ap_bram_oarg_18_dout0),
        .ap_bram_18_we0(ap_bram_oarg_18_we0),
        .ap_bram_18_en0(ap_bram_oarg_18_en0),
        .ap_bram_18_addr1(ap_bram_oarg_18_addr1),
        .ap_bram_18_din1(ap_bram_oarg_18_din1),
        .ap_bram_18_dout1(ap_bram_oarg_18_dout1),
        .ap_bram_18_we1(ap_bram_oarg_18_we1),
        .ap_bram_18_en1(ap_bram_oarg_18_en1),
        .m_axis_bram_19_aclk(m_axis_bram_19_aclk),
        .m_axis_bram_19_aresetn(m_axis_bram_19_aresetn),
        .m_axis_bram_19_tlast(m_axis_bram_19_tlast),
        .m_axis_bram_19_tvalid(m_axis_bram_19_tvalid),
        .m_axis_bram_19_tkeep(m_axis_bram_19_tkeep),
        .m_axis_bram_19_tstrb(m_axis_bram_19_tstrb),
        .m_axis_bram_19_tdata(m_axis_bram_19_tdata),
        .m_axis_bram_19_tready(m_axis_bram_19_tready),
        .ap_bram_19_addr0(ap_bram_oarg_19_addr0),
        .ap_bram_19_din0(ap_bram_oarg_19_din0),
        .ap_bram_19_dout0(ap_bram_oarg_19_dout0),
        .ap_bram_19_we0(ap_bram_oarg_19_we0),
        .ap_bram_19_en0(ap_bram_oarg_19_en0),
        .ap_bram_19_addr1(ap_bram_oarg_19_addr1),
        .ap_bram_19_din1(ap_bram_oarg_19_din1),
        .ap_bram_19_dout1(ap_bram_oarg_19_dout1),
        .ap_bram_19_we1(ap_bram_oarg_19_we1),
        .ap_bram_19_en1(ap_bram_oarg_19_en1),
        .m_axis_bram_20_aclk(m_axis_bram_20_aclk),
        .m_axis_bram_20_aresetn(m_axis_bram_20_aresetn),
        .m_axis_bram_20_tlast(m_axis_bram_20_tlast),
        .m_axis_bram_20_tvalid(m_axis_bram_20_tvalid),
        .m_axis_bram_20_tkeep(m_axis_bram_20_tkeep),
        .m_axis_bram_20_tstrb(m_axis_bram_20_tstrb),
        .m_axis_bram_20_tdata(m_axis_bram_20_tdata),
        .m_axis_bram_20_tready(m_axis_bram_20_tready),
        .ap_bram_20_addr0(ap_bram_oarg_20_addr0),
        .ap_bram_20_din0(ap_bram_oarg_20_din0),
        .ap_bram_20_dout0(ap_bram_oarg_20_dout0),
        .ap_bram_20_we0(ap_bram_oarg_20_we0),
        .ap_bram_20_en0(ap_bram_oarg_20_en0),
        .ap_bram_20_addr1(ap_bram_oarg_20_addr1),
        .ap_bram_20_din1(ap_bram_oarg_20_din1),
        .ap_bram_20_dout1(ap_bram_oarg_20_dout1),
        .ap_bram_20_we1(ap_bram_oarg_20_we1),
        .ap_bram_20_en1(ap_bram_oarg_20_en1),
        .m_axis_bram_21_aclk(m_axis_bram_21_aclk),
        .m_axis_bram_21_aresetn(m_axis_bram_21_aresetn),
        .m_axis_bram_21_tlast(m_axis_bram_21_tlast),
        .m_axis_bram_21_tvalid(m_axis_bram_21_tvalid),
        .m_axis_bram_21_tkeep(m_axis_bram_21_tkeep),
        .m_axis_bram_21_tstrb(m_axis_bram_21_tstrb),
        .m_axis_bram_21_tdata(m_axis_bram_21_tdata),
        .m_axis_bram_21_tready(m_axis_bram_21_tready),
        .ap_bram_21_addr0(ap_bram_oarg_21_addr0),
        .ap_bram_21_din0(ap_bram_oarg_21_din0),
        .ap_bram_21_dout0(ap_bram_oarg_21_dout0),
        .ap_bram_21_we0(ap_bram_oarg_21_we0),
        .ap_bram_21_en0(ap_bram_oarg_21_en0),
        .ap_bram_21_addr1(ap_bram_oarg_21_addr1),
        .ap_bram_21_din1(ap_bram_oarg_21_din1),
        .ap_bram_21_dout1(ap_bram_oarg_21_dout1),
        .ap_bram_21_we1(ap_bram_oarg_21_we1),
        .ap_bram_21_en1(ap_bram_oarg_21_en1),
        .m_axis_bram_22_aclk(m_axis_bram_22_aclk),
        .m_axis_bram_22_aresetn(m_axis_bram_22_aresetn),
        .m_axis_bram_22_tlast(m_axis_bram_22_tlast),
        .m_axis_bram_22_tvalid(m_axis_bram_22_tvalid),
        .m_axis_bram_22_tkeep(m_axis_bram_22_tkeep),
        .m_axis_bram_22_tstrb(m_axis_bram_22_tstrb),
        .m_axis_bram_22_tdata(m_axis_bram_22_tdata),
        .m_axis_bram_22_tready(m_axis_bram_22_tready),
        .ap_bram_22_addr0(ap_bram_oarg_22_addr0),
        .ap_bram_22_din0(ap_bram_oarg_22_din0),
        .ap_bram_22_dout0(ap_bram_oarg_22_dout0),
        .ap_bram_22_we0(ap_bram_oarg_22_we0),
        .ap_bram_22_en0(ap_bram_oarg_22_en0),
        .ap_bram_22_addr1(ap_bram_oarg_22_addr1),
        .ap_bram_22_din1(ap_bram_oarg_22_din1),
        .ap_bram_22_dout1(ap_bram_oarg_22_dout1),
        .ap_bram_22_we1(ap_bram_oarg_22_we1),
        .ap_bram_22_en1(ap_bram_oarg_22_en1),
        .m_axis_bram_23_aclk(m_axis_bram_23_aclk),
        .m_axis_bram_23_aresetn(m_axis_bram_23_aresetn),
        .m_axis_bram_23_tlast(m_axis_bram_23_tlast),
        .m_axis_bram_23_tvalid(m_axis_bram_23_tvalid),
        .m_axis_bram_23_tkeep(m_axis_bram_23_tkeep),
        .m_axis_bram_23_tstrb(m_axis_bram_23_tstrb),
        .m_axis_bram_23_tdata(m_axis_bram_23_tdata),
        .m_axis_bram_23_tready(m_axis_bram_23_tready),
        .ap_bram_23_addr0(ap_bram_oarg_23_addr0),
        .ap_bram_23_din0(ap_bram_oarg_23_din0),
        .ap_bram_23_dout0(ap_bram_oarg_23_dout0),
        .ap_bram_23_we0(ap_bram_oarg_23_we0),
        .ap_bram_23_en0(ap_bram_oarg_23_en0),
        .ap_bram_23_addr1(ap_bram_oarg_23_addr1),
        .ap_bram_23_din1(ap_bram_oarg_23_din1),
        .ap_bram_23_dout1(ap_bram_oarg_23_dout1),
        .ap_bram_23_we1(ap_bram_oarg_23_we1),
        .ap_bram_23_en1(ap_bram_oarg_23_en1),
        .m_axis_bram_24_aclk(m_axis_bram_24_aclk),
        .m_axis_bram_24_aresetn(m_axis_bram_24_aresetn),
        .m_axis_bram_24_tlast(m_axis_bram_24_tlast),
        .m_axis_bram_24_tvalid(m_axis_bram_24_tvalid),
        .m_axis_bram_24_tkeep(m_axis_bram_24_tkeep),
        .m_axis_bram_24_tstrb(m_axis_bram_24_tstrb),
        .m_axis_bram_24_tdata(m_axis_bram_24_tdata),
        .m_axis_bram_24_tready(m_axis_bram_24_tready),
        .ap_bram_24_addr0(ap_bram_oarg_24_addr0),
        .ap_bram_24_din0(ap_bram_oarg_24_din0),
        .ap_bram_24_dout0(ap_bram_oarg_24_dout0),
        .ap_bram_24_we0(ap_bram_oarg_24_we0),
        .ap_bram_24_en0(ap_bram_oarg_24_en0),
        .ap_bram_24_addr1(ap_bram_oarg_24_addr1),
        .ap_bram_24_din1(ap_bram_oarg_24_din1),
        .ap_bram_24_dout1(ap_bram_oarg_24_dout1),
        .ap_bram_24_we1(ap_bram_oarg_24_we1),
        .ap_bram_24_en1(ap_bram_oarg_24_en1),
        .m_axis_bram_25_aclk(m_axis_bram_25_aclk),
        .m_axis_bram_25_aresetn(m_axis_bram_25_aresetn),
        .m_axis_bram_25_tlast(m_axis_bram_25_tlast),
        .m_axis_bram_25_tvalid(m_axis_bram_25_tvalid),
        .m_axis_bram_25_tkeep(m_axis_bram_25_tkeep),
        .m_axis_bram_25_tstrb(m_axis_bram_25_tstrb),
        .m_axis_bram_25_tdata(m_axis_bram_25_tdata),
        .m_axis_bram_25_tready(m_axis_bram_25_tready),
        .ap_bram_25_addr0(ap_bram_oarg_25_addr0),
        .ap_bram_25_din0(ap_bram_oarg_25_din0),
        .ap_bram_25_dout0(ap_bram_oarg_25_dout0),
        .ap_bram_25_we0(ap_bram_oarg_25_we0),
        .ap_bram_25_en0(ap_bram_oarg_25_en0),
        .ap_bram_25_addr1(ap_bram_oarg_25_addr1),
        .ap_bram_25_din1(ap_bram_oarg_25_din1),
        .ap_bram_25_dout1(ap_bram_oarg_25_dout1),
        .ap_bram_25_we1(ap_bram_oarg_25_we1),
        .ap_bram_25_en1(ap_bram_oarg_25_en1),
        .m_axis_bram_26_aclk(m_axis_bram_26_aclk),
        .m_axis_bram_26_aresetn(m_axis_bram_26_aresetn),
        .m_axis_bram_26_tlast(m_axis_bram_26_tlast),
        .m_axis_bram_26_tvalid(m_axis_bram_26_tvalid),
        .m_axis_bram_26_tkeep(m_axis_bram_26_tkeep),
        .m_axis_bram_26_tstrb(m_axis_bram_26_tstrb),
        .m_axis_bram_26_tdata(m_axis_bram_26_tdata),
        .m_axis_bram_26_tready(m_axis_bram_26_tready),
        .ap_bram_26_addr0(ap_bram_oarg_26_addr0),
        .ap_bram_26_din0(ap_bram_oarg_26_din0),
        .ap_bram_26_dout0(ap_bram_oarg_26_dout0),
        .ap_bram_26_we0(ap_bram_oarg_26_we0),
        .ap_bram_26_en0(ap_bram_oarg_26_en0),
        .ap_bram_26_addr1(ap_bram_oarg_26_addr1),
        .ap_bram_26_din1(ap_bram_oarg_26_din1),
        .ap_bram_26_dout1(ap_bram_oarg_26_dout1),
        .ap_bram_26_we1(ap_bram_oarg_26_we1),
        .ap_bram_26_en1(ap_bram_oarg_26_en1),
        .m_axis_bram_27_aclk(m_axis_bram_27_aclk),
        .m_axis_bram_27_aresetn(m_axis_bram_27_aresetn),
        .m_axis_bram_27_tlast(m_axis_bram_27_tlast),
        .m_axis_bram_27_tvalid(m_axis_bram_27_tvalid),
        .m_axis_bram_27_tkeep(m_axis_bram_27_tkeep),
        .m_axis_bram_27_tstrb(m_axis_bram_27_tstrb),
        .m_axis_bram_27_tdata(m_axis_bram_27_tdata),
        .m_axis_bram_27_tready(m_axis_bram_27_tready),
        .ap_bram_27_addr0(ap_bram_oarg_27_addr0),
        .ap_bram_27_din0(ap_bram_oarg_27_din0),
        .ap_bram_27_dout0(ap_bram_oarg_27_dout0),
        .ap_bram_27_we0(ap_bram_oarg_27_we0),
        .ap_bram_27_en0(ap_bram_oarg_27_en0),
        .ap_bram_27_addr1(ap_bram_oarg_27_addr1),
        .ap_bram_27_din1(ap_bram_oarg_27_din1),
        .ap_bram_27_dout1(ap_bram_oarg_27_dout1),
        .ap_bram_27_we1(ap_bram_oarg_27_we1),
        .ap_bram_27_en1(ap_bram_oarg_27_en1),
        .m_axis_bram_28_aclk(m_axis_bram_28_aclk),
        .m_axis_bram_28_aresetn(m_axis_bram_28_aresetn),
        .m_axis_bram_28_tlast(m_axis_bram_28_tlast),
        .m_axis_bram_28_tvalid(m_axis_bram_28_tvalid),
        .m_axis_bram_28_tkeep(m_axis_bram_28_tkeep),
        .m_axis_bram_28_tstrb(m_axis_bram_28_tstrb),
        .m_axis_bram_28_tdata(m_axis_bram_28_tdata),
        .m_axis_bram_28_tready(m_axis_bram_28_tready),
        .ap_bram_28_addr0(ap_bram_oarg_28_addr0),
        .ap_bram_28_din0(ap_bram_oarg_28_din0),
        .ap_bram_28_dout0(ap_bram_oarg_28_dout0),
        .ap_bram_28_we0(ap_bram_oarg_28_we0),
        .ap_bram_28_en0(ap_bram_oarg_28_en0),
        .ap_bram_28_addr1(ap_bram_oarg_28_addr1),
        .ap_bram_28_din1(ap_bram_oarg_28_din1),
        .ap_bram_28_dout1(ap_bram_oarg_28_dout1),
        .ap_bram_28_we1(ap_bram_oarg_28_we1),
        .ap_bram_28_en1(ap_bram_oarg_28_en1),
        .m_axis_bram_29_aclk(m_axis_bram_29_aclk),
        .m_axis_bram_29_aresetn(m_axis_bram_29_aresetn),
        .m_axis_bram_29_tlast(m_axis_bram_29_tlast),
        .m_axis_bram_29_tvalid(m_axis_bram_29_tvalid),
        .m_axis_bram_29_tkeep(m_axis_bram_29_tkeep),
        .m_axis_bram_29_tstrb(m_axis_bram_29_tstrb),
        .m_axis_bram_29_tdata(m_axis_bram_29_tdata),
        .m_axis_bram_29_tready(m_axis_bram_29_tready),
        .ap_bram_29_addr0(ap_bram_oarg_29_addr0),
        .ap_bram_29_din0(ap_bram_oarg_29_din0),
        .ap_bram_29_dout0(ap_bram_oarg_29_dout0),
        .ap_bram_29_we0(ap_bram_oarg_29_we0),
        .ap_bram_29_en0(ap_bram_oarg_29_en0),
        .ap_bram_29_addr1(ap_bram_oarg_29_addr1),
        .ap_bram_29_din1(ap_bram_oarg_29_din1),
        .ap_bram_29_dout1(ap_bram_oarg_29_dout1),
        .ap_bram_29_we1(ap_bram_oarg_29_we1),
        .ap_bram_29_en1(ap_bram_oarg_29_en1),
        .m_axis_bram_30_aclk(m_axis_bram_30_aclk),
        .m_axis_bram_30_aresetn(m_axis_bram_30_aresetn),
        .m_axis_bram_30_tlast(m_axis_bram_30_tlast),
        .m_axis_bram_30_tvalid(m_axis_bram_30_tvalid),
        .m_axis_bram_30_tkeep(m_axis_bram_30_tkeep),
        .m_axis_bram_30_tstrb(m_axis_bram_30_tstrb),
        .m_axis_bram_30_tdata(m_axis_bram_30_tdata),
        .m_axis_bram_30_tready(m_axis_bram_30_tready),
        .ap_bram_30_addr0(ap_bram_oarg_30_addr0),
        .ap_bram_30_din0(ap_bram_oarg_30_din0),
        .ap_bram_30_dout0(ap_bram_oarg_30_dout0),
        .ap_bram_30_we0(ap_bram_oarg_30_we0),
        .ap_bram_30_en0(ap_bram_oarg_30_en0),
        .ap_bram_30_addr1(ap_bram_oarg_30_addr1),
        .ap_bram_30_din1(ap_bram_oarg_30_din1),
        .ap_bram_30_dout1(ap_bram_oarg_30_dout1),
        .ap_bram_30_we1(ap_bram_oarg_30_we1),
        .ap_bram_30_en1(ap_bram_oarg_30_en1),
        .m_axis_bram_31_aclk(m_axis_bram_31_aclk),
        .m_axis_bram_31_aresetn(m_axis_bram_31_aresetn),
        .m_axis_bram_31_tlast(m_axis_bram_31_tlast),
        .m_axis_bram_31_tvalid(m_axis_bram_31_tvalid),
        .m_axis_bram_31_tkeep(m_axis_bram_31_tkeep),
        .m_axis_bram_31_tstrb(m_axis_bram_31_tstrb),
        .m_axis_bram_31_tdata(m_axis_bram_31_tdata),
        .m_axis_bram_31_tready(m_axis_bram_31_tready),
        .ap_bram_31_addr0(ap_bram_oarg_31_addr0),
        .ap_bram_31_din0(ap_bram_oarg_31_din0),
        .ap_bram_31_dout0(ap_bram_oarg_31_dout0),
        .ap_bram_31_we0(ap_bram_oarg_31_we0),
        .ap_bram_31_en0(ap_bram_oarg_31_en0),
        .ap_bram_31_addr1(ap_bram_oarg_31_addr1),
        .ap_bram_31_din1(ap_bram_oarg_31_din1),
        .ap_bram_31_dout1(ap_bram_oarg_31_dout1),
        .ap_bram_31_we1(ap_bram_oarg_31_we1),
        .ap_bram_31_en1(ap_bram_oarg_31_en1),
        .m_axis_bram_32_aclk(m_axis_bram_32_aclk),
        .m_axis_bram_32_aresetn(m_axis_bram_32_aresetn),
        .m_axis_bram_32_tlast(m_axis_bram_32_tlast),
        .m_axis_bram_32_tvalid(m_axis_bram_32_tvalid),
        .m_axis_bram_32_tkeep(m_axis_bram_32_tkeep),
        .m_axis_bram_32_tstrb(m_axis_bram_32_tstrb),
        .m_axis_bram_32_tdata(m_axis_bram_32_tdata),
        .m_axis_bram_32_tready(m_axis_bram_32_tready),
        .ap_bram_32_addr0(ap_bram_oarg_32_addr0),
        .ap_bram_32_din0(ap_bram_oarg_32_din0),
        .ap_bram_32_dout0(ap_bram_oarg_32_dout0),
        .ap_bram_32_we0(ap_bram_oarg_32_we0),
        .ap_bram_32_en0(ap_bram_oarg_32_en0),
        .ap_bram_32_addr1(ap_bram_oarg_32_addr1),
        .ap_bram_32_din1(ap_bram_oarg_32_din1),
        .ap_bram_32_dout1(ap_bram_oarg_32_dout1),
        .ap_bram_32_we1(ap_bram_oarg_32_we1),
        .ap_bram_32_en1(ap_bram_oarg_32_en1),
        .m_axis_bram_33_aclk(m_axis_bram_33_aclk),
        .m_axis_bram_33_aresetn(m_axis_bram_33_aresetn),
        .m_axis_bram_33_tlast(m_axis_bram_33_tlast),
        .m_axis_bram_33_tvalid(m_axis_bram_33_tvalid),
        .m_axis_bram_33_tkeep(m_axis_bram_33_tkeep),
        .m_axis_bram_33_tstrb(m_axis_bram_33_tstrb),
        .m_axis_bram_33_tdata(m_axis_bram_33_tdata),
        .m_axis_bram_33_tready(m_axis_bram_33_tready),
        .ap_bram_33_addr0(ap_bram_oarg_33_addr0),
        .ap_bram_33_din0(ap_bram_oarg_33_din0),
        .ap_bram_33_dout0(ap_bram_oarg_33_dout0),
        .ap_bram_33_we0(ap_bram_oarg_33_we0),
        .ap_bram_33_en0(ap_bram_oarg_33_en0),
        .ap_bram_33_addr1(ap_bram_oarg_33_addr1),
        .ap_bram_33_din1(ap_bram_oarg_33_din1),
        .ap_bram_33_dout1(ap_bram_oarg_33_dout1),
        .ap_bram_33_we1(ap_bram_oarg_33_we1),
        .ap_bram_33_en1(ap_bram_oarg_33_en1),
        .m_axis_bram_34_aclk(m_axis_bram_34_aclk),
        .m_axis_bram_34_aresetn(m_axis_bram_34_aresetn),
        .m_axis_bram_34_tlast(m_axis_bram_34_tlast),
        .m_axis_bram_34_tvalid(m_axis_bram_34_tvalid),
        .m_axis_bram_34_tkeep(m_axis_bram_34_tkeep),
        .m_axis_bram_34_tstrb(m_axis_bram_34_tstrb),
        .m_axis_bram_34_tdata(m_axis_bram_34_tdata),
        .m_axis_bram_34_tready(m_axis_bram_34_tready),
        .ap_bram_34_addr0(ap_bram_oarg_34_addr0),
        .ap_bram_34_din0(ap_bram_oarg_34_din0),
        .ap_bram_34_dout0(ap_bram_oarg_34_dout0),
        .ap_bram_34_we0(ap_bram_oarg_34_we0),
        .ap_bram_34_en0(ap_bram_oarg_34_en0),
        .ap_bram_34_addr1(ap_bram_oarg_34_addr1),
        .ap_bram_34_din1(ap_bram_oarg_34_din1),
        .ap_bram_34_dout1(ap_bram_oarg_34_dout1),
        .ap_bram_34_we1(ap_bram_oarg_34_we1),
        .ap_bram_34_en1(ap_bram_oarg_34_en1),
        .m_axis_bram_35_aclk(m_axis_bram_35_aclk),
        .m_axis_bram_35_aresetn(m_axis_bram_35_aresetn),
        .m_axis_bram_35_tlast(m_axis_bram_35_tlast),
        .m_axis_bram_35_tvalid(m_axis_bram_35_tvalid),
        .m_axis_bram_35_tkeep(m_axis_bram_35_tkeep),
        .m_axis_bram_35_tstrb(m_axis_bram_35_tstrb),
        .m_axis_bram_35_tdata(m_axis_bram_35_tdata),
        .m_axis_bram_35_tready(m_axis_bram_35_tready),
        .ap_bram_35_addr0(ap_bram_oarg_35_addr0),
        .ap_bram_35_din0(ap_bram_oarg_35_din0),
        .ap_bram_35_dout0(ap_bram_oarg_35_dout0),
        .ap_bram_35_we0(ap_bram_oarg_35_we0),
        .ap_bram_35_en0(ap_bram_oarg_35_en0),
        .ap_bram_35_addr1(ap_bram_oarg_35_addr1),
        .ap_bram_35_din1(ap_bram_oarg_35_din1),
        .ap_bram_35_dout1(ap_bram_oarg_35_dout1),
        .ap_bram_35_we1(ap_bram_oarg_35_we1),
        .ap_bram_35_en1(ap_bram_oarg_35_en1),
        .m_axis_bram_36_aclk(m_axis_bram_36_aclk),
        .m_axis_bram_36_aresetn(m_axis_bram_36_aresetn),
        .m_axis_bram_36_tlast(m_axis_bram_36_tlast),
        .m_axis_bram_36_tvalid(m_axis_bram_36_tvalid),
        .m_axis_bram_36_tkeep(m_axis_bram_36_tkeep),
        .m_axis_bram_36_tstrb(m_axis_bram_36_tstrb),
        .m_axis_bram_36_tdata(m_axis_bram_36_tdata),
        .m_axis_bram_36_tready(m_axis_bram_36_tready),
        .ap_bram_36_addr0(ap_bram_oarg_36_addr0),
        .ap_bram_36_din0(ap_bram_oarg_36_din0),
        .ap_bram_36_dout0(ap_bram_oarg_36_dout0),
        .ap_bram_36_we0(ap_bram_oarg_36_we0),
        .ap_bram_36_en0(ap_bram_oarg_36_en0),
        .ap_bram_36_addr1(ap_bram_oarg_36_addr1),
        .ap_bram_36_din1(ap_bram_oarg_36_din1),
        .ap_bram_36_dout1(ap_bram_oarg_36_dout1),
        .ap_bram_36_we1(ap_bram_oarg_36_we1),
        .ap_bram_36_en1(ap_bram_oarg_36_en1),
        .m_axis_bram_37_aclk(m_axis_bram_37_aclk),
        .m_axis_bram_37_aresetn(m_axis_bram_37_aresetn),
        .m_axis_bram_37_tlast(m_axis_bram_37_tlast),
        .m_axis_bram_37_tvalid(m_axis_bram_37_tvalid),
        .m_axis_bram_37_tkeep(m_axis_bram_37_tkeep),
        .m_axis_bram_37_tstrb(m_axis_bram_37_tstrb),
        .m_axis_bram_37_tdata(m_axis_bram_37_tdata),
        .m_axis_bram_37_tready(m_axis_bram_37_tready),
        .ap_bram_37_addr0(ap_bram_oarg_37_addr0),
        .ap_bram_37_din0(ap_bram_oarg_37_din0),
        .ap_bram_37_dout0(ap_bram_oarg_37_dout0),
        .ap_bram_37_we0(ap_bram_oarg_37_we0),
        .ap_bram_37_en0(ap_bram_oarg_37_en0),
        .ap_bram_37_addr1(ap_bram_oarg_37_addr1),
        .ap_bram_37_din1(ap_bram_oarg_37_din1),
        .ap_bram_37_dout1(ap_bram_oarg_37_dout1),
        .ap_bram_37_we1(ap_bram_oarg_37_we1),
        .ap_bram_37_en1(ap_bram_oarg_37_en1),
        .m_axis_bram_38_aclk(m_axis_bram_38_aclk),
        .m_axis_bram_38_aresetn(m_axis_bram_38_aresetn),
        .m_axis_bram_38_tlast(m_axis_bram_38_tlast),
        .m_axis_bram_38_tvalid(m_axis_bram_38_tvalid),
        .m_axis_bram_38_tkeep(m_axis_bram_38_tkeep),
        .m_axis_bram_38_tstrb(m_axis_bram_38_tstrb),
        .m_axis_bram_38_tdata(m_axis_bram_38_tdata),
        .m_axis_bram_38_tready(m_axis_bram_38_tready),
        .ap_bram_38_addr0(ap_bram_oarg_38_addr0),
        .ap_bram_38_din0(ap_bram_oarg_38_din0),
        .ap_bram_38_dout0(ap_bram_oarg_38_dout0),
        .ap_bram_38_we0(ap_bram_oarg_38_we0),
        .ap_bram_38_en0(ap_bram_oarg_38_en0),
        .ap_bram_38_addr1(ap_bram_oarg_38_addr1),
        .ap_bram_38_din1(ap_bram_oarg_38_din1),
        .ap_bram_38_dout1(ap_bram_oarg_38_dout1),
        .ap_bram_38_we1(ap_bram_oarg_38_we1),
        .ap_bram_38_en1(ap_bram_oarg_38_en1),
        .m_axis_bram_39_aclk(m_axis_bram_39_aclk),
        .m_axis_bram_39_aresetn(m_axis_bram_39_aresetn),
        .m_axis_bram_39_tlast(m_axis_bram_39_tlast),
        .m_axis_bram_39_tvalid(m_axis_bram_39_tvalid),
        .m_axis_bram_39_tkeep(m_axis_bram_39_tkeep),
        .m_axis_bram_39_tstrb(m_axis_bram_39_tstrb),
        .m_axis_bram_39_tdata(m_axis_bram_39_tdata),
        .m_axis_bram_39_tready(m_axis_bram_39_tready),
        .ap_bram_39_addr0(ap_bram_oarg_39_addr0),
        .ap_bram_39_din0(ap_bram_oarg_39_din0),
        .ap_bram_39_dout0(ap_bram_oarg_39_dout0),
        .ap_bram_39_we0(ap_bram_oarg_39_we0),
        .ap_bram_39_en0(ap_bram_oarg_39_en0),
        .ap_bram_39_addr1(ap_bram_oarg_39_addr1),
        .ap_bram_39_din1(ap_bram_oarg_39_din1),
        .ap_bram_39_dout1(ap_bram_oarg_39_dout1),
        .ap_bram_39_we1(ap_bram_oarg_39_we1),
        .ap_bram_39_en1(ap_bram_oarg_39_en1),
        .m_axis_bram_40_aclk(m_axis_bram_40_aclk),
        .m_axis_bram_40_aresetn(m_axis_bram_40_aresetn),
        .m_axis_bram_40_tlast(m_axis_bram_40_tlast),
        .m_axis_bram_40_tvalid(m_axis_bram_40_tvalid),
        .m_axis_bram_40_tkeep(m_axis_bram_40_tkeep),
        .m_axis_bram_40_tstrb(m_axis_bram_40_tstrb),
        .m_axis_bram_40_tdata(m_axis_bram_40_tdata),
        .m_axis_bram_40_tready(m_axis_bram_40_tready),
        .ap_bram_40_addr0(ap_bram_oarg_40_addr0),
        .ap_bram_40_din0(ap_bram_oarg_40_din0),
        .ap_bram_40_dout0(ap_bram_oarg_40_dout0),
        .ap_bram_40_we0(ap_bram_oarg_40_we0),
        .ap_bram_40_en0(ap_bram_oarg_40_en0),
        .ap_bram_40_addr1(ap_bram_oarg_40_addr1),
        .ap_bram_40_din1(ap_bram_oarg_40_din1),
        .ap_bram_40_dout1(ap_bram_oarg_40_dout1),
        .ap_bram_40_we1(ap_bram_oarg_40_we1),
        .ap_bram_40_en1(ap_bram_oarg_40_en1),
        .m_axis_bram_41_aclk(m_axis_bram_41_aclk),
        .m_axis_bram_41_aresetn(m_axis_bram_41_aresetn),
        .m_axis_bram_41_tlast(m_axis_bram_41_tlast),
        .m_axis_bram_41_tvalid(m_axis_bram_41_tvalid),
        .m_axis_bram_41_tkeep(m_axis_bram_41_tkeep),
        .m_axis_bram_41_tstrb(m_axis_bram_41_tstrb),
        .m_axis_bram_41_tdata(m_axis_bram_41_tdata),
        .m_axis_bram_41_tready(m_axis_bram_41_tready),
        .ap_bram_41_addr0(ap_bram_oarg_41_addr0),
        .ap_bram_41_din0(ap_bram_oarg_41_din0),
        .ap_bram_41_dout0(ap_bram_oarg_41_dout0),
        .ap_bram_41_we0(ap_bram_oarg_41_we0),
        .ap_bram_41_en0(ap_bram_oarg_41_en0),
        .ap_bram_41_addr1(ap_bram_oarg_41_addr1),
        .ap_bram_41_din1(ap_bram_oarg_41_din1),
        .ap_bram_41_dout1(ap_bram_oarg_41_dout1),
        .ap_bram_41_we1(ap_bram_oarg_41_we1),
        .ap_bram_41_en1(ap_bram_oarg_41_en1),
        .m_axis_bram_42_aclk(m_axis_bram_42_aclk),
        .m_axis_bram_42_aresetn(m_axis_bram_42_aresetn),
        .m_axis_bram_42_tlast(m_axis_bram_42_tlast),
        .m_axis_bram_42_tvalid(m_axis_bram_42_tvalid),
        .m_axis_bram_42_tkeep(m_axis_bram_42_tkeep),
        .m_axis_bram_42_tstrb(m_axis_bram_42_tstrb),
        .m_axis_bram_42_tdata(m_axis_bram_42_tdata),
        .m_axis_bram_42_tready(m_axis_bram_42_tready),
        .ap_bram_42_addr0(ap_bram_oarg_42_addr0),
        .ap_bram_42_din0(ap_bram_oarg_42_din0),
        .ap_bram_42_dout0(ap_bram_oarg_42_dout0),
        .ap_bram_42_we0(ap_bram_oarg_42_we0),
        .ap_bram_42_en0(ap_bram_oarg_42_en0),
        .ap_bram_42_addr1(ap_bram_oarg_42_addr1),
        .ap_bram_42_din1(ap_bram_oarg_42_din1),
        .ap_bram_42_dout1(ap_bram_oarg_42_dout1),
        .ap_bram_42_we1(ap_bram_oarg_42_we1),
        .ap_bram_42_en1(ap_bram_oarg_42_en1),
        .m_axis_bram_43_aclk(m_axis_bram_43_aclk),
        .m_axis_bram_43_aresetn(m_axis_bram_43_aresetn),
        .m_axis_bram_43_tlast(m_axis_bram_43_tlast),
        .m_axis_bram_43_tvalid(m_axis_bram_43_tvalid),
        .m_axis_bram_43_tkeep(m_axis_bram_43_tkeep),
        .m_axis_bram_43_tstrb(m_axis_bram_43_tstrb),
        .m_axis_bram_43_tdata(m_axis_bram_43_tdata),
        .m_axis_bram_43_tready(m_axis_bram_43_tready),
        .ap_bram_43_addr0(ap_bram_oarg_43_addr0),
        .ap_bram_43_din0(ap_bram_oarg_43_din0),
        .ap_bram_43_dout0(ap_bram_oarg_43_dout0),
        .ap_bram_43_we0(ap_bram_oarg_43_we0),
        .ap_bram_43_en0(ap_bram_oarg_43_en0),
        .ap_bram_43_addr1(ap_bram_oarg_43_addr1),
        .ap_bram_43_din1(ap_bram_oarg_43_din1),
        .ap_bram_43_dout1(ap_bram_oarg_43_dout1),
        .ap_bram_43_we1(ap_bram_oarg_43_we1),
        .ap_bram_43_en1(ap_bram_oarg_43_en1),
        .m_axis_bram_44_aclk(m_axis_bram_44_aclk),
        .m_axis_bram_44_aresetn(m_axis_bram_44_aresetn),
        .m_axis_bram_44_tlast(m_axis_bram_44_tlast),
        .m_axis_bram_44_tvalid(m_axis_bram_44_tvalid),
        .m_axis_bram_44_tkeep(m_axis_bram_44_tkeep),
        .m_axis_bram_44_tstrb(m_axis_bram_44_tstrb),
        .m_axis_bram_44_tdata(m_axis_bram_44_tdata),
        .m_axis_bram_44_tready(m_axis_bram_44_tready),
        .ap_bram_44_addr0(ap_bram_oarg_44_addr0),
        .ap_bram_44_din0(ap_bram_oarg_44_din0),
        .ap_bram_44_dout0(ap_bram_oarg_44_dout0),
        .ap_bram_44_we0(ap_bram_oarg_44_we0),
        .ap_bram_44_en0(ap_bram_oarg_44_en0),
        .ap_bram_44_addr1(ap_bram_oarg_44_addr1),
        .ap_bram_44_din1(ap_bram_oarg_44_din1),
        .ap_bram_44_dout1(ap_bram_oarg_44_dout1),
        .ap_bram_44_we1(ap_bram_oarg_44_we1),
        .ap_bram_44_en1(ap_bram_oarg_44_en1),
        .m_axis_bram_45_aclk(m_axis_bram_45_aclk),
        .m_axis_bram_45_aresetn(m_axis_bram_45_aresetn),
        .m_axis_bram_45_tlast(m_axis_bram_45_tlast),
        .m_axis_bram_45_tvalid(m_axis_bram_45_tvalid),
        .m_axis_bram_45_tkeep(m_axis_bram_45_tkeep),
        .m_axis_bram_45_tstrb(m_axis_bram_45_tstrb),
        .m_axis_bram_45_tdata(m_axis_bram_45_tdata),
        .m_axis_bram_45_tready(m_axis_bram_45_tready),
        .ap_bram_45_addr0(ap_bram_oarg_45_addr0),
        .ap_bram_45_din0(ap_bram_oarg_45_din0),
        .ap_bram_45_dout0(ap_bram_oarg_45_dout0),
        .ap_bram_45_we0(ap_bram_oarg_45_we0),
        .ap_bram_45_en0(ap_bram_oarg_45_en0),
        .ap_bram_45_addr1(ap_bram_oarg_45_addr1),
        .ap_bram_45_din1(ap_bram_oarg_45_din1),
        .ap_bram_45_dout1(ap_bram_oarg_45_dout1),
        .ap_bram_45_we1(ap_bram_oarg_45_we1),
        .ap_bram_45_en1(ap_bram_oarg_45_en1),
        .m_axis_bram_46_aclk(m_axis_bram_46_aclk),
        .m_axis_bram_46_aresetn(m_axis_bram_46_aresetn),
        .m_axis_bram_46_tlast(m_axis_bram_46_tlast),
        .m_axis_bram_46_tvalid(m_axis_bram_46_tvalid),
        .m_axis_bram_46_tkeep(m_axis_bram_46_tkeep),
        .m_axis_bram_46_tstrb(m_axis_bram_46_tstrb),
        .m_axis_bram_46_tdata(m_axis_bram_46_tdata),
        .m_axis_bram_46_tready(m_axis_bram_46_tready),
        .ap_bram_46_addr0(ap_bram_oarg_46_addr0),
        .ap_bram_46_din0(ap_bram_oarg_46_din0),
        .ap_bram_46_dout0(ap_bram_oarg_46_dout0),
        .ap_bram_46_we0(ap_bram_oarg_46_we0),
        .ap_bram_46_en0(ap_bram_oarg_46_en0),
        .ap_bram_46_addr1(ap_bram_oarg_46_addr1),
        .ap_bram_46_din1(ap_bram_oarg_46_din1),
        .ap_bram_46_dout1(ap_bram_oarg_46_dout1),
        .ap_bram_46_we1(ap_bram_oarg_46_we1),
        .ap_bram_46_en1(ap_bram_oarg_46_en1),
        .m_axis_bram_47_aclk(m_axis_bram_47_aclk),
        .m_axis_bram_47_aresetn(m_axis_bram_47_aresetn),
        .m_axis_bram_47_tlast(m_axis_bram_47_tlast),
        .m_axis_bram_47_tvalid(m_axis_bram_47_tvalid),
        .m_axis_bram_47_tkeep(m_axis_bram_47_tkeep),
        .m_axis_bram_47_tstrb(m_axis_bram_47_tstrb),
        .m_axis_bram_47_tdata(m_axis_bram_47_tdata),
        .m_axis_bram_47_tready(m_axis_bram_47_tready),
        .ap_bram_47_addr0(ap_bram_oarg_47_addr0),
        .ap_bram_47_din0(ap_bram_oarg_47_din0),
        .ap_bram_47_dout0(ap_bram_oarg_47_dout0),
        .ap_bram_47_we0(ap_bram_oarg_47_we0),
        .ap_bram_47_en0(ap_bram_oarg_47_en0),
        .ap_bram_47_addr1(ap_bram_oarg_47_addr1),
        .ap_bram_47_din1(ap_bram_oarg_47_din1),
        .ap_bram_47_dout1(ap_bram_oarg_47_dout1),
        .ap_bram_47_we1(ap_bram_oarg_47_we1),
        .ap_bram_47_en1(ap_bram_oarg_47_en1),
        .m_axis_bram_48_aclk(m_axis_bram_48_aclk),
        .m_axis_bram_48_aresetn(m_axis_bram_48_aresetn),
        .m_axis_bram_48_tlast(m_axis_bram_48_tlast),
        .m_axis_bram_48_tvalid(m_axis_bram_48_tvalid),
        .m_axis_bram_48_tkeep(m_axis_bram_48_tkeep),
        .m_axis_bram_48_tstrb(m_axis_bram_48_tstrb),
        .m_axis_bram_48_tdata(m_axis_bram_48_tdata),
        .m_axis_bram_48_tready(m_axis_bram_48_tready),
        .ap_bram_48_addr0(ap_bram_oarg_48_addr0),
        .ap_bram_48_din0(ap_bram_oarg_48_din0),
        .ap_bram_48_dout0(ap_bram_oarg_48_dout0),
        .ap_bram_48_we0(ap_bram_oarg_48_we0),
        .ap_bram_48_en0(ap_bram_oarg_48_en0),
        .ap_bram_48_addr1(ap_bram_oarg_48_addr1),
        .ap_bram_48_din1(ap_bram_oarg_48_din1),
        .ap_bram_48_dout1(ap_bram_oarg_48_dout1),
        .ap_bram_48_we1(ap_bram_oarg_48_we1),
        .ap_bram_48_en1(ap_bram_oarg_48_en1),
        .m_axis_bram_49_aclk(m_axis_bram_49_aclk),
        .m_axis_bram_49_aresetn(m_axis_bram_49_aresetn),
        .m_axis_bram_49_tlast(m_axis_bram_49_tlast),
        .m_axis_bram_49_tvalid(m_axis_bram_49_tvalid),
        .m_axis_bram_49_tkeep(m_axis_bram_49_tkeep),
        .m_axis_bram_49_tstrb(m_axis_bram_49_tstrb),
        .m_axis_bram_49_tdata(m_axis_bram_49_tdata),
        .m_axis_bram_49_tready(m_axis_bram_49_tready),
        .ap_bram_49_addr0(ap_bram_oarg_49_addr0),
        .ap_bram_49_din0(ap_bram_oarg_49_din0),
        .ap_bram_49_dout0(ap_bram_oarg_49_dout0),
        .ap_bram_49_we0(ap_bram_oarg_49_we0),
        .ap_bram_49_en0(ap_bram_oarg_49_en0),
        .ap_bram_49_addr1(ap_bram_oarg_49_addr1),
        .ap_bram_49_din1(ap_bram_oarg_49_din1),
        .ap_bram_49_dout1(ap_bram_oarg_49_dout1),
        .ap_bram_49_we1(ap_bram_oarg_49_we1),
        .ap_bram_49_en1(ap_bram_oarg_49_en1),
        .m_axis_bram_50_aclk(m_axis_bram_50_aclk),
        .m_axis_bram_50_aresetn(m_axis_bram_50_aresetn),
        .m_axis_bram_50_tlast(m_axis_bram_50_tlast),
        .m_axis_bram_50_tvalid(m_axis_bram_50_tvalid),
        .m_axis_bram_50_tkeep(m_axis_bram_50_tkeep),
        .m_axis_bram_50_tstrb(m_axis_bram_50_tstrb),
        .m_axis_bram_50_tdata(m_axis_bram_50_tdata),
        .m_axis_bram_50_tready(m_axis_bram_50_tready),
        .ap_bram_50_addr0(ap_bram_oarg_50_addr0),
        .ap_bram_50_din0(ap_bram_oarg_50_din0),
        .ap_bram_50_dout0(ap_bram_oarg_50_dout0),
        .ap_bram_50_we0(ap_bram_oarg_50_we0),
        .ap_bram_50_en0(ap_bram_oarg_50_en0),
        .ap_bram_50_addr1(ap_bram_oarg_50_addr1),
        .ap_bram_50_din1(ap_bram_oarg_50_din1),
        .ap_bram_50_dout1(ap_bram_oarg_50_dout1),
        .ap_bram_50_we1(ap_bram_oarg_50_we1),
        .ap_bram_50_en1(ap_bram_oarg_50_en1),
        .m_axis_bram_51_aclk(m_axis_bram_51_aclk),
        .m_axis_bram_51_aresetn(m_axis_bram_51_aresetn),
        .m_axis_bram_51_tlast(m_axis_bram_51_tlast),
        .m_axis_bram_51_tvalid(m_axis_bram_51_tvalid),
        .m_axis_bram_51_tkeep(m_axis_bram_51_tkeep),
        .m_axis_bram_51_tstrb(m_axis_bram_51_tstrb),
        .m_axis_bram_51_tdata(m_axis_bram_51_tdata),
        .m_axis_bram_51_tready(m_axis_bram_51_tready),
        .ap_bram_51_addr0(ap_bram_oarg_51_addr0),
        .ap_bram_51_din0(ap_bram_oarg_51_din0),
        .ap_bram_51_dout0(ap_bram_oarg_51_dout0),
        .ap_bram_51_we0(ap_bram_oarg_51_we0),
        .ap_bram_51_en0(ap_bram_oarg_51_en0),
        .ap_bram_51_addr1(ap_bram_oarg_51_addr1),
        .ap_bram_51_din1(ap_bram_oarg_51_din1),
        .ap_bram_51_dout1(ap_bram_oarg_51_dout1),
        .ap_bram_51_we1(ap_bram_oarg_51_we1),
        .ap_bram_51_en1(ap_bram_oarg_51_en1),
        .m_axis_bram_52_aclk(m_axis_bram_52_aclk),
        .m_axis_bram_52_aresetn(m_axis_bram_52_aresetn),
        .m_axis_bram_52_tlast(m_axis_bram_52_tlast),
        .m_axis_bram_52_tvalid(m_axis_bram_52_tvalid),
        .m_axis_bram_52_tkeep(m_axis_bram_52_tkeep),
        .m_axis_bram_52_tstrb(m_axis_bram_52_tstrb),
        .m_axis_bram_52_tdata(m_axis_bram_52_tdata),
        .m_axis_bram_52_tready(m_axis_bram_52_tready),
        .ap_bram_52_addr0(ap_bram_oarg_52_addr0),
        .ap_bram_52_din0(ap_bram_oarg_52_din0),
        .ap_bram_52_dout0(ap_bram_oarg_52_dout0),
        .ap_bram_52_we0(ap_bram_oarg_52_we0),
        .ap_bram_52_en0(ap_bram_oarg_52_en0),
        .ap_bram_52_addr1(ap_bram_oarg_52_addr1),
        .ap_bram_52_din1(ap_bram_oarg_52_din1),
        .ap_bram_52_dout1(ap_bram_oarg_52_dout1),
        .ap_bram_52_we1(ap_bram_oarg_52_we1),
        .ap_bram_52_en1(ap_bram_oarg_52_en1),
        .m_axis_bram_53_aclk(m_axis_bram_53_aclk),
        .m_axis_bram_53_aresetn(m_axis_bram_53_aresetn),
        .m_axis_bram_53_tlast(m_axis_bram_53_tlast),
        .m_axis_bram_53_tvalid(m_axis_bram_53_tvalid),
        .m_axis_bram_53_tkeep(m_axis_bram_53_tkeep),
        .m_axis_bram_53_tstrb(m_axis_bram_53_tstrb),
        .m_axis_bram_53_tdata(m_axis_bram_53_tdata),
        .m_axis_bram_53_tready(m_axis_bram_53_tready),
        .ap_bram_53_addr0(ap_bram_oarg_53_addr0),
        .ap_bram_53_din0(ap_bram_oarg_53_din0),
        .ap_bram_53_dout0(ap_bram_oarg_53_dout0),
        .ap_bram_53_we0(ap_bram_oarg_53_we0),
        .ap_bram_53_en0(ap_bram_oarg_53_en0),
        .ap_bram_53_addr1(ap_bram_oarg_53_addr1),
        .ap_bram_53_din1(ap_bram_oarg_53_din1),
        .ap_bram_53_dout1(ap_bram_oarg_53_dout1),
        .ap_bram_53_we1(ap_bram_oarg_53_we1),
        .ap_bram_53_en1(ap_bram_oarg_53_en1),
        .m_axis_bram_54_aclk(m_axis_bram_54_aclk),
        .m_axis_bram_54_aresetn(m_axis_bram_54_aresetn),
        .m_axis_bram_54_tlast(m_axis_bram_54_tlast),
        .m_axis_bram_54_tvalid(m_axis_bram_54_tvalid),
        .m_axis_bram_54_tkeep(m_axis_bram_54_tkeep),
        .m_axis_bram_54_tstrb(m_axis_bram_54_tstrb),
        .m_axis_bram_54_tdata(m_axis_bram_54_tdata),
        .m_axis_bram_54_tready(m_axis_bram_54_tready),
        .ap_bram_54_addr0(ap_bram_oarg_54_addr0),
        .ap_bram_54_din0(ap_bram_oarg_54_din0),
        .ap_bram_54_dout0(ap_bram_oarg_54_dout0),
        .ap_bram_54_we0(ap_bram_oarg_54_we0),
        .ap_bram_54_en0(ap_bram_oarg_54_en0),
        .ap_bram_54_addr1(ap_bram_oarg_54_addr1),
        .ap_bram_54_din1(ap_bram_oarg_54_din1),
        .ap_bram_54_dout1(ap_bram_oarg_54_dout1),
        .ap_bram_54_we1(ap_bram_oarg_54_we1),
        .ap_bram_54_en1(ap_bram_oarg_54_en1),
        .m_axis_bram_55_aclk(m_axis_bram_55_aclk),
        .m_axis_bram_55_aresetn(m_axis_bram_55_aresetn),
        .m_axis_bram_55_tlast(m_axis_bram_55_tlast),
        .m_axis_bram_55_tvalid(m_axis_bram_55_tvalid),
        .m_axis_bram_55_tkeep(m_axis_bram_55_tkeep),
        .m_axis_bram_55_tstrb(m_axis_bram_55_tstrb),
        .m_axis_bram_55_tdata(m_axis_bram_55_tdata),
        .m_axis_bram_55_tready(m_axis_bram_55_tready),
        .ap_bram_55_addr0(ap_bram_oarg_55_addr0),
        .ap_bram_55_din0(ap_bram_oarg_55_din0),
        .ap_bram_55_dout0(ap_bram_oarg_55_dout0),
        .ap_bram_55_we0(ap_bram_oarg_55_we0),
        .ap_bram_55_en0(ap_bram_oarg_55_en0),
        .ap_bram_55_addr1(ap_bram_oarg_55_addr1),
        .ap_bram_55_din1(ap_bram_oarg_55_din1),
        .ap_bram_55_dout1(ap_bram_oarg_55_dout1),
        .ap_bram_55_we1(ap_bram_oarg_55_we1),
        .ap_bram_55_en1(ap_bram_oarg_55_en1),
        .m_axis_bram_56_aclk(m_axis_bram_56_aclk),
        .m_axis_bram_56_aresetn(m_axis_bram_56_aresetn),
        .m_axis_bram_56_tlast(m_axis_bram_56_tlast),
        .m_axis_bram_56_tvalid(m_axis_bram_56_tvalid),
        .m_axis_bram_56_tkeep(m_axis_bram_56_tkeep),
        .m_axis_bram_56_tstrb(m_axis_bram_56_tstrb),
        .m_axis_bram_56_tdata(m_axis_bram_56_tdata),
        .m_axis_bram_56_tready(m_axis_bram_56_tready),
        .ap_bram_56_addr0(ap_bram_oarg_56_addr0),
        .ap_bram_56_din0(ap_bram_oarg_56_din0),
        .ap_bram_56_dout0(ap_bram_oarg_56_dout0),
        .ap_bram_56_we0(ap_bram_oarg_56_we0),
        .ap_bram_56_en0(ap_bram_oarg_56_en0),
        .ap_bram_56_addr1(ap_bram_oarg_56_addr1),
        .ap_bram_56_din1(ap_bram_oarg_56_din1),
        .ap_bram_56_dout1(ap_bram_oarg_56_dout1),
        .ap_bram_56_we1(ap_bram_oarg_56_we1),
        .ap_bram_56_en1(ap_bram_oarg_56_en1),
        .m_axis_bram_57_aclk(m_axis_bram_57_aclk),
        .m_axis_bram_57_aresetn(m_axis_bram_57_aresetn),
        .m_axis_bram_57_tlast(m_axis_bram_57_tlast),
        .m_axis_bram_57_tvalid(m_axis_bram_57_tvalid),
        .m_axis_bram_57_tkeep(m_axis_bram_57_tkeep),
        .m_axis_bram_57_tstrb(m_axis_bram_57_tstrb),
        .m_axis_bram_57_tdata(m_axis_bram_57_tdata),
        .m_axis_bram_57_tready(m_axis_bram_57_tready),
        .ap_bram_57_addr0(ap_bram_oarg_57_addr0),
        .ap_bram_57_din0(ap_bram_oarg_57_din0),
        .ap_bram_57_dout0(ap_bram_oarg_57_dout0),
        .ap_bram_57_we0(ap_bram_oarg_57_we0),
        .ap_bram_57_en0(ap_bram_oarg_57_en0),
        .ap_bram_57_addr1(ap_bram_oarg_57_addr1),
        .ap_bram_57_din1(ap_bram_oarg_57_din1),
        .ap_bram_57_dout1(ap_bram_oarg_57_dout1),
        .ap_bram_57_we1(ap_bram_oarg_57_we1),
        .ap_bram_57_en1(ap_bram_oarg_57_en1),
        .m_axis_bram_58_aclk(m_axis_bram_58_aclk),
        .m_axis_bram_58_aresetn(m_axis_bram_58_aresetn),
        .m_axis_bram_58_tlast(m_axis_bram_58_tlast),
        .m_axis_bram_58_tvalid(m_axis_bram_58_tvalid),
        .m_axis_bram_58_tkeep(m_axis_bram_58_tkeep),
        .m_axis_bram_58_tstrb(m_axis_bram_58_tstrb),
        .m_axis_bram_58_tdata(m_axis_bram_58_tdata),
        .m_axis_bram_58_tready(m_axis_bram_58_tready),
        .ap_bram_58_addr0(ap_bram_oarg_58_addr0),
        .ap_bram_58_din0(ap_bram_oarg_58_din0),
        .ap_bram_58_dout0(ap_bram_oarg_58_dout0),
        .ap_bram_58_we0(ap_bram_oarg_58_we0),
        .ap_bram_58_en0(ap_bram_oarg_58_en0),
        .ap_bram_58_addr1(ap_bram_oarg_58_addr1),
        .ap_bram_58_din1(ap_bram_oarg_58_din1),
        .ap_bram_58_dout1(ap_bram_oarg_58_dout1),
        .ap_bram_58_we1(ap_bram_oarg_58_we1),
        .ap_bram_58_en1(ap_bram_oarg_58_en1),
        .m_axis_bram_59_aclk(m_axis_bram_59_aclk),
        .m_axis_bram_59_aresetn(m_axis_bram_59_aresetn),
        .m_axis_bram_59_tlast(m_axis_bram_59_tlast),
        .m_axis_bram_59_tvalid(m_axis_bram_59_tvalid),
        .m_axis_bram_59_tkeep(m_axis_bram_59_tkeep),
        .m_axis_bram_59_tstrb(m_axis_bram_59_tstrb),
        .m_axis_bram_59_tdata(m_axis_bram_59_tdata),
        .m_axis_bram_59_tready(m_axis_bram_59_tready),
        .ap_bram_59_addr0(ap_bram_oarg_59_addr0),
        .ap_bram_59_din0(ap_bram_oarg_59_din0),
        .ap_bram_59_dout0(ap_bram_oarg_59_dout0),
        .ap_bram_59_we0(ap_bram_oarg_59_we0),
        .ap_bram_59_en0(ap_bram_oarg_59_en0),
        .ap_bram_59_addr1(ap_bram_oarg_59_addr1),
        .ap_bram_59_din1(ap_bram_oarg_59_din1),
        .ap_bram_59_dout1(ap_bram_oarg_59_dout1),
        .ap_bram_59_we1(ap_bram_oarg_59_we1),
        .ap_bram_59_en1(ap_bram_oarg_59_en1),
        .m_axis_bram_60_aclk(m_axis_bram_60_aclk),
        .m_axis_bram_60_aresetn(m_axis_bram_60_aresetn),
        .m_axis_bram_60_tlast(m_axis_bram_60_tlast),
        .m_axis_bram_60_tvalid(m_axis_bram_60_tvalid),
        .m_axis_bram_60_tkeep(m_axis_bram_60_tkeep),
        .m_axis_bram_60_tstrb(m_axis_bram_60_tstrb),
        .m_axis_bram_60_tdata(m_axis_bram_60_tdata),
        .m_axis_bram_60_tready(m_axis_bram_60_tready),
        .ap_bram_60_addr0(ap_bram_oarg_60_addr0),
        .ap_bram_60_din0(ap_bram_oarg_60_din0),
        .ap_bram_60_dout0(ap_bram_oarg_60_dout0),
        .ap_bram_60_we0(ap_bram_oarg_60_we0),
        .ap_bram_60_en0(ap_bram_oarg_60_en0),
        .ap_bram_60_addr1(ap_bram_oarg_60_addr1),
        .ap_bram_60_din1(ap_bram_oarg_60_din1),
        .ap_bram_60_dout1(ap_bram_oarg_60_dout1),
        .ap_bram_60_we1(ap_bram_oarg_60_we1),
        .ap_bram_60_en1(ap_bram_oarg_60_en1),
        .m_axis_bram_61_aclk(m_axis_bram_61_aclk),
        .m_axis_bram_61_aresetn(m_axis_bram_61_aresetn),
        .m_axis_bram_61_tlast(m_axis_bram_61_tlast),
        .m_axis_bram_61_tvalid(m_axis_bram_61_tvalid),
        .m_axis_bram_61_tkeep(m_axis_bram_61_tkeep),
        .m_axis_bram_61_tstrb(m_axis_bram_61_tstrb),
        .m_axis_bram_61_tdata(m_axis_bram_61_tdata),
        .m_axis_bram_61_tready(m_axis_bram_61_tready),
        .ap_bram_61_addr0(ap_bram_oarg_61_addr0),
        .ap_bram_61_din0(ap_bram_oarg_61_din0),
        .ap_bram_61_dout0(ap_bram_oarg_61_dout0),
        .ap_bram_61_we0(ap_bram_oarg_61_we0),
        .ap_bram_61_en0(ap_bram_oarg_61_en0),
        .ap_bram_61_addr1(ap_bram_oarg_61_addr1),
        .ap_bram_61_din1(ap_bram_oarg_61_din1),
        .ap_bram_61_dout1(ap_bram_oarg_61_dout1),
        .ap_bram_61_we1(ap_bram_oarg_61_we1),
        .ap_bram_61_en1(ap_bram_oarg_61_en1),
        .m_axis_bram_62_aclk(m_axis_bram_62_aclk),
        .m_axis_bram_62_aresetn(m_axis_bram_62_aresetn),
        .m_axis_bram_62_tlast(m_axis_bram_62_tlast),
        .m_axis_bram_62_tvalid(m_axis_bram_62_tvalid),
        .m_axis_bram_62_tkeep(m_axis_bram_62_tkeep),
        .m_axis_bram_62_tstrb(m_axis_bram_62_tstrb),
        .m_axis_bram_62_tdata(m_axis_bram_62_tdata),
        .m_axis_bram_62_tready(m_axis_bram_62_tready),
        .ap_bram_62_addr0(ap_bram_oarg_62_addr0),
        .ap_bram_62_din0(ap_bram_oarg_62_din0),
        .ap_bram_62_dout0(ap_bram_oarg_62_dout0),
        .ap_bram_62_we0(ap_bram_oarg_62_we0),
        .ap_bram_62_en0(ap_bram_oarg_62_en0),
        .ap_bram_62_addr1(ap_bram_oarg_62_addr1),
        .ap_bram_62_din1(ap_bram_oarg_62_din1),
        .ap_bram_62_dout1(ap_bram_oarg_62_dout1),
        .ap_bram_62_we1(ap_bram_oarg_62_we1),
        .ap_bram_62_en1(ap_bram_oarg_62_en1),
        .m_axis_bram_63_aclk(m_axis_bram_63_aclk),
        .m_axis_bram_63_aresetn(m_axis_bram_63_aresetn),
        .m_axis_bram_63_tlast(m_axis_bram_63_tlast),
        .m_axis_bram_63_tvalid(m_axis_bram_63_tvalid),
        .m_axis_bram_63_tkeep(m_axis_bram_63_tkeep),
        .m_axis_bram_63_tstrb(m_axis_bram_63_tstrb),
        .m_axis_bram_63_tdata(m_axis_bram_63_tdata),
        .m_axis_bram_63_tready(m_axis_bram_63_tready),
        .ap_bram_63_addr0(ap_bram_oarg_63_addr0),
        .ap_bram_63_din0(ap_bram_oarg_63_din0),
        .ap_bram_63_dout0(ap_bram_oarg_63_dout0),
        .ap_bram_63_we0(ap_bram_oarg_63_we0),
        .ap_bram_63_en0(ap_bram_oarg_63_en0),
        .ap_bram_63_addr1(ap_bram_oarg_63_addr1),
        .ap_bram_63_din1(ap_bram_oarg_63_din1),
        .ap_bram_63_dout1(ap_bram_oarg_63_dout1),
        .ap_bram_63_we1(ap_bram_oarg_63_we1),
        .ap_bram_63_en1(ap_bram_oarg_63_en1),
        .m_axis_bram_64_aclk(m_axis_bram_64_aclk),
        .m_axis_bram_64_aresetn(m_axis_bram_64_aresetn),
        .m_axis_bram_64_tlast(m_axis_bram_64_tlast),
        .m_axis_bram_64_tvalid(m_axis_bram_64_tvalid),
        .m_axis_bram_64_tkeep(m_axis_bram_64_tkeep),
        .m_axis_bram_64_tstrb(m_axis_bram_64_tstrb),
        .m_axis_bram_64_tdata(m_axis_bram_64_tdata),
        .m_axis_bram_64_tready(m_axis_bram_64_tready),
        .ap_bram_64_addr0(ap_bram_oarg_64_addr0),
        .ap_bram_64_din0(ap_bram_oarg_64_din0),
        .ap_bram_64_dout0(ap_bram_oarg_64_dout0),
        .ap_bram_64_we0(ap_bram_oarg_64_we0),
        .ap_bram_64_en0(ap_bram_oarg_64_en0),
        .ap_bram_64_addr1(ap_bram_oarg_64_addr1),
        .ap_bram_64_din1(ap_bram_oarg_64_din1),
        .ap_bram_64_dout1(ap_bram_oarg_64_dout1),
        .ap_bram_64_we1(ap_bram_oarg_64_we1),
        .ap_bram_64_en1(ap_bram_oarg_64_en1),
        .m_axis_bram_65_aclk(m_axis_bram_65_aclk),
        .m_axis_bram_65_aresetn(m_axis_bram_65_aresetn),
        .m_axis_bram_65_tlast(m_axis_bram_65_tlast),
        .m_axis_bram_65_tvalid(m_axis_bram_65_tvalid),
        .m_axis_bram_65_tkeep(m_axis_bram_65_tkeep),
        .m_axis_bram_65_tstrb(m_axis_bram_65_tstrb),
        .m_axis_bram_65_tdata(m_axis_bram_65_tdata),
        .m_axis_bram_65_tready(m_axis_bram_65_tready),
        .ap_bram_65_addr0(ap_bram_oarg_65_addr0),
        .ap_bram_65_din0(ap_bram_oarg_65_din0),
        .ap_bram_65_dout0(ap_bram_oarg_65_dout0),
        .ap_bram_65_we0(ap_bram_oarg_65_we0),
        .ap_bram_65_en0(ap_bram_oarg_65_en0),
        .ap_bram_65_addr1(ap_bram_oarg_65_addr1),
        .ap_bram_65_din1(ap_bram_oarg_65_din1),
        .ap_bram_65_dout1(ap_bram_oarg_65_dout1),
        .ap_bram_65_we1(ap_bram_oarg_65_we1),
        .ap_bram_65_en1(ap_bram_oarg_65_en1),
        .m_axis_bram_66_aclk(m_axis_bram_66_aclk),
        .m_axis_bram_66_aresetn(m_axis_bram_66_aresetn),
        .m_axis_bram_66_tlast(m_axis_bram_66_tlast),
        .m_axis_bram_66_tvalid(m_axis_bram_66_tvalid),
        .m_axis_bram_66_tkeep(m_axis_bram_66_tkeep),
        .m_axis_bram_66_tstrb(m_axis_bram_66_tstrb),
        .m_axis_bram_66_tdata(m_axis_bram_66_tdata),
        .m_axis_bram_66_tready(m_axis_bram_66_tready),
        .ap_bram_66_addr0(ap_bram_oarg_66_addr0),
        .ap_bram_66_din0(ap_bram_oarg_66_din0),
        .ap_bram_66_dout0(ap_bram_oarg_66_dout0),
        .ap_bram_66_we0(ap_bram_oarg_66_we0),
        .ap_bram_66_en0(ap_bram_oarg_66_en0),
        .ap_bram_66_addr1(ap_bram_oarg_66_addr1),
        .ap_bram_66_din1(ap_bram_oarg_66_din1),
        .ap_bram_66_dout1(ap_bram_oarg_66_dout1),
        .ap_bram_66_we1(ap_bram_oarg_66_we1),
        .ap_bram_66_en1(ap_bram_oarg_66_en1),
        .m_axis_bram_67_aclk(m_axis_bram_67_aclk),
        .m_axis_bram_67_aresetn(m_axis_bram_67_aresetn),
        .m_axis_bram_67_tlast(m_axis_bram_67_tlast),
        .m_axis_bram_67_tvalid(m_axis_bram_67_tvalid),
        .m_axis_bram_67_tkeep(m_axis_bram_67_tkeep),
        .m_axis_bram_67_tstrb(m_axis_bram_67_tstrb),
        .m_axis_bram_67_tdata(m_axis_bram_67_tdata),
        .m_axis_bram_67_tready(m_axis_bram_67_tready),
        .ap_bram_67_addr0(ap_bram_oarg_67_addr0),
        .ap_bram_67_din0(ap_bram_oarg_67_din0),
        .ap_bram_67_dout0(ap_bram_oarg_67_dout0),
        .ap_bram_67_we0(ap_bram_oarg_67_we0),
        .ap_bram_67_en0(ap_bram_oarg_67_en0),
        .ap_bram_67_addr1(ap_bram_oarg_67_addr1),
        .ap_bram_67_din1(ap_bram_oarg_67_din1),
        .ap_bram_67_dout1(ap_bram_oarg_67_dout1),
        .ap_bram_67_we1(ap_bram_oarg_67_we1),
        .ap_bram_67_en1(ap_bram_oarg_67_en1),
        .m_axis_bram_68_aclk(m_axis_bram_68_aclk),
        .m_axis_bram_68_aresetn(m_axis_bram_68_aresetn),
        .m_axis_bram_68_tlast(m_axis_bram_68_tlast),
        .m_axis_bram_68_tvalid(m_axis_bram_68_tvalid),
        .m_axis_bram_68_tkeep(m_axis_bram_68_tkeep),
        .m_axis_bram_68_tstrb(m_axis_bram_68_tstrb),
        .m_axis_bram_68_tdata(m_axis_bram_68_tdata),
        .m_axis_bram_68_tready(m_axis_bram_68_tready),
        .ap_bram_68_addr0(ap_bram_oarg_68_addr0),
        .ap_bram_68_din0(ap_bram_oarg_68_din0),
        .ap_bram_68_dout0(ap_bram_oarg_68_dout0),
        .ap_bram_68_we0(ap_bram_oarg_68_we0),
        .ap_bram_68_en0(ap_bram_oarg_68_en0),
        .ap_bram_68_addr1(ap_bram_oarg_68_addr1),
        .ap_bram_68_din1(ap_bram_oarg_68_din1),
        .ap_bram_68_dout1(ap_bram_oarg_68_dout1),
        .ap_bram_68_we1(ap_bram_oarg_68_we1),
        .ap_bram_68_en1(ap_bram_oarg_68_en1),
        .m_axis_bram_69_aclk(m_axis_bram_69_aclk),
        .m_axis_bram_69_aresetn(m_axis_bram_69_aresetn),
        .m_axis_bram_69_tlast(m_axis_bram_69_tlast),
        .m_axis_bram_69_tvalid(m_axis_bram_69_tvalid),
        .m_axis_bram_69_tkeep(m_axis_bram_69_tkeep),
        .m_axis_bram_69_tstrb(m_axis_bram_69_tstrb),
        .m_axis_bram_69_tdata(m_axis_bram_69_tdata),
        .m_axis_bram_69_tready(m_axis_bram_69_tready),
        .ap_bram_69_addr0(ap_bram_oarg_69_addr0),
        .ap_bram_69_din0(ap_bram_oarg_69_din0),
        .ap_bram_69_dout0(ap_bram_oarg_69_dout0),
        .ap_bram_69_we0(ap_bram_oarg_69_we0),
        .ap_bram_69_en0(ap_bram_oarg_69_en0),
        .ap_bram_69_addr1(ap_bram_oarg_69_addr1),
        .ap_bram_69_din1(ap_bram_oarg_69_din1),
        .ap_bram_69_dout1(ap_bram_oarg_69_dout1),
        .ap_bram_69_we1(ap_bram_oarg_69_we1),
        .ap_bram_69_en1(ap_bram_oarg_69_en1),
        .m_axis_bram_70_aclk(m_axis_bram_70_aclk),
        .m_axis_bram_70_aresetn(m_axis_bram_70_aresetn),
        .m_axis_bram_70_tlast(m_axis_bram_70_tlast),
        .m_axis_bram_70_tvalid(m_axis_bram_70_tvalid),
        .m_axis_bram_70_tkeep(m_axis_bram_70_tkeep),
        .m_axis_bram_70_tstrb(m_axis_bram_70_tstrb),
        .m_axis_bram_70_tdata(m_axis_bram_70_tdata),
        .m_axis_bram_70_tready(m_axis_bram_70_tready),
        .ap_bram_70_addr0(ap_bram_oarg_70_addr0),
        .ap_bram_70_din0(ap_bram_oarg_70_din0),
        .ap_bram_70_dout0(ap_bram_oarg_70_dout0),
        .ap_bram_70_we0(ap_bram_oarg_70_we0),
        .ap_bram_70_en0(ap_bram_oarg_70_en0),
        .ap_bram_70_addr1(ap_bram_oarg_70_addr1),
        .ap_bram_70_din1(ap_bram_oarg_70_din1),
        .ap_bram_70_dout1(ap_bram_oarg_70_dout1),
        .ap_bram_70_we1(ap_bram_oarg_70_we1),
        .ap_bram_70_en1(ap_bram_oarg_70_en1),
        .m_axis_bram_71_aclk(m_axis_bram_71_aclk),
        .m_axis_bram_71_aresetn(m_axis_bram_71_aresetn),
        .m_axis_bram_71_tlast(m_axis_bram_71_tlast),
        .m_axis_bram_71_tvalid(m_axis_bram_71_tvalid),
        .m_axis_bram_71_tkeep(m_axis_bram_71_tkeep),
        .m_axis_bram_71_tstrb(m_axis_bram_71_tstrb),
        .m_axis_bram_71_tdata(m_axis_bram_71_tdata),
        .m_axis_bram_71_tready(m_axis_bram_71_tready),
        .ap_bram_71_addr0(ap_bram_oarg_71_addr0),
        .ap_bram_71_din0(ap_bram_oarg_71_din0),
        .ap_bram_71_dout0(ap_bram_oarg_71_dout0),
        .ap_bram_71_we0(ap_bram_oarg_71_we0),
        .ap_bram_71_en0(ap_bram_oarg_71_en0),
        .ap_bram_71_addr1(ap_bram_oarg_71_addr1),
        .ap_bram_71_din1(ap_bram_oarg_71_din1),
        .ap_bram_71_dout1(ap_bram_oarg_71_dout1),
        .ap_bram_71_we1(ap_bram_oarg_71_we1),
        .ap_bram_71_en1(ap_bram_oarg_71_en1),
        .m_axis_bram_72_aclk(m_axis_bram_72_aclk),
        .m_axis_bram_72_aresetn(m_axis_bram_72_aresetn),
        .m_axis_bram_72_tlast(m_axis_bram_72_tlast),
        .m_axis_bram_72_tvalid(m_axis_bram_72_tvalid),
        .m_axis_bram_72_tkeep(m_axis_bram_72_tkeep),
        .m_axis_bram_72_tstrb(m_axis_bram_72_tstrb),
        .m_axis_bram_72_tdata(m_axis_bram_72_tdata),
        .m_axis_bram_72_tready(m_axis_bram_72_tready),
        .ap_bram_72_addr0(ap_bram_oarg_72_addr0),
        .ap_bram_72_din0(ap_bram_oarg_72_din0),
        .ap_bram_72_dout0(ap_bram_oarg_72_dout0),
        .ap_bram_72_we0(ap_bram_oarg_72_we0),
        .ap_bram_72_en0(ap_bram_oarg_72_en0),
        .ap_bram_72_addr1(ap_bram_oarg_72_addr1),
        .ap_bram_72_din1(ap_bram_oarg_72_din1),
        .ap_bram_72_dout1(ap_bram_oarg_72_dout1),
        .ap_bram_72_we1(ap_bram_oarg_72_we1),
        .ap_bram_72_en1(ap_bram_oarg_72_en1),
        .m_axis_bram_73_aclk(m_axis_bram_73_aclk),
        .m_axis_bram_73_aresetn(m_axis_bram_73_aresetn),
        .m_axis_bram_73_tlast(m_axis_bram_73_tlast),
        .m_axis_bram_73_tvalid(m_axis_bram_73_tvalid),
        .m_axis_bram_73_tkeep(m_axis_bram_73_tkeep),
        .m_axis_bram_73_tstrb(m_axis_bram_73_tstrb),
        .m_axis_bram_73_tdata(m_axis_bram_73_tdata),
        .m_axis_bram_73_tready(m_axis_bram_73_tready),
        .ap_bram_73_addr0(ap_bram_oarg_73_addr0),
        .ap_bram_73_din0(ap_bram_oarg_73_din0),
        .ap_bram_73_dout0(ap_bram_oarg_73_dout0),
        .ap_bram_73_we0(ap_bram_oarg_73_we0),
        .ap_bram_73_en0(ap_bram_oarg_73_en0),
        .ap_bram_73_addr1(ap_bram_oarg_73_addr1),
        .ap_bram_73_din1(ap_bram_oarg_73_din1),
        .ap_bram_73_dout1(ap_bram_oarg_73_dout1),
        .ap_bram_73_we1(ap_bram_oarg_73_we1),
        .ap_bram_73_en1(ap_bram_oarg_73_en1),
        .m_axis_bram_74_aclk(m_axis_bram_74_aclk),
        .m_axis_bram_74_aresetn(m_axis_bram_74_aresetn),
        .m_axis_bram_74_tlast(m_axis_bram_74_tlast),
        .m_axis_bram_74_tvalid(m_axis_bram_74_tvalid),
        .m_axis_bram_74_tkeep(m_axis_bram_74_tkeep),
        .m_axis_bram_74_tstrb(m_axis_bram_74_tstrb),
        .m_axis_bram_74_tdata(m_axis_bram_74_tdata),
        .m_axis_bram_74_tready(m_axis_bram_74_tready),
        .ap_bram_74_addr0(ap_bram_oarg_74_addr0),
        .ap_bram_74_din0(ap_bram_oarg_74_din0),
        .ap_bram_74_dout0(ap_bram_oarg_74_dout0),
        .ap_bram_74_we0(ap_bram_oarg_74_we0),
        .ap_bram_74_en0(ap_bram_oarg_74_en0),
        .ap_bram_74_addr1(ap_bram_oarg_74_addr1),
        .ap_bram_74_din1(ap_bram_oarg_74_din1),
        .ap_bram_74_dout1(ap_bram_oarg_74_dout1),
        .ap_bram_74_we1(ap_bram_oarg_74_we1),
        .ap_bram_74_en1(ap_bram_oarg_74_en1),
        .m_axis_bram_75_aclk(m_axis_bram_75_aclk),
        .m_axis_bram_75_aresetn(m_axis_bram_75_aresetn),
        .m_axis_bram_75_tlast(m_axis_bram_75_tlast),
        .m_axis_bram_75_tvalid(m_axis_bram_75_tvalid),
        .m_axis_bram_75_tkeep(m_axis_bram_75_tkeep),
        .m_axis_bram_75_tstrb(m_axis_bram_75_tstrb),
        .m_axis_bram_75_tdata(m_axis_bram_75_tdata),
        .m_axis_bram_75_tready(m_axis_bram_75_tready),
        .ap_bram_75_addr0(ap_bram_oarg_75_addr0),
        .ap_bram_75_din0(ap_bram_oarg_75_din0),
        .ap_bram_75_dout0(ap_bram_oarg_75_dout0),
        .ap_bram_75_we0(ap_bram_oarg_75_we0),
        .ap_bram_75_en0(ap_bram_oarg_75_en0),
        .ap_bram_75_addr1(ap_bram_oarg_75_addr1),
        .ap_bram_75_din1(ap_bram_oarg_75_din1),
        .ap_bram_75_dout1(ap_bram_oarg_75_dout1),
        .ap_bram_75_we1(ap_bram_oarg_75_we1),
        .ap_bram_75_en1(ap_bram_oarg_75_en1),
        .m_axis_bram_76_aclk(m_axis_bram_76_aclk),
        .m_axis_bram_76_aresetn(m_axis_bram_76_aresetn),
        .m_axis_bram_76_tlast(m_axis_bram_76_tlast),
        .m_axis_bram_76_tvalid(m_axis_bram_76_tvalid),
        .m_axis_bram_76_tkeep(m_axis_bram_76_tkeep),
        .m_axis_bram_76_tstrb(m_axis_bram_76_tstrb),
        .m_axis_bram_76_tdata(m_axis_bram_76_tdata),
        .m_axis_bram_76_tready(m_axis_bram_76_tready),
        .ap_bram_76_addr0(ap_bram_oarg_76_addr0),
        .ap_bram_76_din0(ap_bram_oarg_76_din0),
        .ap_bram_76_dout0(ap_bram_oarg_76_dout0),
        .ap_bram_76_we0(ap_bram_oarg_76_we0),
        .ap_bram_76_en0(ap_bram_oarg_76_en0),
        .ap_bram_76_addr1(ap_bram_oarg_76_addr1),
        .ap_bram_76_din1(ap_bram_oarg_76_din1),
        .ap_bram_76_dout1(ap_bram_oarg_76_dout1),
        .ap_bram_76_we1(ap_bram_oarg_76_we1),
        .ap_bram_76_en1(ap_bram_oarg_76_en1),
        .m_axis_bram_77_aclk(m_axis_bram_77_aclk),
        .m_axis_bram_77_aresetn(m_axis_bram_77_aresetn),
        .m_axis_bram_77_tlast(m_axis_bram_77_tlast),
        .m_axis_bram_77_tvalid(m_axis_bram_77_tvalid),
        .m_axis_bram_77_tkeep(m_axis_bram_77_tkeep),
        .m_axis_bram_77_tstrb(m_axis_bram_77_tstrb),
        .m_axis_bram_77_tdata(m_axis_bram_77_tdata),
        .m_axis_bram_77_tready(m_axis_bram_77_tready),
        .ap_bram_77_addr0(ap_bram_oarg_77_addr0),
        .ap_bram_77_din0(ap_bram_oarg_77_din0),
        .ap_bram_77_dout0(ap_bram_oarg_77_dout0),
        .ap_bram_77_we0(ap_bram_oarg_77_we0),
        .ap_bram_77_en0(ap_bram_oarg_77_en0),
        .ap_bram_77_addr1(ap_bram_oarg_77_addr1),
        .ap_bram_77_din1(ap_bram_oarg_77_din1),
        .ap_bram_77_dout1(ap_bram_oarg_77_dout1),
        .ap_bram_77_we1(ap_bram_oarg_77_we1),
        .ap_bram_77_en1(ap_bram_oarg_77_en1),
        .m_axis_bram_78_aclk(m_axis_bram_78_aclk),
        .m_axis_bram_78_aresetn(m_axis_bram_78_aresetn),
        .m_axis_bram_78_tlast(m_axis_bram_78_tlast),
        .m_axis_bram_78_tvalid(m_axis_bram_78_tvalid),
        .m_axis_bram_78_tkeep(m_axis_bram_78_tkeep),
        .m_axis_bram_78_tstrb(m_axis_bram_78_tstrb),
        .m_axis_bram_78_tdata(m_axis_bram_78_tdata),
        .m_axis_bram_78_tready(m_axis_bram_78_tready),
        .ap_bram_78_addr0(ap_bram_oarg_78_addr0),
        .ap_bram_78_din0(ap_bram_oarg_78_din0),
        .ap_bram_78_dout0(ap_bram_oarg_78_dout0),
        .ap_bram_78_we0(ap_bram_oarg_78_we0),
        .ap_bram_78_en0(ap_bram_oarg_78_en0),
        .ap_bram_78_addr1(ap_bram_oarg_78_addr1),
        .ap_bram_78_din1(ap_bram_oarg_78_din1),
        .ap_bram_78_dout1(ap_bram_oarg_78_dout1),
        .ap_bram_78_we1(ap_bram_oarg_78_we1),
        .ap_bram_78_en1(ap_bram_oarg_78_en1),
        .m_axis_bram_79_aclk(m_axis_bram_79_aclk),
        .m_axis_bram_79_aresetn(m_axis_bram_79_aresetn),
        .m_axis_bram_79_tlast(m_axis_bram_79_tlast),
        .m_axis_bram_79_tvalid(m_axis_bram_79_tvalid),
        .m_axis_bram_79_tkeep(m_axis_bram_79_tkeep),
        .m_axis_bram_79_tstrb(m_axis_bram_79_tstrb),
        .m_axis_bram_79_tdata(m_axis_bram_79_tdata),
        .m_axis_bram_79_tready(m_axis_bram_79_tready),
        .ap_bram_79_addr0(ap_bram_oarg_79_addr0),
        .ap_bram_79_din0(ap_bram_oarg_79_din0),
        .ap_bram_79_dout0(ap_bram_oarg_79_dout0),
        .ap_bram_79_we0(ap_bram_oarg_79_we0),
        .ap_bram_79_en0(ap_bram_oarg_79_en0),
        .ap_bram_79_addr1(ap_bram_oarg_79_addr1),
        .ap_bram_79_din1(ap_bram_oarg_79_din1),
        .ap_bram_79_dout1(ap_bram_oarg_79_dout1),
        .ap_bram_79_we1(ap_bram_oarg_79_we1),
        .ap_bram_79_en1(ap_bram_oarg_79_en1),
        .m_axis_bram_80_aclk(m_axis_bram_80_aclk),
        .m_axis_bram_80_aresetn(m_axis_bram_80_aresetn),
        .m_axis_bram_80_tlast(m_axis_bram_80_tlast),
        .m_axis_bram_80_tvalid(m_axis_bram_80_tvalid),
        .m_axis_bram_80_tkeep(m_axis_bram_80_tkeep),
        .m_axis_bram_80_tstrb(m_axis_bram_80_tstrb),
        .m_axis_bram_80_tdata(m_axis_bram_80_tdata),
        .m_axis_bram_80_tready(m_axis_bram_80_tready),
        .ap_bram_80_addr0(ap_bram_oarg_80_addr0),
        .ap_bram_80_din0(ap_bram_oarg_80_din0),
        .ap_bram_80_dout0(ap_bram_oarg_80_dout0),
        .ap_bram_80_we0(ap_bram_oarg_80_we0),
        .ap_bram_80_en0(ap_bram_oarg_80_en0),
        .ap_bram_80_addr1(ap_bram_oarg_80_addr1),
        .ap_bram_80_din1(ap_bram_oarg_80_din1),
        .ap_bram_80_dout1(ap_bram_oarg_80_dout1),
        .ap_bram_80_we1(ap_bram_oarg_80_we1),
        .ap_bram_80_en1(ap_bram_oarg_80_en1),
        .m_axis_bram_81_aclk(m_axis_bram_81_aclk),
        .m_axis_bram_81_aresetn(m_axis_bram_81_aresetn),
        .m_axis_bram_81_tlast(m_axis_bram_81_tlast),
        .m_axis_bram_81_tvalid(m_axis_bram_81_tvalid),
        .m_axis_bram_81_tkeep(m_axis_bram_81_tkeep),
        .m_axis_bram_81_tstrb(m_axis_bram_81_tstrb),
        .m_axis_bram_81_tdata(m_axis_bram_81_tdata),
        .m_axis_bram_81_tready(m_axis_bram_81_tready),
        .ap_bram_81_addr0(ap_bram_oarg_81_addr0),
        .ap_bram_81_din0(ap_bram_oarg_81_din0),
        .ap_bram_81_dout0(ap_bram_oarg_81_dout0),
        .ap_bram_81_we0(ap_bram_oarg_81_we0),
        .ap_bram_81_en0(ap_bram_oarg_81_en0),
        .ap_bram_81_addr1(ap_bram_oarg_81_addr1),
        .ap_bram_81_din1(ap_bram_oarg_81_din1),
        .ap_bram_81_dout1(ap_bram_oarg_81_dout1),
        .ap_bram_81_we1(ap_bram_oarg_81_we1),
        .ap_bram_81_en1(ap_bram_oarg_81_en1),
        .m_axis_bram_82_aclk(m_axis_bram_82_aclk),
        .m_axis_bram_82_aresetn(m_axis_bram_82_aresetn),
        .m_axis_bram_82_tlast(m_axis_bram_82_tlast),
        .m_axis_bram_82_tvalid(m_axis_bram_82_tvalid),
        .m_axis_bram_82_tkeep(m_axis_bram_82_tkeep),
        .m_axis_bram_82_tstrb(m_axis_bram_82_tstrb),
        .m_axis_bram_82_tdata(m_axis_bram_82_tdata),
        .m_axis_bram_82_tready(m_axis_bram_82_tready),
        .ap_bram_82_addr0(ap_bram_oarg_82_addr0),
        .ap_bram_82_din0(ap_bram_oarg_82_din0),
        .ap_bram_82_dout0(ap_bram_oarg_82_dout0),
        .ap_bram_82_we0(ap_bram_oarg_82_we0),
        .ap_bram_82_en0(ap_bram_oarg_82_en0),
        .ap_bram_82_addr1(ap_bram_oarg_82_addr1),
        .ap_bram_82_din1(ap_bram_oarg_82_din1),
        .ap_bram_82_dout1(ap_bram_oarg_82_dout1),
        .ap_bram_82_we1(ap_bram_oarg_82_we1),
        .ap_bram_82_en1(ap_bram_oarg_82_en1),
        .m_axis_bram_83_aclk(m_axis_bram_83_aclk),
        .m_axis_bram_83_aresetn(m_axis_bram_83_aresetn),
        .m_axis_bram_83_tlast(m_axis_bram_83_tlast),
        .m_axis_bram_83_tvalid(m_axis_bram_83_tvalid),
        .m_axis_bram_83_tkeep(m_axis_bram_83_tkeep),
        .m_axis_bram_83_tstrb(m_axis_bram_83_tstrb),
        .m_axis_bram_83_tdata(m_axis_bram_83_tdata),
        .m_axis_bram_83_tready(m_axis_bram_83_tready),
        .ap_bram_83_addr0(ap_bram_oarg_83_addr0),
        .ap_bram_83_din0(ap_bram_oarg_83_din0),
        .ap_bram_83_dout0(ap_bram_oarg_83_dout0),
        .ap_bram_83_we0(ap_bram_oarg_83_we0),
        .ap_bram_83_en0(ap_bram_oarg_83_en0),
        .ap_bram_83_addr1(ap_bram_oarg_83_addr1),
        .ap_bram_83_din1(ap_bram_oarg_83_din1),
        .ap_bram_83_dout1(ap_bram_oarg_83_dout1),
        .ap_bram_83_we1(ap_bram_oarg_83_we1),
        .ap_bram_83_en1(ap_bram_oarg_83_en1),
        .m_axis_bram_84_aclk(m_axis_bram_84_aclk),
        .m_axis_bram_84_aresetn(m_axis_bram_84_aresetn),
        .m_axis_bram_84_tlast(m_axis_bram_84_tlast),
        .m_axis_bram_84_tvalid(m_axis_bram_84_tvalid),
        .m_axis_bram_84_tkeep(m_axis_bram_84_tkeep),
        .m_axis_bram_84_tstrb(m_axis_bram_84_tstrb),
        .m_axis_bram_84_tdata(m_axis_bram_84_tdata),
        .m_axis_bram_84_tready(m_axis_bram_84_tready),
        .ap_bram_84_addr0(ap_bram_oarg_84_addr0),
        .ap_bram_84_din0(ap_bram_oarg_84_din0),
        .ap_bram_84_dout0(ap_bram_oarg_84_dout0),
        .ap_bram_84_we0(ap_bram_oarg_84_we0),
        .ap_bram_84_en0(ap_bram_oarg_84_en0),
        .ap_bram_84_addr1(ap_bram_oarg_84_addr1),
        .ap_bram_84_din1(ap_bram_oarg_84_din1),
        .ap_bram_84_dout1(ap_bram_oarg_84_dout1),
        .ap_bram_84_we1(ap_bram_oarg_84_we1),
        .ap_bram_84_en1(ap_bram_oarg_84_en1),
        .m_axis_bram_85_aclk(m_axis_bram_85_aclk),
        .m_axis_bram_85_aresetn(m_axis_bram_85_aresetn),
        .m_axis_bram_85_tlast(m_axis_bram_85_tlast),
        .m_axis_bram_85_tvalid(m_axis_bram_85_tvalid),
        .m_axis_bram_85_tkeep(m_axis_bram_85_tkeep),
        .m_axis_bram_85_tstrb(m_axis_bram_85_tstrb),
        .m_axis_bram_85_tdata(m_axis_bram_85_tdata),
        .m_axis_bram_85_tready(m_axis_bram_85_tready),
        .ap_bram_85_addr0(ap_bram_oarg_85_addr0),
        .ap_bram_85_din0(ap_bram_oarg_85_din0),
        .ap_bram_85_dout0(ap_bram_oarg_85_dout0),
        .ap_bram_85_we0(ap_bram_oarg_85_we0),
        .ap_bram_85_en0(ap_bram_oarg_85_en0),
        .ap_bram_85_addr1(ap_bram_oarg_85_addr1),
        .ap_bram_85_din1(ap_bram_oarg_85_din1),
        .ap_bram_85_dout1(ap_bram_oarg_85_dout1),
        .ap_bram_85_we1(ap_bram_oarg_85_we1),
        .ap_bram_85_en1(ap_bram_oarg_85_en1),
        .m_axis_bram_86_aclk(m_axis_bram_86_aclk),
        .m_axis_bram_86_aresetn(m_axis_bram_86_aresetn),
        .m_axis_bram_86_tlast(m_axis_bram_86_tlast),
        .m_axis_bram_86_tvalid(m_axis_bram_86_tvalid),
        .m_axis_bram_86_tkeep(m_axis_bram_86_tkeep),
        .m_axis_bram_86_tstrb(m_axis_bram_86_tstrb),
        .m_axis_bram_86_tdata(m_axis_bram_86_tdata),
        .m_axis_bram_86_tready(m_axis_bram_86_tready),
        .ap_bram_86_addr0(ap_bram_oarg_86_addr0),
        .ap_bram_86_din0(ap_bram_oarg_86_din0),
        .ap_bram_86_dout0(ap_bram_oarg_86_dout0),
        .ap_bram_86_we0(ap_bram_oarg_86_we0),
        .ap_bram_86_en0(ap_bram_oarg_86_en0),
        .ap_bram_86_addr1(ap_bram_oarg_86_addr1),
        .ap_bram_86_din1(ap_bram_oarg_86_din1),
        .ap_bram_86_dout1(ap_bram_oarg_86_dout1),
        .ap_bram_86_we1(ap_bram_oarg_86_we1),
        .ap_bram_86_en1(ap_bram_oarg_86_en1),
        .m_axis_bram_87_aclk(m_axis_bram_87_aclk),
        .m_axis_bram_87_aresetn(m_axis_bram_87_aresetn),
        .m_axis_bram_87_tlast(m_axis_bram_87_tlast),
        .m_axis_bram_87_tvalid(m_axis_bram_87_tvalid),
        .m_axis_bram_87_tkeep(m_axis_bram_87_tkeep),
        .m_axis_bram_87_tstrb(m_axis_bram_87_tstrb),
        .m_axis_bram_87_tdata(m_axis_bram_87_tdata),
        .m_axis_bram_87_tready(m_axis_bram_87_tready),
        .ap_bram_87_addr0(ap_bram_oarg_87_addr0),
        .ap_bram_87_din0(ap_bram_oarg_87_din0),
        .ap_bram_87_dout0(ap_bram_oarg_87_dout0),
        .ap_bram_87_we0(ap_bram_oarg_87_we0),
        .ap_bram_87_en0(ap_bram_oarg_87_en0),
        .ap_bram_87_addr1(ap_bram_oarg_87_addr1),
        .ap_bram_87_din1(ap_bram_oarg_87_din1),
        .ap_bram_87_dout1(ap_bram_oarg_87_dout1),
        .ap_bram_87_we1(ap_bram_oarg_87_we1),
        .ap_bram_87_en1(ap_bram_oarg_87_en1),
        .m_axis_bram_88_aclk(m_axis_bram_88_aclk),
        .m_axis_bram_88_aresetn(m_axis_bram_88_aresetn),
        .m_axis_bram_88_tlast(m_axis_bram_88_tlast),
        .m_axis_bram_88_tvalid(m_axis_bram_88_tvalid),
        .m_axis_bram_88_tkeep(m_axis_bram_88_tkeep),
        .m_axis_bram_88_tstrb(m_axis_bram_88_tstrb),
        .m_axis_bram_88_tdata(m_axis_bram_88_tdata),
        .m_axis_bram_88_tready(m_axis_bram_88_tready),
        .ap_bram_88_addr0(ap_bram_oarg_88_addr0),
        .ap_bram_88_din0(ap_bram_oarg_88_din0),
        .ap_bram_88_dout0(ap_bram_oarg_88_dout0),
        .ap_bram_88_we0(ap_bram_oarg_88_we0),
        .ap_bram_88_en0(ap_bram_oarg_88_en0),
        .ap_bram_88_addr1(ap_bram_oarg_88_addr1),
        .ap_bram_88_din1(ap_bram_oarg_88_din1),
        .ap_bram_88_dout1(ap_bram_oarg_88_dout1),
        .ap_bram_88_we1(ap_bram_oarg_88_we1),
        .ap_bram_88_en1(ap_bram_oarg_88_en1),
        .m_axis_bram_89_aclk(m_axis_bram_89_aclk),
        .m_axis_bram_89_aresetn(m_axis_bram_89_aresetn),
        .m_axis_bram_89_tlast(m_axis_bram_89_tlast),
        .m_axis_bram_89_tvalid(m_axis_bram_89_tvalid),
        .m_axis_bram_89_tkeep(m_axis_bram_89_tkeep),
        .m_axis_bram_89_tstrb(m_axis_bram_89_tstrb),
        .m_axis_bram_89_tdata(m_axis_bram_89_tdata),
        .m_axis_bram_89_tready(m_axis_bram_89_tready),
        .ap_bram_89_addr0(ap_bram_oarg_89_addr0),
        .ap_bram_89_din0(ap_bram_oarg_89_din0),
        .ap_bram_89_dout0(ap_bram_oarg_89_dout0),
        .ap_bram_89_we0(ap_bram_oarg_89_we0),
        .ap_bram_89_en0(ap_bram_oarg_89_en0),
        .ap_bram_89_addr1(ap_bram_oarg_89_addr1),
        .ap_bram_89_din1(ap_bram_oarg_89_din1),
        .ap_bram_89_dout1(ap_bram_oarg_89_dout1),
        .ap_bram_89_we1(ap_bram_oarg_89_we1),
        .ap_bram_89_en1(ap_bram_oarg_89_en1),
        .m_axis_bram_90_aclk(m_axis_bram_90_aclk),
        .m_axis_bram_90_aresetn(m_axis_bram_90_aresetn),
        .m_axis_bram_90_tlast(m_axis_bram_90_tlast),
        .m_axis_bram_90_tvalid(m_axis_bram_90_tvalid),
        .m_axis_bram_90_tkeep(m_axis_bram_90_tkeep),
        .m_axis_bram_90_tstrb(m_axis_bram_90_tstrb),
        .m_axis_bram_90_tdata(m_axis_bram_90_tdata),
        .m_axis_bram_90_tready(m_axis_bram_90_tready),
        .ap_bram_90_addr0(ap_bram_oarg_90_addr0),
        .ap_bram_90_din0(ap_bram_oarg_90_din0),
        .ap_bram_90_dout0(ap_bram_oarg_90_dout0),
        .ap_bram_90_we0(ap_bram_oarg_90_we0),
        .ap_bram_90_en0(ap_bram_oarg_90_en0),
        .ap_bram_90_addr1(ap_bram_oarg_90_addr1),
        .ap_bram_90_din1(ap_bram_oarg_90_din1),
        .ap_bram_90_dout1(ap_bram_oarg_90_dout1),
        .ap_bram_90_we1(ap_bram_oarg_90_we1),
        .ap_bram_90_en1(ap_bram_oarg_90_en1),
        .m_axis_bram_91_aclk(m_axis_bram_91_aclk),
        .m_axis_bram_91_aresetn(m_axis_bram_91_aresetn),
        .m_axis_bram_91_tlast(m_axis_bram_91_tlast),
        .m_axis_bram_91_tvalid(m_axis_bram_91_tvalid),
        .m_axis_bram_91_tkeep(m_axis_bram_91_tkeep),
        .m_axis_bram_91_tstrb(m_axis_bram_91_tstrb),
        .m_axis_bram_91_tdata(m_axis_bram_91_tdata),
        .m_axis_bram_91_tready(m_axis_bram_91_tready),
        .ap_bram_91_addr0(ap_bram_oarg_91_addr0),
        .ap_bram_91_din0(ap_bram_oarg_91_din0),
        .ap_bram_91_dout0(ap_bram_oarg_91_dout0),
        .ap_bram_91_we0(ap_bram_oarg_91_we0),
        .ap_bram_91_en0(ap_bram_oarg_91_en0),
        .ap_bram_91_addr1(ap_bram_oarg_91_addr1),
        .ap_bram_91_din1(ap_bram_oarg_91_din1),
        .ap_bram_91_dout1(ap_bram_oarg_91_dout1),
        .ap_bram_91_we1(ap_bram_oarg_91_we1),
        .ap_bram_91_en1(ap_bram_oarg_91_en1),
        .m_axis_bram_92_aclk(m_axis_bram_92_aclk),
        .m_axis_bram_92_aresetn(m_axis_bram_92_aresetn),
        .m_axis_bram_92_tlast(m_axis_bram_92_tlast),
        .m_axis_bram_92_tvalid(m_axis_bram_92_tvalid),
        .m_axis_bram_92_tkeep(m_axis_bram_92_tkeep),
        .m_axis_bram_92_tstrb(m_axis_bram_92_tstrb),
        .m_axis_bram_92_tdata(m_axis_bram_92_tdata),
        .m_axis_bram_92_tready(m_axis_bram_92_tready),
        .ap_bram_92_addr0(ap_bram_oarg_92_addr0),
        .ap_bram_92_din0(ap_bram_oarg_92_din0),
        .ap_bram_92_dout0(ap_bram_oarg_92_dout0),
        .ap_bram_92_we0(ap_bram_oarg_92_we0),
        .ap_bram_92_en0(ap_bram_oarg_92_en0),
        .ap_bram_92_addr1(ap_bram_oarg_92_addr1),
        .ap_bram_92_din1(ap_bram_oarg_92_din1),
        .ap_bram_92_dout1(ap_bram_oarg_92_dout1),
        .ap_bram_92_we1(ap_bram_oarg_92_we1),
        .ap_bram_92_en1(ap_bram_oarg_92_en1),
        .m_axis_bram_93_aclk(m_axis_bram_93_aclk),
        .m_axis_bram_93_aresetn(m_axis_bram_93_aresetn),
        .m_axis_bram_93_tlast(m_axis_bram_93_tlast),
        .m_axis_bram_93_tvalid(m_axis_bram_93_tvalid),
        .m_axis_bram_93_tkeep(m_axis_bram_93_tkeep),
        .m_axis_bram_93_tstrb(m_axis_bram_93_tstrb),
        .m_axis_bram_93_tdata(m_axis_bram_93_tdata),
        .m_axis_bram_93_tready(m_axis_bram_93_tready),
        .ap_bram_93_addr0(ap_bram_oarg_93_addr0),
        .ap_bram_93_din0(ap_bram_oarg_93_din0),
        .ap_bram_93_dout0(ap_bram_oarg_93_dout0),
        .ap_bram_93_we0(ap_bram_oarg_93_we0),
        .ap_bram_93_en0(ap_bram_oarg_93_en0),
        .ap_bram_93_addr1(ap_bram_oarg_93_addr1),
        .ap_bram_93_din1(ap_bram_oarg_93_din1),
        .ap_bram_93_dout1(ap_bram_oarg_93_dout1),
        .ap_bram_93_we1(ap_bram_oarg_93_we1),
        .ap_bram_93_en1(ap_bram_oarg_93_en1),
        .m_axis_bram_94_aclk(m_axis_bram_94_aclk),
        .m_axis_bram_94_aresetn(m_axis_bram_94_aresetn),
        .m_axis_bram_94_tlast(m_axis_bram_94_tlast),
        .m_axis_bram_94_tvalid(m_axis_bram_94_tvalid),
        .m_axis_bram_94_tkeep(m_axis_bram_94_tkeep),
        .m_axis_bram_94_tstrb(m_axis_bram_94_tstrb),
        .m_axis_bram_94_tdata(m_axis_bram_94_tdata),
        .m_axis_bram_94_tready(m_axis_bram_94_tready),
        .ap_bram_94_addr0(ap_bram_oarg_94_addr0),
        .ap_bram_94_din0(ap_bram_oarg_94_din0),
        .ap_bram_94_dout0(ap_bram_oarg_94_dout0),
        .ap_bram_94_we0(ap_bram_oarg_94_we0),
        .ap_bram_94_en0(ap_bram_oarg_94_en0),
        .ap_bram_94_addr1(ap_bram_oarg_94_addr1),
        .ap_bram_94_din1(ap_bram_oarg_94_din1),
        .ap_bram_94_dout1(ap_bram_oarg_94_dout1),
        .ap_bram_94_we1(ap_bram_oarg_94_we1),
        .ap_bram_94_en1(ap_bram_oarg_94_en1),
        .m_axis_bram_95_aclk(m_axis_bram_95_aclk),
        .m_axis_bram_95_aresetn(m_axis_bram_95_aresetn),
        .m_axis_bram_95_tlast(m_axis_bram_95_tlast),
        .m_axis_bram_95_tvalid(m_axis_bram_95_tvalid),
        .m_axis_bram_95_tkeep(m_axis_bram_95_tkeep),
        .m_axis_bram_95_tstrb(m_axis_bram_95_tstrb),
        .m_axis_bram_95_tdata(m_axis_bram_95_tdata),
        .m_axis_bram_95_tready(m_axis_bram_95_tready),
        .ap_bram_95_addr0(ap_bram_oarg_95_addr0),
        .ap_bram_95_din0(ap_bram_oarg_95_din0),
        .ap_bram_95_dout0(ap_bram_oarg_95_dout0),
        .ap_bram_95_we0(ap_bram_oarg_95_we0),
        .ap_bram_95_en0(ap_bram_oarg_95_en0),
        .ap_bram_95_addr1(ap_bram_oarg_95_addr1),
        .ap_bram_95_din1(ap_bram_oarg_95_din1),
        .ap_bram_95_dout1(ap_bram_oarg_95_dout1),
        .ap_bram_95_we1(ap_bram_oarg_95_we1),
        .ap_bram_95_en1(ap_bram_oarg_95_en1),
        .m_axis_bram_96_aclk(m_axis_bram_96_aclk),
        .m_axis_bram_96_aresetn(m_axis_bram_96_aresetn),
        .m_axis_bram_96_tlast(m_axis_bram_96_tlast),
        .m_axis_bram_96_tvalid(m_axis_bram_96_tvalid),
        .m_axis_bram_96_tkeep(m_axis_bram_96_tkeep),
        .m_axis_bram_96_tstrb(m_axis_bram_96_tstrb),
        .m_axis_bram_96_tdata(m_axis_bram_96_tdata),
        .m_axis_bram_96_tready(m_axis_bram_96_tready),
        .ap_bram_96_addr0(ap_bram_oarg_96_addr0),
        .ap_bram_96_din0(ap_bram_oarg_96_din0),
        .ap_bram_96_dout0(ap_bram_oarg_96_dout0),
        .ap_bram_96_we0(ap_bram_oarg_96_we0),
        .ap_bram_96_en0(ap_bram_oarg_96_en0),
        .ap_bram_96_addr1(ap_bram_oarg_96_addr1),
        .ap_bram_96_din1(ap_bram_oarg_96_din1),
        .ap_bram_96_dout1(ap_bram_oarg_96_dout1),
        .ap_bram_96_we1(ap_bram_oarg_96_we1),
        .ap_bram_96_en1(ap_bram_oarg_96_en1),
        .m_axis_bram_97_aclk(m_axis_bram_97_aclk),
        .m_axis_bram_97_aresetn(m_axis_bram_97_aresetn),
        .m_axis_bram_97_tlast(m_axis_bram_97_tlast),
        .m_axis_bram_97_tvalid(m_axis_bram_97_tvalid),
        .m_axis_bram_97_tkeep(m_axis_bram_97_tkeep),
        .m_axis_bram_97_tstrb(m_axis_bram_97_tstrb),
        .m_axis_bram_97_tdata(m_axis_bram_97_tdata),
        .m_axis_bram_97_tready(m_axis_bram_97_tready),
        .ap_bram_97_addr0(ap_bram_oarg_97_addr0),
        .ap_bram_97_din0(ap_bram_oarg_97_din0),
        .ap_bram_97_dout0(ap_bram_oarg_97_dout0),
        .ap_bram_97_we0(ap_bram_oarg_97_we0),
        .ap_bram_97_en0(ap_bram_oarg_97_en0),
        .ap_bram_97_addr1(ap_bram_oarg_97_addr1),
        .ap_bram_97_din1(ap_bram_oarg_97_din1),
        .ap_bram_97_dout1(ap_bram_oarg_97_dout1),
        .ap_bram_97_we1(ap_bram_oarg_97_we1),
        .ap_bram_97_en1(ap_bram_oarg_97_en1),
        .m_axis_bram_98_aclk(m_axis_bram_98_aclk),
        .m_axis_bram_98_aresetn(m_axis_bram_98_aresetn),
        .m_axis_bram_98_tlast(m_axis_bram_98_tlast),
        .m_axis_bram_98_tvalid(m_axis_bram_98_tvalid),
        .m_axis_bram_98_tkeep(m_axis_bram_98_tkeep),
        .m_axis_bram_98_tstrb(m_axis_bram_98_tstrb),
        .m_axis_bram_98_tdata(m_axis_bram_98_tdata),
        .m_axis_bram_98_tready(m_axis_bram_98_tready),
        .ap_bram_98_addr0(ap_bram_oarg_98_addr0),
        .ap_bram_98_din0(ap_bram_oarg_98_din0),
        .ap_bram_98_dout0(ap_bram_oarg_98_dout0),
        .ap_bram_98_we0(ap_bram_oarg_98_we0),
        .ap_bram_98_en0(ap_bram_oarg_98_en0),
        .ap_bram_98_addr1(ap_bram_oarg_98_addr1),
        .ap_bram_98_din1(ap_bram_oarg_98_din1),
        .ap_bram_98_dout1(ap_bram_oarg_98_dout1),
        .ap_bram_98_we1(ap_bram_oarg_98_we1),
        .ap_bram_98_en1(ap_bram_oarg_98_en1),
        .m_axis_bram_99_aclk(m_axis_bram_99_aclk),
        .m_axis_bram_99_aresetn(m_axis_bram_99_aresetn),
        .m_axis_bram_99_tlast(m_axis_bram_99_tlast),
        .m_axis_bram_99_tvalid(m_axis_bram_99_tvalid),
        .m_axis_bram_99_tkeep(m_axis_bram_99_tkeep),
        .m_axis_bram_99_tstrb(m_axis_bram_99_tstrb),
        .m_axis_bram_99_tdata(m_axis_bram_99_tdata),
        .m_axis_bram_99_tready(m_axis_bram_99_tready),
        .ap_bram_99_addr0(ap_bram_oarg_99_addr0),
        .ap_bram_99_din0(ap_bram_oarg_99_din0),
        .ap_bram_99_dout0(ap_bram_oarg_99_dout0),
        .ap_bram_99_we0(ap_bram_oarg_99_we0),
        .ap_bram_99_en0(ap_bram_oarg_99_en0),
        .ap_bram_99_addr1(ap_bram_oarg_99_addr1),
        .ap_bram_99_din1(ap_bram_oarg_99_din1),
        .ap_bram_99_dout1(ap_bram_oarg_99_dout1),
        .ap_bram_99_we1(ap_bram_oarg_99_we1),
        .ap_bram_99_en1(ap_bram_oarg_99_en1),
        .m_axis_bram_100_aclk(m_axis_bram_100_aclk),
        .m_axis_bram_100_aresetn(m_axis_bram_100_aresetn),
        .m_axis_bram_100_tlast(m_axis_bram_100_tlast),
        .m_axis_bram_100_tvalid(m_axis_bram_100_tvalid),
        .m_axis_bram_100_tkeep(m_axis_bram_100_tkeep),
        .m_axis_bram_100_tstrb(m_axis_bram_100_tstrb),
        .m_axis_bram_100_tdata(m_axis_bram_100_tdata),
        .m_axis_bram_100_tready(m_axis_bram_100_tready),
        .ap_bram_100_addr0(ap_bram_oarg_100_addr0),
        .ap_bram_100_din0(ap_bram_oarg_100_din0),
        .ap_bram_100_dout0(ap_bram_oarg_100_dout0),
        .ap_bram_100_we0(ap_bram_oarg_100_we0),
        .ap_bram_100_en0(ap_bram_oarg_100_en0),
        .ap_bram_100_addr1(ap_bram_oarg_100_addr1),
        .ap_bram_100_din1(ap_bram_oarg_100_din1),
        .ap_bram_100_dout1(ap_bram_oarg_100_dout1),
        .ap_bram_100_we1(ap_bram_oarg_100_we1),
        .ap_bram_100_en1(ap_bram_oarg_100_en1),
        .m_axis_bram_101_aclk(m_axis_bram_101_aclk),
        .m_axis_bram_101_aresetn(m_axis_bram_101_aresetn),
        .m_axis_bram_101_tlast(m_axis_bram_101_tlast),
        .m_axis_bram_101_tvalid(m_axis_bram_101_tvalid),
        .m_axis_bram_101_tkeep(m_axis_bram_101_tkeep),
        .m_axis_bram_101_tstrb(m_axis_bram_101_tstrb),
        .m_axis_bram_101_tdata(m_axis_bram_101_tdata),
        .m_axis_bram_101_tready(m_axis_bram_101_tready),
        .ap_bram_101_addr0(ap_bram_oarg_101_addr0),
        .ap_bram_101_din0(ap_bram_oarg_101_din0),
        .ap_bram_101_dout0(ap_bram_oarg_101_dout0),
        .ap_bram_101_we0(ap_bram_oarg_101_we0),
        .ap_bram_101_en0(ap_bram_oarg_101_en0),
        .ap_bram_101_addr1(ap_bram_oarg_101_addr1),
        .ap_bram_101_din1(ap_bram_oarg_101_din1),
        .ap_bram_101_dout1(ap_bram_oarg_101_dout1),
        .ap_bram_101_we1(ap_bram_oarg_101_we1),
        .ap_bram_101_en1(ap_bram_oarg_101_en1),
        .m_axis_bram_102_aclk(m_axis_bram_102_aclk),
        .m_axis_bram_102_aresetn(m_axis_bram_102_aresetn),
        .m_axis_bram_102_tlast(m_axis_bram_102_tlast),
        .m_axis_bram_102_tvalid(m_axis_bram_102_tvalid),
        .m_axis_bram_102_tkeep(m_axis_bram_102_tkeep),
        .m_axis_bram_102_tstrb(m_axis_bram_102_tstrb),
        .m_axis_bram_102_tdata(m_axis_bram_102_tdata),
        .m_axis_bram_102_tready(m_axis_bram_102_tready),
        .ap_bram_102_addr0(ap_bram_oarg_102_addr0),
        .ap_bram_102_din0(ap_bram_oarg_102_din0),
        .ap_bram_102_dout0(ap_bram_oarg_102_dout0),
        .ap_bram_102_we0(ap_bram_oarg_102_we0),
        .ap_bram_102_en0(ap_bram_oarg_102_en0),
        .ap_bram_102_addr1(ap_bram_oarg_102_addr1),
        .ap_bram_102_din1(ap_bram_oarg_102_din1),
        .ap_bram_102_dout1(ap_bram_oarg_102_dout1),
        .ap_bram_102_we1(ap_bram_oarg_102_we1),
        .ap_bram_102_en1(ap_bram_oarg_102_en1),
        .m_axis_bram_103_aclk(m_axis_bram_103_aclk),
        .m_axis_bram_103_aresetn(m_axis_bram_103_aresetn),
        .m_axis_bram_103_tlast(m_axis_bram_103_tlast),
        .m_axis_bram_103_tvalid(m_axis_bram_103_tvalid),
        .m_axis_bram_103_tkeep(m_axis_bram_103_tkeep),
        .m_axis_bram_103_tstrb(m_axis_bram_103_tstrb),
        .m_axis_bram_103_tdata(m_axis_bram_103_tdata),
        .m_axis_bram_103_tready(m_axis_bram_103_tready),
        .ap_bram_103_addr0(ap_bram_oarg_103_addr0),
        .ap_bram_103_din0(ap_bram_oarg_103_din0),
        .ap_bram_103_dout0(ap_bram_oarg_103_dout0),
        .ap_bram_103_we0(ap_bram_oarg_103_we0),
        .ap_bram_103_en0(ap_bram_oarg_103_en0),
        .ap_bram_103_addr1(ap_bram_oarg_103_addr1),
        .ap_bram_103_din1(ap_bram_oarg_103_din1),
        .ap_bram_103_dout1(ap_bram_oarg_103_dout1),
        .ap_bram_103_we1(ap_bram_oarg_103_we1),
        .ap_bram_103_en1(ap_bram_oarg_103_en1),
        .m_axis_bram_104_aclk(m_axis_bram_104_aclk),
        .m_axis_bram_104_aresetn(m_axis_bram_104_aresetn),
        .m_axis_bram_104_tlast(m_axis_bram_104_tlast),
        .m_axis_bram_104_tvalid(m_axis_bram_104_tvalid),
        .m_axis_bram_104_tkeep(m_axis_bram_104_tkeep),
        .m_axis_bram_104_tstrb(m_axis_bram_104_tstrb),
        .m_axis_bram_104_tdata(m_axis_bram_104_tdata),
        .m_axis_bram_104_tready(m_axis_bram_104_tready),
        .ap_bram_104_addr0(ap_bram_oarg_104_addr0),
        .ap_bram_104_din0(ap_bram_oarg_104_din0),
        .ap_bram_104_dout0(ap_bram_oarg_104_dout0),
        .ap_bram_104_we0(ap_bram_oarg_104_we0),
        .ap_bram_104_en0(ap_bram_oarg_104_en0),
        .ap_bram_104_addr1(ap_bram_oarg_104_addr1),
        .ap_bram_104_din1(ap_bram_oarg_104_din1),
        .ap_bram_104_dout1(ap_bram_oarg_104_dout1),
        .ap_bram_104_we1(ap_bram_oarg_104_we1),
        .ap_bram_104_en1(ap_bram_oarg_104_en1),
        .m_axis_bram_105_aclk(m_axis_bram_105_aclk),
        .m_axis_bram_105_aresetn(m_axis_bram_105_aresetn),
        .m_axis_bram_105_tlast(m_axis_bram_105_tlast),
        .m_axis_bram_105_tvalid(m_axis_bram_105_tvalid),
        .m_axis_bram_105_tkeep(m_axis_bram_105_tkeep),
        .m_axis_bram_105_tstrb(m_axis_bram_105_tstrb),
        .m_axis_bram_105_tdata(m_axis_bram_105_tdata),
        .m_axis_bram_105_tready(m_axis_bram_105_tready),
        .ap_bram_105_addr0(ap_bram_oarg_105_addr0),
        .ap_bram_105_din0(ap_bram_oarg_105_din0),
        .ap_bram_105_dout0(ap_bram_oarg_105_dout0),
        .ap_bram_105_we0(ap_bram_oarg_105_we0),
        .ap_bram_105_en0(ap_bram_oarg_105_en0),
        .ap_bram_105_addr1(ap_bram_oarg_105_addr1),
        .ap_bram_105_din1(ap_bram_oarg_105_din1),
        .ap_bram_105_dout1(ap_bram_oarg_105_dout1),
        .ap_bram_105_we1(ap_bram_oarg_105_we1),
        .ap_bram_105_en1(ap_bram_oarg_105_en1),
        .m_axis_bram_106_aclk(m_axis_bram_106_aclk),
        .m_axis_bram_106_aresetn(m_axis_bram_106_aresetn),
        .m_axis_bram_106_tlast(m_axis_bram_106_tlast),
        .m_axis_bram_106_tvalid(m_axis_bram_106_tvalid),
        .m_axis_bram_106_tkeep(m_axis_bram_106_tkeep),
        .m_axis_bram_106_tstrb(m_axis_bram_106_tstrb),
        .m_axis_bram_106_tdata(m_axis_bram_106_tdata),
        .m_axis_bram_106_tready(m_axis_bram_106_tready),
        .ap_bram_106_addr0(ap_bram_oarg_106_addr0),
        .ap_bram_106_din0(ap_bram_oarg_106_din0),
        .ap_bram_106_dout0(ap_bram_oarg_106_dout0),
        .ap_bram_106_we0(ap_bram_oarg_106_we0),
        .ap_bram_106_en0(ap_bram_oarg_106_en0),
        .ap_bram_106_addr1(ap_bram_oarg_106_addr1),
        .ap_bram_106_din1(ap_bram_oarg_106_din1),
        .ap_bram_106_dout1(ap_bram_oarg_106_dout1),
        .ap_bram_106_we1(ap_bram_oarg_106_we1),
        .ap_bram_106_en1(ap_bram_oarg_106_en1),
        .m_axis_bram_107_aclk(m_axis_bram_107_aclk),
        .m_axis_bram_107_aresetn(m_axis_bram_107_aresetn),
        .m_axis_bram_107_tlast(m_axis_bram_107_tlast),
        .m_axis_bram_107_tvalid(m_axis_bram_107_tvalid),
        .m_axis_bram_107_tkeep(m_axis_bram_107_tkeep),
        .m_axis_bram_107_tstrb(m_axis_bram_107_tstrb),
        .m_axis_bram_107_tdata(m_axis_bram_107_tdata),
        .m_axis_bram_107_tready(m_axis_bram_107_tready),
        .ap_bram_107_addr0(ap_bram_oarg_107_addr0),
        .ap_bram_107_din0(ap_bram_oarg_107_din0),
        .ap_bram_107_dout0(ap_bram_oarg_107_dout0),
        .ap_bram_107_we0(ap_bram_oarg_107_we0),
        .ap_bram_107_en0(ap_bram_oarg_107_en0),
        .ap_bram_107_addr1(ap_bram_oarg_107_addr1),
        .ap_bram_107_din1(ap_bram_oarg_107_din1),
        .ap_bram_107_dout1(ap_bram_oarg_107_dout1),
        .ap_bram_107_we1(ap_bram_oarg_107_we1),
        .ap_bram_107_en1(ap_bram_oarg_107_en1),
        .m_axis_bram_108_aclk(m_axis_bram_108_aclk),
        .m_axis_bram_108_aresetn(m_axis_bram_108_aresetn),
        .m_axis_bram_108_tlast(m_axis_bram_108_tlast),
        .m_axis_bram_108_tvalid(m_axis_bram_108_tvalid),
        .m_axis_bram_108_tkeep(m_axis_bram_108_tkeep),
        .m_axis_bram_108_tstrb(m_axis_bram_108_tstrb),
        .m_axis_bram_108_tdata(m_axis_bram_108_tdata),
        .m_axis_bram_108_tready(m_axis_bram_108_tready),
        .ap_bram_108_addr0(ap_bram_oarg_108_addr0),
        .ap_bram_108_din0(ap_bram_oarg_108_din0),
        .ap_bram_108_dout0(ap_bram_oarg_108_dout0),
        .ap_bram_108_we0(ap_bram_oarg_108_we0),
        .ap_bram_108_en0(ap_bram_oarg_108_en0),
        .ap_bram_108_addr1(ap_bram_oarg_108_addr1),
        .ap_bram_108_din1(ap_bram_oarg_108_din1),
        .ap_bram_108_dout1(ap_bram_oarg_108_dout1),
        .ap_bram_108_we1(ap_bram_oarg_108_we1),
        .ap_bram_108_en1(ap_bram_oarg_108_en1),
        .m_axis_bram_109_aclk(m_axis_bram_109_aclk),
        .m_axis_bram_109_aresetn(m_axis_bram_109_aresetn),
        .m_axis_bram_109_tlast(m_axis_bram_109_tlast),
        .m_axis_bram_109_tvalid(m_axis_bram_109_tvalid),
        .m_axis_bram_109_tkeep(m_axis_bram_109_tkeep),
        .m_axis_bram_109_tstrb(m_axis_bram_109_tstrb),
        .m_axis_bram_109_tdata(m_axis_bram_109_tdata),
        .m_axis_bram_109_tready(m_axis_bram_109_tready),
        .ap_bram_109_addr0(ap_bram_oarg_109_addr0),
        .ap_bram_109_din0(ap_bram_oarg_109_din0),
        .ap_bram_109_dout0(ap_bram_oarg_109_dout0),
        .ap_bram_109_we0(ap_bram_oarg_109_we0),
        .ap_bram_109_en0(ap_bram_oarg_109_en0),
        .ap_bram_109_addr1(ap_bram_oarg_109_addr1),
        .ap_bram_109_din1(ap_bram_oarg_109_din1),
        .ap_bram_109_dout1(ap_bram_oarg_109_dout1),
        .ap_bram_109_we1(ap_bram_oarg_109_we1),
        .ap_bram_109_en1(ap_bram_oarg_109_en1),
        .m_axis_bram_110_aclk(m_axis_bram_110_aclk),
        .m_axis_bram_110_aresetn(m_axis_bram_110_aresetn),
        .m_axis_bram_110_tlast(m_axis_bram_110_tlast),
        .m_axis_bram_110_tvalid(m_axis_bram_110_tvalid),
        .m_axis_bram_110_tkeep(m_axis_bram_110_tkeep),
        .m_axis_bram_110_tstrb(m_axis_bram_110_tstrb),
        .m_axis_bram_110_tdata(m_axis_bram_110_tdata),
        .m_axis_bram_110_tready(m_axis_bram_110_tready),
        .ap_bram_110_addr0(ap_bram_oarg_110_addr0),
        .ap_bram_110_din0(ap_bram_oarg_110_din0),
        .ap_bram_110_dout0(ap_bram_oarg_110_dout0),
        .ap_bram_110_we0(ap_bram_oarg_110_we0),
        .ap_bram_110_en0(ap_bram_oarg_110_en0),
        .ap_bram_110_addr1(ap_bram_oarg_110_addr1),
        .ap_bram_110_din1(ap_bram_oarg_110_din1),
        .ap_bram_110_dout1(ap_bram_oarg_110_dout1),
        .ap_bram_110_we1(ap_bram_oarg_110_we1),
        .ap_bram_110_en1(ap_bram_oarg_110_en1),
        .m_axis_bram_111_aclk(m_axis_bram_111_aclk),
        .m_axis_bram_111_aresetn(m_axis_bram_111_aresetn),
        .m_axis_bram_111_tlast(m_axis_bram_111_tlast),
        .m_axis_bram_111_tvalid(m_axis_bram_111_tvalid),
        .m_axis_bram_111_tkeep(m_axis_bram_111_tkeep),
        .m_axis_bram_111_tstrb(m_axis_bram_111_tstrb),
        .m_axis_bram_111_tdata(m_axis_bram_111_tdata),
        .m_axis_bram_111_tready(m_axis_bram_111_tready),
        .ap_bram_111_addr0(ap_bram_oarg_111_addr0),
        .ap_bram_111_din0(ap_bram_oarg_111_din0),
        .ap_bram_111_dout0(ap_bram_oarg_111_dout0),
        .ap_bram_111_we0(ap_bram_oarg_111_we0),
        .ap_bram_111_en0(ap_bram_oarg_111_en0),
        .ap_bram_111_addr1(ap_bram_oarg_111_addr1),
        .ap_bram_111_din1(ap_bram_oarg_111_din1),
        .ap_bram_111_dout1(ap_bram_oarg_111_dout1),
        .ap_bram_111_we1(ap_bram_oarg_111_we1),
        .ap_bram_111_en1(ap_bram_oarg_111_en1),
        .m_axis_bram_112_aclk(m_axis_bram_112_aclk),
        .m_axis_bram_112_aresetn(m_axis_bram_112_aresetn),
        .m_axis_bram_112_tlast(m_axis_bram_112_tlast),
        .m_axis_bram_112_tvalid(m_axis_bram_112_tvalid),
        .m_axis_bram_112_tkeep(m_axis_bram_112_tkeep),
        .m_axis_bram_112_tstrb(m_axis_bram_112_tstrb),
        .m_axis_bram_112_tdata(m_axis_bram_112_tdata),
        .m_axis_bram_112_tready(m_axis_bram_112_tready),
        .ap_bram_112_addr0(ap_bram_oarg_112_addr0),
        .ap_bram_112_din0(ap_bram_oarg_112_din0),
        .ap_bram_112_dout0(ap_bram_oarg_112_dout0),
        .ap_bram_112_we0(ap_bram_oarg_112_we0),
        .ap_bram_112_en0(ap_bram_oarg_112_en0),
        .ap_bram_112_addr1(ap_bram_oarg_112_addr1),
        .ap_bram_112_din1(ap_bram_oarg_112_din1),
        .ap_bram_112_dout1(ap_bram_oarg_112_dout1),
        .ap_bram_112_we1(ap_bram_oarg_112_we1),
        .ap_bram_112_en1(ap_bram_oarg_112_en1),
        .m_axis_bram_113_aclk(m_axis_bram_113_aclk),
        .m_axis_bram_113_aresetn(m_axis_bram_113_aresetn),
        .m_axis_bram_113_tlast(m_axis_bram_113_tlast),
        .m_axis_bram_113_tvalid(m_axis_bram_113_tvalid),
        .m_axis_bram_113_tkeep(m_axis_bram_113_tkeep),
        .m_axis_bram_113_tstrb(m_axis_bram_113_tstrb),
        .m_axis_bram_113_tdata(m_axis_bram_113_tdata),
        .m_axis_bram_113_tready(m_axis_bram_113_tready),
        .ap_bram_113_addr0(ap_bram_oarg_113_addr0),
        .ap_bram_113_din0(ap_bram_oarg_113_din0),
        .ap_bram_113_dout0(ap_bram_oarg_113_dout0),
        .ap_bram_113_we0(ap_bram_oarg_113_we0),
        .ap_bram_113_en0(ap_bram_oarg_113_en0),
        .ap_bram_113_addr1(ap_bram_oarg_113_addr1),
        .ap_bram_113_din1(ap_bram_oarg_113_din1),
        .ap_bram_113_dout1(ap_bram_oarg_113_dout1),
        .ap_bram_113_we1(ap_bram_oarg_113_we1),
        .ap_bram_113_en1(ap_bram_oarg_113_en1),
        .m_axis_bram_114_aclk(m_axis_bram_114_aclk),
        .m_axis_bram_114_aresetn(m_axis_bram_114_aresetn),
        .m_axis_bram_114_tlast(m_axis_bram_114_tlast),
        .m_axis_bram_114_tvalid(m_axis_bram_114_tvalid),
        .m_axis_bram_114_tkeep(m_axis_bram_114_tkeep),
        .m_axis_bram_114_tstrb(m_axis_bram_114_tstrb),
        .m_axis_bram_114_tdata(m_axis_bram_114_tdata),
        .m_axis_bram_114_tready(m_axis_bram_114_tready),
        .ap_bram_114_addr0(ap_bram_oarg_114_addr0),
        .ap_bram_114_din0(ap_bram_oarg_114_din0),
        .ap_bram_114_dout0(ap_bram_oarg_114_dout0),
        .ap_bram_114_we0(ap_bram_oarg_114_we0),
        .ap_bram_114_en0(ap_bram_oarg_114_en0),
        .ap_bram_114_addr1(ap_bram_oarg_114_addr1),
        .ap_bram_114_din1(ap_bram_oarg_114_din1),
        .ap_bram_114_dout1(ap_bram_oarg_114_dout1),
        .ap_bram_114_we1(ap_bram_oarg_114_we1),
        .ap_bram_114_en1(ap_bram_oarg_114_en1),
        .m_axis_bram_115_aclk(m_axis_bram_115_aclk),
        .m_axis_bram_115_aresetn(m_axis_bram_115_aresetn),
        .m_axis_bram_115_tlast(m_axis_bram_115_tlast),
        .m_axis_bram_115_tvalid(m_axis_bram_115_tvalid),
        .m_axis_bram_115_tkeep(m_axis_bram_115_tkeep),
        .m_axis_bram_115_tstrb(m_axis_bram_115_tstrb),
        .m_axis_bram_115_tdata(m_axis_bram_115_tdata),
        .m_axis_bram_115_tready(m_axis_bram_115_tready),
        .ap_bram_115_addr0(ap_bram_oarg_115_addr0),
        .ap_bram_115_din0(ap_bram_oarg_115_din0),
        .ap_bram_115_dout0(ap_bram_oarg_115_dout0),
        .ap_bram_115_we0(ap_bram_oarg_115_we0),
        .ap_bram_115_en0(ap_bram_oarg_115_en0),
        .ap_bram_115_addr1(ap_bram_oarg_115_addr1),
        .ap_bram_115_din1(ap_bram_oarg_115_din1),
        .ap_bram_115_dout1(ap_bram_oarg_115_dout1),
        .ap_bram_115_we1(ap_bram_oarg_115_we1),
        .ap_bram_115_en1(ap_bram_oarg_115_en1),
        .m_axis_bram_116_aclk(m_axis_bram_116_aclk),
        .m_axis_bram_116_aresetn(m_axis_bram_116_aresetn),
        .m_axis_bram_116_tlast(m_axis_bram_116_tlast),
        .m_axis_bram_116_tvalid(m_axis_bram_116_tvalid),
        .m_axis_bram_116_tkeep(m_axis_bram_116_tkeep),
        .m_axis_bram_116_tstrb(m_axis_bram_116_tstrb),
        .m_axis_bram_116_tdata(m_axis_bram_116_tdata),
        .m_axis_bram_116_tready(m_axis_bram_116_tready),
        .ap_bram_116_addr0(ap_bram_oarg_116_addr0),
        .ap_bram_116_din0(ap_bram_oarg_116_din0),
        .ap_bram_116_dout0(ap_bram_oarg_116_dout0),
        .ap_bram_116_we0(ap_bram_oarg_116_we0),
        .ap_bram_116_en0(ap_bram_oarg_116_en0),
        .ap_bram_116_addr1(ap_bram_oarg_116_addr1),
        .ap_bram_116_din1(ap_bram_oarg_116_din1),
        .ap_bram_116_dout1(ap_bram_oarg_116_dout1),
        .ap_bram_116_we1(ap_bram_oarg_116_we1),
        .ap_bram_116_en1(ap_bram_oarg_116_en1),
        .m_axis_bram_117_aclk(m_axis_bram_117_aclk),
        .m_axis_bram_117_aresetn(m_axis_bram_117_aresetn),
        .m_axis_bram_117_tlast(m_axis_bram_117_tlast),
        .m_axis_bram_117_tvalid(m_axis_bram_117_tvalid),
        .m_axis_bram_117_tkeep(m_axis_bram_117_tkeep),
        .m_axis_bram_117_tstrb(m_axis_bram_117_tstrb),
        .m_axis_bram_117_tdata(m_axis_bram_117_tdata),
        .m_axis_bram_117_tready(m_axis_bram_117_tready),
        .ap_bram_117_addr0(ap_bram_oarg_117_addr0),
        .ap_bram_117_din0(ap_bram_oarg_117_din0),
        .ap_bram_117_dout0(ap_bram_oarg_117_dout0),
        .ap_bram_117_we0(ap_bram_oarg_117_we0),
        .ap_bram_117_en0(ap_bram_oarg_117_en0),
        .ap_bram_117_addr1(ap_bram_oarg_117_addr1),
        .ap_bram_117_din1(ap_bram_oarg_117_din1),
        .ap_bram_117_dout1(ap_bram_oarg_117_dout1),
        .ap_bram_117_we1(ap_bram_oarg_117_we1),
        .ap_bram_117_en1(ap_bram_oarg_117_en1),
        .m_axis_bram_118_aclk(m_axis_bram_118_aclk),
        .m_axis_bram_118_aresetn(m_axis_bram_118_aresetn),
        .m_axis_bram_118_tlast(m_axis_bram_118_tlast),
        .m_axis_bram_118_tvalid(m_axis_bram_118_tvalid),
        .m_axis_bram_118_tkeep(m_axis_bram_118_tkeep),
        .m_axis_bram_118_tstrb(m_axis_bram_118_tstrb),
        .m_axis_bram_118_tdata(m_axis_bram_118_tdata),
        .m_axis_bram_118_tready(m_axis_bram_118_tready),
        .ap_bram_118_addr0(ap_bram_oarg_118_addr0),
        .ap_bram_118_din0(ap_bram_oarg_118_din0),
        .ap_bram_118_dout0(ap_bram_oarg_118_dout0),
        .ap_bram_118_we0(ap_bram_oarg_118_we0),
        .ap_bram_118_en0(ap_bram_oarg_118_en0),
        .ap_bram_118_addr1(ap_bram_oarg_118_addr1),
        .ap_bram_118_din1(ap_bram_oarg_118_din1),
        .ap_bram_118_dout1(ap_bram_oarg_118_dout1),
        .ap_bram_118_we1(ap_bram_oarg_118_we1),
        .ap_bram_118_en1(ap_bram_oarg_118_en1),
        .m_axis_bram_119_aclk(m_axis_bram_119_aclk),
        .m_axis_bram_119_aresetn(m_axis_bram_119_aresetn),
        .m_axis_bram_119_tlast(m_axis_bram_119_tlast),
        .m_axis_bram_119_tvalid(m_axis_bram_119_tvalid),
        .m_axis_bram_119_tkeep(m_axis_bram_119_tkeep),
        .m_axis_bram_119_tstrb(m_axis_bram_119_tstrb),
        .m_axis_bram_119_tdata(m_axis_bram_119_tdata),
        .m_axis_bram_119_tready(m_axis_bram_119_tready),
        .ap_bram_119_addr0(ap_bram_oarg_119_addr0),
        .ap_bram_119_din0(ap_bram_oarg_119_din0),
        .ap_bram_119_dout0(ap_bram_oarg_119_dout0),
        .ap_bram_119_we0(ap_bram_oarg_119_we0),
        .ap_bram_119_en0(ap_bram_oarg_119_en0),
        .ap_bram_119_addr1(ap_bram_oarg_119_addr1),
        .ap_bram_119_din1(ap_bram_oarg_119_din1),
        .ap_bram_119_dout1(ap_bram_oarg_119_dout1),
        .ap_bram_119_we1(ap_bram_oarg_119_we1),
        .ap_bram_119_en1(ap_bram_oarg_119_en1),
        .m_axis_bram_120_aclk(m_axis_bram_120_aclk),
        .m_axis_bram_120_aresetn(m_axis_bram_120_aresetn),
        .m_axis_bram_120_tlast(m_axis_bram_120_tlast),
        .m_axis_bram_120_tvalid(m_axis_bram_120_tvalid),
        .m_axis_bram_120_tkeep(m_axis_bram_120_tkeep),
        .m_axis_bram_120_tstrb(m_axis_bram_120_tstrb),
        .m_axis_bram_120_tdata(m_axis_bram_120_tdata),
        .m_axis_bram_120_tready(m_axis_bram_120_tready),
        .ap_bram_120_addr0(ap_bram_oarg_120_addr0),
        .ap_bram_120_din0(ap_bram_oarg_120_din0),
        .ap_bram_120_dout0(ap_bram_oarg_120_dout0),
        .ap_bram_120_we0(ap_bram_oarg_120_we0),
        .ap_bram_120_en0(ap_bram_oarg_120_en0),
        .ap_bram_120_addr1(ap_bram_oarg_120_addr1),
        .ap_bram_120_din1(ap_bram_oarg_120_din1),
        .ap_bram_120_dout1(ap_bram_oarg_120_dout1),
        .ap_bram_120_we1(ap_bram_oarg_120_we1),
        .ap_bram_120_en1(ap_bram_oarg_120_en1),
        .m_axis_bram_121_aclk(m_axis_bram_121_aclk),
        .m_axis_bram_121_aresetn(m_axis_bram_121_aresetn),
        .m_axis_bram_121_tlast(m_axis_bram_121_tlast),
        .m_axis_bram_121_tvalid(m_axis_bram_121_tvalid),
        .m_axis_bram_121_tkeep(m_axis_bram_121_tkeep),
        .m_axis_bram_121_tstrb(m_axis_bram_121_tstrb),
        .m_axis_bram_121_tdata(m_axis_bram_121_tdata),
        .m_axis_bram_121_tready(m_axis_bram_121_tready),
        .ap_bram_121_addr0(ap_bram_oarg_121_addr0),
        .ap_bram_121_din0(ap_bram_oarg_121_din0),
        .ap_bram_121_dout0(ap_bram_oarg_121_dout0),
        .ap_bram_121_we0(ap_bram_oarg_121_we0),
        .ap_bram_121_en0(ap_bram_oarg_121_en0),
        .ap_bram_121_addr1(ap_bram_oarg_121_addr1),
        .ap_bram_121_din1(ap_bram_oarg_121_din1),
        .ap_bram_121_dout1(ap_bram_oarg_121_dout1),
        .ap_bram_121_we1(ap_bram_oarg_121_we1),
        .ap_bram_121_en1(ap_bram_oarg_121_en1),
        .m_axis_bram_122_aclk(m_axis_bram_122_aclk),
        .m_axis_bram_122_aresetn(m_axis_bram_122_aresetn),
        .m_axis_bram_122_tlast(m_axis_bram_122_tlast),
        .m_axis_bram_122_tvalid(m_axis_bram_122_tvalid),
        .m_axis_bram_122_tkeep(m_axis_bram_122_tkeep),
        .m_axis_bram_122_tstrb(m_axis_bram_122_tstrb),
        .m_axis_bram_122_tdata(m_axis_bram_122_tdata),
        .m_axis_bram_122_tready(m_axis_bram_122_tready),
        .ap_bram_122_addr0(ap_bram_oarg_122_addr0),
        .ap_bram_122_din0(ap_bram_oarg_122_din0),
        .ap_bram_122_dout0(ap_bram_oarg_122_dout0),
        .ap_bram_122_we0(ap_bram_oarg_122_we0),
        .ap_bram_122_en0(ap_bram_oarg_122_en0),
        .ap_bram_122_addr1(ap_bram_oarg_122_addr1),
        .ap_bram_122_din1(ap_bram_oarg_122_din1),
        .ap_bram_122_dout1(ap_bram_oarg_122_dout1),
        .ap_bram_122_we1(ap_bram_oarg_122_we1),
        .ap_bram_122_en1(ap_bram_oarg_122_en1),
        .m_axis_bram_123_aclk(m_axis_bram_123_aclk),
        .m_axis_bram_123_aresetn(m_axis_bram_123_aresetn),
        .m_axis_bram_123_tlast(m_axis_bram_123_tlast),
        .m_axis_bram_123_tvalid(m_axis_bram_123_tvalid),
        .m_axis_bram_123_tkeep(m_axis_bram_123_tkeep),
        .m_axis_bram_123_tstrb(m_axis_bram_123_tstrb),
        .m_axis_bram_123_tdata(m_axis_bram_123_tdata),
        .m_axis_bram_123_tready(m_axis_bram_123_tready),
        .ap_bram_123_addr0(ap_bram_oarg_123_addr0),
        .ap_bram_123_din0(ap_bram_oarg_123_din0),
        .ap_bram_123_dout0(ap_bram_oarg_123_dout0),
        .ap_bram_123_we0(ap_bram_oarg_123_we0),
        .ap_bram_123_en0(ap_bram_oarg_123_en0),
        .ap_bram_123_addr1(ap_bram_oarg_123_addr1),
        .ap_bram_123_din1(ap_bram_oarg_123_din1),
        .ap_bram_123_dout1(ap_bram_oarg_123_dout1),
        .ap_bram_123_we1(ap_bram_oarg_123_we1),
        .ap_bram_123_en1(ap_bram_oarg_123_en1),
        .m_axis_bram_124_aclk(m_axis_bram_124_aclk),
        .m_axis_bram_124_aresetn(m_axis_bram_124_aresetn),
        .m_axis_bram_124_tlast(m_axis_bram_124_tlast),
        .m_axis_bram_124_tvalid(m_axis_bram_124_tvalid),
        .m_axis_bram_124_tkeep(m_axis_bram_124_tkeep),
        .m_axis_bram_124_tstrb(m_axis_bram_124_tstrb),
        .m_axis_bram_124_tdata(m_axis_bram_124_tdata),
        .m_axis_bram_124_tready(m_axis_bram_124_tready),
        .ap_bram_124_addr0(ap_bram_oarg_124_addr0),
        .ap_bram_124_din0(ap_bram_oarg_124_din0),
        .ap_bram_124_dout0(ap_bram_oarg_124_dout0),
        .ap_bram_124_we0(ap_bram_oarg_124_we0),
        .ap_bram_124_en0(ap_bram_oarg_124_en0),
        .ap_bram_124_addr1(ap_bram_oarg_124_addr1),
        .ap_bram_124_din1(ap_bram_oarg_124_din1),
        .ap_bram_124_dout1(ap_bram_oarg_124_dout1),
        .ap_bram_124_we1(ap_bram_oarg_124_we1),
        .ap_bram_124_en1(ap_bram_oarg_124_en1),
        .m_axis_bram_125_aclk(m_axis_bram_125_aclk),
        .m_axis_bram_125_aresetn(m_axis_bram_125_aresetn),
        .m_axis_bram_125_tlast(m_axis_bram_125_tlast),
        .m_axis_bram_125_tvalid(m_axis_bram_125_tvalid),
        .m_axis_bram_125_tkeep(m_axis_bram_125_tkeep),
        .m_axis_bram_125_tstrb(m_axis_bram_125_tstrb),
        .m_axis_bram_125_tdata(m_axis_bram_125_tdata),
        .m_axis_bram_125_tready(m_axis_bram_125_tready),
        .ap_bram_125_addr0(ap_bram_oarg_125_addr0),
        .ap_bram_125_din0(ap_bram_oarg_125_din0),
        .ap_bram_125_dout0(ap_bram_oarg_125_dout0),
        .ap_bram_125_we0(ap_bram_oarg_125_we0),
        .ap_bram_125_en0(ap_bram_oarg_125_en0),
        .ap_bram_125_addr1(ap_bram_oarg_125_addr1),
        .ap_bram_125_din1(ap_bram_oarg_125_din1),
        .ap_bram_125_dout1(ap_bram_oarg_125_dout1),
        .ap_bram_125_we1(ap_bram_oarg_125_we1),
        .ap_bram_125_en1(ap_bram_oarg_125_en1),
        .m_axis_bram_126_aclk(m_axis_bram_126_aclk),
        .m_axis_bram_126_aresetn(m_axis_bram_126_aresetn),
        .m_axis_bram_126_tlast(m_axis_bram_126_tlast),
        .m_axis_bram_126_tvalid(m_axis_bram_126_tvalid),
        .m_axis_bram_126_tkeep(m_axis_bram_126_tkeep),
        .m_axis_bram_126_tstrb(m_axis_bram_126_tstrb),
        .m_axis_bram_126_tdata(m_axis_bram_126_tdata),
        .m_axis_bram_126_tready(m_axis_bram_126_tready),
        .ap_bram_126_addr0(ap_bram_oarg_126_addr0),
        .ap_bram_126_din0(ap_bram_oarg_126_din0),
        .ap_bram_126_dout0(ap_bram_oarg_126_dout0),
        .ap_bram_126_we0(ap_bram_oarg_126_we0),
        .ap_bram_126_en0(ap_bram_oarg_126_en0),
        .ap_bram_126_addr1(ap_bram_oarg_126_addr1),
        .ap_bram_126_din1(ap_bram_oarg_126_din1),
        .ap_bram_126_dout1(ap_bram_oarg_126_dout1),
        .ap_bram_126_we1(ap_bram_oarg_126_we1),
        .ap_bram_126_en1(ap_bram_oarg_126_en1),
        .m_axis_bram_127_aclk(m_axis_bram_127_aclk),
        .m_axis_bram_127_aresetn(m_axis_bram_127_aresetn),
        .m_axis_bram_127_tlast(m_axis_bram_127_tlast),
        .m_axis_bram_127_tvalid(m_axis_bram_127_tvalid),
        .m_axis_bram_127_tkeep(m_axis_bram_127_tkeep),
        .m_axis_bram_127_tstrb(m_axis_bram_127_tstrb),
        .m_axis_bram_127_tdata(m_axis_bram_127_tdata),
        .m_axis_bram_127_tready(m_axis_bram_127_tready),
        .ap_bram_127_addr0(ap_bram_oarg_127_addr0),
        .ap_bram_127_din0(ap_bram_oarg_127_din0),
        .ap_bram_127_dout0(ap_bram_oarg_127_dout0),
        .ap_bram_127_we0(ap_bram_oarg_127_we0),
        .ap_bram_127_en0(ap_bram_oarg_127_en0),
        .ap_bram_127_addr1(ap_bram_oarg_127_addr1),
        .ap_bram_127_din1(ap_bram_oarg_127_din1),
        .ap_bram_127_dout1(ap_bram_oarg_127_dout1),
        .ap_bram_127_we1(ap_bram_oarg_127_we1),
        .ap_bram_127_en1(ap_bram_oarg_127_en1)
    );

endmodule
