// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689
`timescale 1ns / 1ps

module aximm_args #(
    parameter C_NUM_AXIMMs = 0,
    parameter M_AXIMM_ADDR_WIDTH = 32,
    parameter M_AXIMM_0_DATA_WIDTH = 32,
    parameter M_AXIMM_1_DATA_WIDTH = 32,
    parameter M_AXIMM_2_DATA_WIDTH = 32,
    parameter M_AXIMM_3_DATA_WIDTH = 32,
    parameter M_AXIMM_4_DATA_WIDTH = 32,
    parameter M_AXIMM_5_DATA_WIDTH = 32,
    parameter M_AXIMM_6_DATA_WIDTH = 32,
    parameter M_AXIMM_7_DATA_WIDTH = 32,
    parameter M_AXIMM_8_DATA_WIDTH = 32,
    parameter M_AXIMM_9_DATA_WIDTH = 32,
    parameter M_AXIMM_10_DATA_WIDTH = 32,
    parameter M_AXIMM_11_DATA_WIDTH = 32,
    parameter M_AXIMM_12_DATA_WIDTH = 32,
    parameter M_AXIMM_13_DATA_WIDTH = 32,
    parameter M_AXIMM_14_DATA_WIDTH = 32,
    parameter M_AXIMM_15_DATA_WIDTH = 32,
    parameter M_AXIMM_16_DATA_WIDTH = 32,
    parameter M_AXIMM_17_DATA_WIDTH = 32,
    parameter M_AXIMM_18_DATA_WIDTH = 32,
    parameter M_AXIMM_19_DATA_WIDTH = 32,
    parameter M_AXIMM_20_DATA_WIDTH = 32,
    parameter M_AXIMM_21_DATA_WIDTH = 32,
    parameter M_AXIMM_22_DATA_WIDTH = 32,
    parameter M_AXIMM_23_DATA_WIDTH = 32,
    parameter M_AXIMM_24_DATA_WIDTH = 32,
    parameter M_AXIMM_25_DATA_WIDTH = 32,
    parameter M_AXIMM_26_DATA_WIDTH = 32,
    parameter M_AXIMM_27_DATA_WIDTH = 32,
    parameter M_AXIMM_28_DATA_WIDTH = 32,
    parameter M_AXIMM_29_DATA_WIDTH = 32,
    parameter M_AXIMM_30_DATA_WIDTH = 32,
    parameter M_AXIMM_31_DATA_WIDTH = 32,
    parameter M_AXIMM_32_DATA_WIDTH = 32,
    parameter M_AXIMM_33_DATA_WIDTH = 32,
    parameter M_AXIMM_34_DATA_WIDTH = 32,
    parameter M_AXIMM_35_DATA_WIDTH = 32,
    parameter M_AXIMM_36_DATA_WIDTH = 32,
    parameter M_AXIMM_37_DATA_WIDTH = 32,
    parameter M_AXIMM_38_DATA_WIDTH = 32,
    parameter M_AXIMM_39_DATA_WIDTH = 32,
    parameter M_AXIMM_40_DATA_WIDTH = 32,
    parameter M_AXIMM_41_DATA_WIDTH = 32,
    parameter M_AXIMM_42_DATA_WIDTH = 32,
    parameter M_AXIMM_43_DATA_WIDTH = 32,
    parameter M_AXIMM_44_DATA_WIDTH = 32,
    parameter M_AXIMM_45_DATA_WIDTH = 32,
    parameter M_AXIMM_46_DATA_WIDTH = 32,
    parameter M_AXIMM_47_DATA_WIDTH = 32,
    parameter M_AXIMM_48_DATA_WIDTH = 32,
    parameter M_AXIMM_49_DATA_WIDTH = 32,
    parameter M_AXIMM_50_DATA_WIDTH = 32,
    parameter M_AXIMM_51_DATA_WIDTH = 32,
    parameter M_AXIMM_52_DATA_WIDTH = 32,
    parameter M_AXIMM_53_DATA_WIDTH = 32,
    parameter M_AXIMM_54_DATA_WIDTH = 32,
    parameter M_AXIMM_55_DATA_WIDTH = 32,
    parameter M_AXIMM_56_DATA_WIDTH = 32,
    parameter M_AXIMM_57_DATA_WIDTH = 32,
    parameter M_AXIMM_58_DATA_WIDTH = 32,
    parameter M_AXIMM_59_DATA_WIDTH = 32,
    parameter M_AXIMM_60_DATA_WIDTH = 32,
    parameter M_AXIMM_61_DATA_WIDTH = 32,
    parameter M_AXIMM_62_DATA_WIDTH = 32,
    parameter M_AXIMM_63_DATA_WIDTH = 32,
    parameter M_AXIMM_64_DATA_WIDTH = 32,
    parameter M_AXIMM_65_DATA_WIDTH = 32,
    parameter M_AXIMM_66_DATA_WIDTH = 32,
    parameter M_AXIMM_67_DATA_WIDTH = 32,
    parameter M_AXIMM_68_DATA_WIDTH = 32,
    parameter M_AXIMM_69_DATA_WIDTH = 32,
    parameter M_AXIMM_70_DATA_WIDTH = 32,
    parameter M_AXIMM_71_DATA_WIDTH = 32,
    parameter M_AXIMM_72_DATA_WIDTH = 32,
    parameter M_AXIMM_73_DATA_WIDTH = 32,
    parameter M_AXIMM_74_DATA_WIDTH = 32,
    parameter M_AXIMM_75_DATA_WIDTH = 32,
    parameter M_AXIMM_76_DATA_WIDTH = 32,
    parameter M_AXIMM_77_DATA_WIDTH = 32,
    parameter M_AXIMM_78_DATA_WIDTH = 32,
    parameter M_AXIMM_79_DATA_WIDTH = 32,
    parameter M_AXIMM_80_DATA_WIDTH = 32,
    parameter M_AXIMM_81_DATA_WIDTH = 32,
    parameter M_AXIMM_82_DATA_WIDTH = 32,
    parameter M_AXIMM_83_DATA_WIDTH = 32,
    parameter M_AXIMM_84_DATA_WIDTH = 32,
    parameter M_AXIMM_85_DATA_WIDTH = 32,
    parameter M_AXIMM_86_DATA_WIDTH = 32,
    parameter M_AXIMM_87_DATA_WIDTH = 32,
    parameter M_AXIMM_88_DATA_WIDTH = 32,
    parameter M_AXIMM_89_DATA_WIDTH = 32,
    parameter M_AXIMM_90_DATA_WIDTH = 32,
    parameter M_AXIMM_91_DATA_WIDTH = 32,
    parameter M_AXIMM_92_DATA_WIDTH = 32,
    parameter M_AXIMM_93_DATA_WIDTH = 32,
    parameter M_AXIMM_94_DATA_WIDTH = 32,
    parameter M_AXIMM_95_DATA_WIDTH = 32,
    parameter M_AXIMM_96_DATA_WIDTH = 32,
    parameter M_AXIMM_97_DATA_WIDTH = 32,
    parameter M_AXIMM_98_DATA_WIDTH = 32,
    parameter M_AXIMM_99_DATA_WIDTH = 32,
    parameter M_AXIMM_100_DATA_WIDTH = 32,
    parameter M_AXIMM_101_DATA_WIDTH = 32,
    parameter M_AXIMM_102_DATA_WIDTH = 32,
    parameter M_AXIMM_103_DATA_WIDTH = 32,
    parameter M_AXIMM_104_DATA_WIDTH = 32,
    parameter M_AXIMM_105_DATA_WIDTH = 32,
    parameter M_AXIMM_106_DATA_WIDTH = 32,
    parameter M_AXIMM_107_DATA_WIDTH = 32,
    parameter M_AXIMM_108_DATA_WIDTH = 32,
    parameter M_AXIMM_109_DATA_WIDTH = 32,
    parameter M_AXIMM_110_DATA_WIDTH = 32,
    parameter M_AXIMM_111_DATA_WIDTH = 32,
    parameter M_AXIMM_112_DATA_WIDTH = 32,
    parameter M_AXIMM_113_DATA_WIDTH = 32,
    parameter M_AXIMM_114_DATA_WIDTH = 32,
    parameter M_AXIMM_115_DATA_WIDTH = 32,
    parameter M_AXIMM_116_DATA_WIDTH = 32,
    parameter M_AXIMM_117_DATA_WIDTH = 32,
    parameter M_AXIMM_118_DATA_WIDTH = 32,
    parameter M_AXIMM_119_DATA_WIDTH = 32,
    parameter M_AXIMM_120_DATA_WIDTH = 32,
    parameter M_AXIMM_121_DATA_WIDTH = 32,
    parameter M_AXIMM_122_DATA_WIDTH = 32,
    parameter M_AXIMM_123_DATA_WIDTH = 32,
    parameter M_AXIMM_124_DATA_WIDTH = 32,
    parameter M_AXIMM_125_DATA_WIDTH = 32,
    parameter M_AXIMM_126_DATA_WIDTH = 32,
    parameter M_AXIMM_127_DATA_WIDTH = 32,
    parameter [0:0] M_AXIMM_0_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_ARUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_AWUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_BUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_RUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_WUSER_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_ARID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_AWID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_BID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_RID_WIDTH = 0,
    parameter [0:0] M_AXIMM_0_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_1_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_2_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_3_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_4_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_5_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_6_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_7_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_8_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_9_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_10_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_11_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_12_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_13_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_14_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_15_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_16_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_17_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_18_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_19_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_20_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_21_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_22_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_23_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_24_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_25_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_26_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_27_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_28_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_29_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_30_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_31_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_32_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_33_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_34_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_35_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_36_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_37_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_38_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_39_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_40_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_41_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_42_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_43_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_44_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_45_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_46_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_47_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_48_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_49_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_50_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_51_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_52_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_53_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_54_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_55_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_56_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_57_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_58_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_59_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_60_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_61_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_62_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_63_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_64_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_65_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_66_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_67_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_68_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_69_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_70_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_71_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_72_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_73_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_74_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_75_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_76_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_77_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_78_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_79_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_80_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_81_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_82_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_83_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_84_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_85_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_86_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_87_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_88_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_89_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_90_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_91_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_92_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_93_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_94_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_95_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_96_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_97_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_98_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_99_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_100_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_101_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_102_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_103_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_104_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_105_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_106_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_107_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_108_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_109_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_110_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_111_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_112_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_113_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_114_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_115_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_116_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_117_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_118_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_119_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_120_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_121_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_122_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_123_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_124_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_125_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_126_WID_WIDTH = 0,
    parameter [0:0] M_AXIMM_127_WID_WIDTH = 0
 ) (
    input acc_clk,
    input dm_clk,
    //control interface
    input aresetn,
    //AXI-MM pass-through interface 0
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_0_AWADDR,
    input wire [7:0]                      AP_AXIMM_0_AWLEN,
    input wire [2:0]                      AP_AXIMM_0_AWSIZE,
    input wire [1:0]                      AP_AXIMM_0_AWBURST,
    input wire [1:0]                      AP_AXIMM_0_AWLOCK,
    input wire [3:0]                      AP_AXIMM_0_AWCACHE,
    input wire [2:0]                      AP_AXIMM_0_AWPROT,
    input wire [3:0]                      AP_AXIMM_0_AWREGION,
    input wire [3:0]                      AP_AXIMM_0_AWQOS,
    input wire                            AP_AXIMM_0_AWVALID,
    output  wire                            AP_AXIMM_0_AWREADY,
    input wire [M_AXIMM_0_DATA_WIDTH-1:0]   AP_AXIMM_0_WDATA,
    input wire [M_AXIMM_0_DATA_WIDTH/8-1:0] AP_AXIMM_0_WSTRB,
    input wire                            AP_AXIMM_0_WLAST,
    input wire                            AP_AXIMM_0_WVALID,
    output  wire                            AP_AXIMM_0_WREADY,
    output  wire [1:0]                      AP_AXIMM_0_BRESP,
    output  wire                            AP_AXIMM_0_BVALID,
    input wire                            AP_AXIMM_0_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_0_ARADDR,
    input wire [7:0]                      AP_AXIMM_0_ARLEN,
    input wire [2:0]                      AP_AXIMM_0_ARSIZE,
    input wire [1:0]                      AP_AXIMM_0_ARBURST,
    input wire [1:0]                      AP_AXIMM_0_ARLOCK,
    input wire [3:0]                      AP_AXIMM_0_ARCACHE,
    input wire [2:0]                      AP_AXIMM_0_ARPROT,
    input wire [3:0]                      AP_AXIMM_0_ARREGION,
    input wire [3:0]                      AP_AXIMM_0_ARQOS,
    input wire                            AP_AXIMM_0_ARVALID,
    output  wire                            AP_AXIMM_0_ARREADY,
    output  wire [M_AXIMM_0_DATA_WIDTH-1:0]   AP_AXIMM_0_RDATA,
    output  wire [1:0]                      AP_AXIMM_0_RRESP,
    output  wire                            AP_AXIMM_0_RLAST,
    output  wire                            AP_AXIMM_0_RVALID,
    input  wire                            AP_AXIMM_0_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_0_AWADDR,
    output wire [7:0]                      M_AXIMM_0_AWLEN,
    output wire [2:0]                      M_AXIMM_0_AWSIZE,
    output wire [1:0]                      M_AXIMM_0_AWBURST,
    output wire [1:0]                      M_AXIMM_0_AWLOCK,
    output wire [3:0]                      M_AXIMM_0_AWCACHE,
    output wire [2:0]                      M_AXIMM_0_AWPROT,
    output wire [3:0]                      M_AXIMM_0_AWREGION,
    output wire [3:0]                      M_AXIMM_0_AWQOS,
    output wire                            M_AXIMM_0_AWVALID,
    input  wire                            M_AXIMM_0_AWREADY,
    output wire [M_AXIMM_0_DATA_WIDTH-1:0]   M_AXIMM_0_WDATA,
    output wire [M_AXIMM_0_DATA_WIDTH/8-1:0] M_AXIMM_0_WSTRB,
    output wire                            M_AXIMM_0_WLAST,
    output wire                            M_AXIMM_0_WVALID,
    input  wire                            M_AXIMM_0_WREADY,
    input  wire [1:0]                      M_AXIMM_0_BRESP,
    input  wire                            M_AXIMM_0_BVALID,
    output wire                            M_AXIMM_0_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_0_ARADDR,
    output wire [7:0]                      M_AXIMM_0_ARLEN,
    output wire [2:0]                      M_AXIMM_0_ARSIZE,
    output wire [1:0]                      M_AXIMM_0_ARBURST,
    output wire [1:0]                      M_AXIMM_0_ARLOCK,
    output wire [3:0]                      M_AXIMM_0_ARCACHE,
    output wire [2:0]                      M_AXIMM_0_ARPROT,
    output wire [3:0]                      M_AXIMM_0_ARREGION,
    output wire [3:0]                      M_AXIMM_0_ARQOS,
    output wire                            M_AXIMM_0_ARVALID,
    input  wire                            M_AXIMM_0_ARREADY,
    input  wire [M_AXIMM_0_DATA_WIDTH-1:0]   M_AXIMM_0_RDATA,
    input  wire [1:0]                      M_AXIMM_0_RRESP,
    input  wire                            M_AXIMM_0_RLAST,
    input  wire                            M_AXIMM_0_RVALID,
    output wire                            M_AXIMM_0_RREADY,
    //AXI-MM pass-through interface 1
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_1_AWADDR,
    input wire [7:0]                      AP_AXIMM_1_AWLEN,
    input wire [2:0]                      AP_AXIMM_1_AWSIZE,
    input wire [1:0]                      AP_AXIMM_1_AWBURST,
    input wire [1:0]                      AP_AXIMM_1_AWLOCK,
    input wire [3:0]                      AP_AXIMM_1_AWCACHE,
    input wire [2:0]                      AP_AXIMM_1_AWPROT,
    input wire [3:0]                      AP_AXIMM_1_AWREGION,
    input wire [3:0]                      AP_AXIMM_1_AWQOS,
    input wire                            AP_AXIMM_1_AWVALID,
    output  wire                            AP_AXIMM_1_AWREADY,
    input wire [M_AXIMM_1_DATA_WIDTH-1:0]   AP_AXIMM_1_WDATA,
    input wire [M_AXIMM_1_DATA_WIDTH/8-1:0] AP_AXIMM_1_WSTRB,
    input wire                            AP_AXIMM_1_WLAST,
    input wire                            AP_AXIMM_1_WVALID,
    output  wire                            AP_AXIMM_1_WREADY,
    output  wire [1:0]                      AP_AXIMM_1_BRESP,
    output  wire                            AP_AXIMM_1_BVALID,
    input wire                            AP_AXIMM_1_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_1_ARADDR,
    input wire [7:0]                      AP_AXIMM_1_ARLEN,
    input wire [2:0]                      AP_AXIMM_1_ARSIZE,
    input wire [1:0]                      AP_AXIMM_1_ARBURST,
    input wire [1:0]                      AP_AXIMM_1_ARLOCK,
    input wire [3:0]                      AP_AXIMM_1_ARCACHE,
    input wire [2:0]                      AP_AXIMM_1_ARPROT,
    input wire [3:0]                      AP_AXIMM_1_ARREGION,
    input wire [3:0]                      AP_AXIMM_1_ARQOS,
    input wire                            AP_AXIMM_1_ARVALID,
    output  wire                            AP_AXIMM_1_ARREADY,
    output  wire [M_AXIMM_1_DATA_WIDTH-1:0]   AP_AXIMM_1_RDATA,
    output  wire [1:0]                      AP_AXIMM_1_RRESP,
    output  wire                            AP_AXIMM_1_RLAST,
    output  wire                            AP_AXIMM_1_RVALID,
    input  wire                            AP_AXIMM_1_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_1_AWADDR,
    output wire [7:0]                      M_AXIMM_1_AWLEN,
    output wire [2:0]                      M_AXIMM_1_AWSIZE,
    output wire [1:0]                      M_AXIMM_1_AWBURST,
    output wire [1:0]                      M_AXIMM_1_AWLOCK,
    output wire [3:0]                      M_AXIMM_1_AWCACHE,
    output wire [2:0]                      M_AXIMM_1_AWPROT,
    output wire [3:0]                      M_AXIMM_1_AWREGION,
    output wire [3:0]                      M_AXIMM_1_AWQOS,
    output wire                            M_AXIMM_1_AWVALID,
    input  wire                            M_AXIMM_1_AWREADY,
    output wire [M_AXIMM_1_DATA_WIDTH-1:0]   M_AXIMM_1_WDATA,
    output wire [M_AXIMM_1_DATA_WIDTH/8-1:0] M_AXIMM_1_WSTRB,
    output wire                            M_AXIMM_1_WLAST,
    output wire                            M_AXIMM_1_WVALID,
    input  wire                            M_AXIMM_1_WREADY,
    input  wire [1:0]                      M_AXIMM_1_BRESP,
    input  wire                            M_AXIMM_1_BVALID,
    output wire                            M_AXIMM_1_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_1_ARADDR,
    output wire [7:0]                      M_AXIMM_1_ARLEN,
    output wire [2:0]                      M_AXIMM_1_ARSIZE,
    output wire [1:0]                      M_AXIMM_1_ARBURST,
    output wire [1:0]                      M_AXIMM_1_ARLOCK,
    output wire [3:0]                      M_AXIMM_1_ARCACHE,
    output wire [2:0]                      M_AXIMM_1_ARPROT,
    output wire [3:0]                      M_AXIMM_1_ARREGION,
    output wire [3:0]                      M_AXIMM_1_ARQOS,
    output wire                            M_AXIMM_1_ARVALID,
    input  wire                            M_AXIMM_1_ARREADY,
    input  wire [M_AXIMM_1_DATA_WIDTH-1:0]   M_AXIMM_1_RDATA,
    input  wire [1:0]                      M_AXIMM_1_RRESP,
    input  wire                            M_AXIMM_1_RLAST,
    input  wire                            M_AXIMM_1_RVALID,
    output wire                            M_AXIMM_1_RREADY,
    //AXI-MM pass-through interface 2
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_2_AWADDR,
    input wire [7:0]                      AP_AXIMM_2_AWLEN,
    input wire [2:0]                      AP_AXIMM_2_AWSIZE,
    input wire [1:0]                      AP_AXIMM_2_AWBURST,
    input wire [1:0]                      AP_AXIMM_2_AWLOCK,
    input wire [3:0]                      AP_AXIMM_2_AWCACHE,
    input wire [2:0]                      AP_AXIMM_2_AWPROT,
    input wire [3:0]                      AP_AXIMM_2_AWREGION,
    input wire [3:0]                      AP_AXIMM_2_AWQOS,
    input wire                            AP_AXIMM_2_AWVALID,
    output  wire                            AP_AXIMM_2_AWREADY,
    input wire [M_AXIMM_2_DATA_WIDTH-1:0]   AP_AXIMM_2_WDATA,
    input wire [M_AXIMM_2_DATA_WIDTH/8-1:0] AP_AXIMM_2_WSTRB,
    input wire                            AP_AXIMM_2_WLAST,
    input wire                            AP_AXIMM_2_WVALID,
    output  wire                            AP_AXIMM_2_WREADY,
    output  wire [1:0]                      AP_AXIMM_2_BRESP,
    output  wire                            AP_AXIMM_2_BVALID,
    input wire                            AP_AXIMM_2_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_2_ARADDR,
    input wire [7:0]                      AP_AXIMM_2_ARLEN,
    input wire [2:0]                      AP_AXIMM_2_ARSIZE,
    input wire [1:0]                      AP_AXIMM_2_ARBURST,
    input wire [1:0]                      AP_AXIMM_2_ARLOCK,
    input wire [3:0]                      AP_AXIMM_2_ARCACHE,
    input wire [2:0]                      AP_AXIMM_2_ARPROT,
    input wire [3:0]                      AP_AXIMM_2_ARREGION,
    input wire [3:0]                      AP_AXIMM_2_ARQOS,
    input wire                            AP_AXIMM_2_ARVALID,
    output  wire                            AP_AXIMM_2_ARREADY,
    output  wire [M_AXIMM_2_DATA_WIDTH-1:0]   AP_AXIMM_2_RDATA,
    output  wire [1:0]                      AP_AXIMM_2_RRESP,
    output  wire                            AP_AXIMM_2_RLAST,
    output  wire                            AP_AXIMM_2_RVALID,
    input  wire                            AP_AXIMM_2_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_2_AWADDR,
    output wire [7:0]                      M_AXIMM_2_AWLEN,
    output wire [2:0]                      M_AXIMM_2_AWSIZE,
    output wire [1:0]                      M_AXIMM_2_AWBURST,
    output wire [1:0]                      M_AXIMM_2_AWLOCK,
    output wire [3:0]                      M_AXIMM_2_AWCACHE,
    output wire [2:0]                      M_AXIMM_2_AWPROT,
    output wire [3:0]                      M_AXIMM_2_AWREGION,
    output wire [3:0]                      M_AXIMM_2_AWQOS,
    output wire                            M_AXIMM_2_AWVALID,
    input  wire                            M_AXIMM_2_AWREADY,
    output wire [M_AXIMM_2_DATA_WIDTH-1:0]   M_AXIMM_2_WDATA,
    output wire [M_AXIMM_2_DATA_WIDTH/8-1:0] M_AXIMM_2_WSTRB,
    output wire                            M_AXIMM_2_WLAST,
    output wire                            M_AXIMM_2_WVALID,
    input  wire                            M_AXIMM_2_WREADY,
    input  wire [1:0]                      M_AXIMM_2_BRESP,
    input  wire                            M_AXIMM_2_BVALID,
    output wire                            M_AXIMM_2_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_2_ARADDR,
    output wire [7:0]                      M_AXIMM_2_ARLEN,
    output wire [2:0]                      M_AXIMM_2_ARSIZE,
    output wire [1:0]                      M_AXIMM_2_ARBURST,
    output wire [1:0]                      M_AXIMM_2_ARLOCK,
    output wire [3:0]                      M_AXIMM_2_ARCACHE,
    output wire [2:0]                      M_AXIMM_2_ARPROT,
    output wire [3:0]                      M_AXIMM_2_ARREGION,
    output wire [3:0]                      M_AXIMM_2_ARQOS,
    output wire                            M_AXIMM_2_ARVALID,
    input  wire                            M_AXIMM_2_ARREADY,
    input  wire [M_AXIMM_2_DATA_WIDTH-1:0]   M_AXIMM_2_RDATA,
    input  wire [1:0]                      M_AXIMM_2_RRESP,
    input  wire                            M_AXIMM_2_RLAST,
    input  wire                            M_AXIMM_2_RVALID,
    output wire                            M_AXIMM_2_RREADY,
    //AXI-MM pass-through interface 3
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_3_AWADDR,
    input wire [7:0]                      AP_AXIMM_3_AWLEN,
    input wire [2:0]                      AP_AXIMM_3_AWSIZE,
    input wire [1:0]                      AP_AXIMM_3_AWBURST,
    input wire [1:0]                      AP_AXIMM_3_AWLOCK,
    input wire [3:0]                      AP_AXIMM_3_AWCACHE,
    input wire [2:0]                      AP_AXIMM_3_AWPROT,
    input wire [3:0]                      AP_AXIMM_3_AWREGION,
    input wire [3:0]                      AP_AXIMM_3_AWQOS,
    input wire                            AP_AXIMM_3_AWVALID,
    output  wire                            AP_AXIMM_3_AWREADY,
    input wire [M_AXIMM_3_DATA_WIDTH-1:0]   AP_AXIMM_3_WDATA,
    input wire [M_AXIMM_3_DATA_WIDTH/8-1:0] AP_AXIMM_3_WSTRB,
    input wire                            AP_AXIMM_3_WLAST,
    input wire                            AP_AXIMM_3_WVALID,
    output  wire                            AP_AXIMM_3_WREADY,
    output  wire [1:0]                      AP_AXIMM_3_BRESP,
    output  wire                            AP_AXIMM_3_BVALID,
    input wire                            AP_AXIMM_3_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_3_ARADDR,
    input wire [7:0]                      AP_AXIMM_3_ARLEN,
    input wire [2:0]                      AP_AXIMM_3_ARSIZE,
    input wire [1:0]                      AP_AXIMM_3_ARBURST,
    input wire [1:0]                      AP_AXIMM_3_ARLOCK,
    input wire [3:0]                      AP_AXIMM_3_ARCACHE,
    input wire [2:0]                      AP_AXIMM_3_ARPROT,
    input wire [3:0]                      AP_AXIMM_3_ARREGION,
    input wire [3:0]                      AP_AXIMM_3_ARQOS,
    input wire                            AP_AXIMM_3_ARVALID,
    output  wire                            AP_AXIMM_3_ARREADY,
    output  wire [M_AXIMM_3_DATA_WIDTH-1:0]   AP_AXIMM_3_RDATA,
    output  wire [1:0]                      AP_AXIMM_3_RRESP,
    output  wire                            AP_AXIMM_3_RLAST,
    output  wire                            AP_AXIMM_3_RVALID,
    input  wire                            AP_AXIMM_3_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_3_AWADDR,
    output wire [7:0]                      M_AXIMM_3_AWLEN,
    output wire [2:0]                      M_AXIMM_3_AWSIZE,
    output wire [1:0]                      M_AXIMM_3_AWBURST,
    output wire [1:0]                      M_AXIMM_3_AWLOCK,
    output wire [3:0]                      M_AXIMM_3_AWCACHE,
    output wire [2:0]                      M_AXIMM_3_AWPROT,
    output wire [3:0]                      M_AXIMM_3_AWREGION,
    output wire [3:0]                      M_AXIMM_3_AWQOS,
    output wire                            M_AXIMM_3_AWVALID,
    input  wire                            M_AXIMM_3_AWREADY,
    output wire [M_AXIMM_3_DATA_WIDTH-1:0]   M_AXIMM_3_WDATA,
    output wire [M_AXIMM_3_DATA_WIDTH/8-1:0] M_AXIMM_3_WSTRB,
    output wire                            M_AXIMM_3_WLAST,
    output wire                            M_AXIMM_3_WVALID,
    input  wire                            M_AXIMM_3_WREADY,
    input  wire [1:0]                      M_AXIMM_3_BRESP,
    input  wire                            M_AXIMM_3_BVALID,
    output wire                            M_AXIMM_3_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_3_ARADDR,
    output wire [7:0]                      M_AXIMM_3_ARLEN,
    output wire [2:0]                      M_AXIMM_3_ARSIZE,
    output wire [1:0]                      M_AXIMM_3_ARBURST,
    output wire [1:0]                      M_AXIMM_3_ARLOCK,
    output wire [3:0]                      M_AXIMM_3_ARCACHE,
    output wire [2:0]                      M_AXIMM_3_ARPROT,
    output wire [3:0]                      M_AXIMM_3_ARREGION,
    output wire [3:0]                      M_AXIMM_3_ARQOS,
    output wire                            M_AXIMM_3_ARVALID,
    input  wire                            M_AXIMM_3_ARREADY,
    input  wire [M_AXIMM_3_DATA_WIDTH-1:0]   M_AXIMM_3_RDATA,
    input  wire [1:0]                      M_AXIMM_3_RRESP,
    input  wire                            M_AXIMM_3_RLAST,
    input  wire                            M_AXIMM_3_RVALID,
    output wire                            M_AXIMM_3_RREADY,
    //AXI-MM pass-through interface 4
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_4_AWADDR,
    input wire [7:0]                      AP_AXIMM_4_AWLEN,
    input wire [2:0]                      AP_AXIMM_4_AWSIZE,
    input wire [1:0]                      AP_AXIMM_4_AWBURST,
    input wire [1:0]                      AP_AXIMM_4_AWLOCK,
    input wire [3:0]                      AP_AXIMM_4_AWCACHE,
    input wire [2:0]                      AP_AXIMM_4_AWPROT,
    input wire [3:0]                      AP_AXIMM_4_AWREGION,
    input wire [3:0]                      AP_AXIMM_4_AWQOS,
    input wire                            AP_AXIMM_4_AWVALID,
    output  wire                            AP_AXIMM_4_AWREADY,
    input wire [M_AXIMM_4_DATA_WIDTH-1:0]   AP_AXIMM_4_WDATA,
    input wire [M_AXIMM_4_DATA_WIDTH/8-1:0] AP_AXIMM_4_WSTRB,
    input wire                            AP_AXIMM_4_WLAST,
    input wire                            AP_AXIMM_4_WVALID,
    output  wire                            AP_AXIMM_4_WREADY,
    output  wire [1:0]                      AP_AXIMM_4_BRESP,
    output  wire                            AP_AXIMM_4_BVALID,
    input wire                            AP_AXIMM_4_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_4_ARADDR,
    input wire [7:0]                      AP_AXIMM_4_ARLEN,
    input wire [2:0]                      AP_AXIMM_4_ARSIZE,
    input wire [1:0]                      AP_AXIMM_4_ARBURST,
    input wire [1:0]                      AP_AXIMM_4_ARLOCK,
    input wire [3:0]                      AP_AXIMM_4_ARCACHE,
    input wire [2:0]                      AP_AXIMM_4_ARPROT,
    input wire [3:0]                      AP_AXIMM_4_ARREGION,
    input wire [3:0]                      AP_AXIMM_4_ARQOS,
    input wire                            AP_AXIMM_4_ARVALID,
    output  wire                            AP_AXIMM_4_ARREADY,
    output  wire [M_AXIMM_4_DATA_WIDTH-1:0]   AP_AXIMM_4_RDATA,
    output  wire [1:0]                      AP_AXIMM_4_RRESP,
    output  wire                            AP_AXIMM_4_RLAST,
    output  wire                            AP_AXIMM_4_RVALID,
    input  wire                            AP_AXIMM_4_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_4_AWADDR,
    output wire [7:0]                      M_AXIMM_4_AWLEN,
    output wire [2:0]                      M_AXIMM_4_AWSIZE,
    output wire [1:0]                      M_AXIMM_4_AWBURST,
    output wire [1:0]                      M_AXIMM_4_AWLOCK,
    output wire [3:0]                      M_AXIMM_4_AWCACHE,
    output wire [2:0]                      M_AXIMM_4_AWPROT,
    output wire [3:0]                      M_AXIMM_4_AWREGION,
    output wire [3:0]                      M_AXIMM_4_AWQOS,
    output wire                            M_AXIMM_4_AWVALID,
    input  wire                            M_AXIMM_4_AWREADY,
    output wire [M_AXIMM_4_DATA_WIDTH-1:0]   M_AXIMM_4_WDATA,
    output wire [M_AXIMM_4_DATA_WIDTH/8-1:0] M_AXIMM_4_WSTRB,
    output wire                            M_AXIMM_4_WLAST,
    output wire                            M_AXIMM_4_WVALID,
    input  wire                            M_AXIMM_4_WREADY,
    input  wire [1:0]                      M_AXIMM_4_BRESP,
    input  wire                            M_AXIMM_4_BVALID,
    output wire                            M_AXIMM_4_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_4_ARADDR,
    output wire [7:0]                      M_AXIMM_4_ARLEN,
    output wire [2:0]                      M_AXIMM_4_ARSIZE,
    output wire [1:0]                      M_AXIMM_4_ARBURST,
    output wire [1:0]                      M_AXIMM_4_ARLOCK,
    output wire [3:0]                      M_AXIMM_4_ARCACHE,
    output wire [2:0]                      M_AXIMM_4_ARPROT,
    output wire [3:0]                      M_AXIMM_4_ARREGION,
    output wire [3:0]                      M_AXIMM_4_ARQOS,
    output wire                            M_AXIMM_4_ARVALID,
    input  wire                            M_AXIMM_4_ARREADY,
    input  wire [M_AXIMM_4_DATA_WIDTH-1:0]   M_AXIMM_4_RDATA,
    input  wire [1:0]                      M_AXIMM_4_RRESP,
    input  wire                            M_AXIMM_4_RLAST,
    input  wire                            M_AXIMM_4_RVALID,
    output wire                            M_AXIMM_4_RREADY,
    //AXI-MM pass-through interface 5
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_5_AWADDR,
    input wire [7:0]                      AP_AXIMM_5_AWLEN,
    input wire [2:0]                      AP_AXIMM_5_AWSIZE,
    input wire [1:0]                      AP_AXIMM_5_AWBURST,
    input wire [1:0]                      AP_AXIMM_5_AWLOCK,
    input wire [3:0]                      AP_AXIMM_5_AWCACHE,
    input wire [2:0]                      AP_AXIMM_5_AWPROT,
    input wire [3:0]                      AP_AXIMM_5_AWREGION,
    input wire [3:0]                      AP_AXIMM_5_AWQOS,
    input wire                            AP_AXIMM_5_AWVALID,
    output  wire                            AP_AXIMM_5_AWREADY,
    input wire [M_AXIMM_5_DATA_WIDTH-1:0]   AP_AXIMM_5_WDATA,
    input wire [M_AXIMM_5_DATA_WIDTH/8-1:0] AP_AXIMM_5_WSTRB,
    input wire                            AP_AXIMM_5_WLAST,
    input wire                            AP_AXIMM_5_WVALID,
    output  wire                            AP_AXIMM_5_WREADY,
    output  wire [1:0]                      AP_AXIMM_5_BRESP,
    output  wire                            AP_AXIMM_5_BVALID,
    input wire                            AP_AXIMM_5_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_5_ARADDR,
    input wire [7:0]                      AP_AXIMM_5_ARLEN,
    input wire [2:0]                      AP_AXIMM_5_ARSIZE,
    input wire [1:0]                      AP_AXIMM_5_ARBURST,
    input wire [1:0]                      AP_AXIMM_5_ARLOCK,
    input wire [3:0]                      AP_AXIMM_5_ARCACHE,
    input wire [2:0]                      AP_AXIMM_5_ARPROT,
    input wire [3:0]                      AP_AXIMM_5_ARREGION,
    input wire [3:0]                      AP_AXIMM_5_ARQOS,
    input wire                            AP_AXIMM_5_ARVALID,
    output  wire                            AP_AXIMM_5_ARREADY,
    output  wire [M_AXIMM_5_DATA_WIDTH-1:0]   AP_AXIMM_5_RDATA,
    output  wire [1:0]                      AP_AXIMM_5_RRESP,
    output  wire                            AP_AXIMM_5_RLAST,
    output  wire                            AP_AXIMM_5_RVALID,
    input  wire                            AP_AXIMM_5_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_5_AWADDR,
    output wire [7:0]                      M_AXIMM_5_AWLEN,
    output wire [2:0]                      M_AXIMM_5_AWSIZE,
    output wire [1:0]                      M_AXIMM_5_AWBURST,
    output wire [1:0]                      M_AXIMM_5_AWLOCK,
    output wire [3:0]                      M_AXIMM_5_AWCACHE,
    output wire [2:0]                      M_AXIMM_5_AWPROT,
    output wire [3:0]                      M_AXIMM_5_AWREGION,
    output wire [3:0]                      M_AXIMM_5_AWQOS,
    output wire                            M_AXIMM_5_AWVALID,
    input  wire                            M_AXIMM_5_AWREADY,
    output wire [M_AXIMM_5_DATA_WIDTH-1:0]   M_AXIMM_5_WDATA,
    output wire [M_AXIMM_5_DATA_WIDTH/8-1:0] M_AXIMM_5_WSTRB,
    output wire                            M_AXIMM_5_WLAST,
    output wire                            M_AXIMM_5_WVALID,
    input  wire                            M_AXIMM_5_WREADY,
    input  wire [1:0]                      M_AXIMM_5_BRESP,
    input  wire                            M_AXIMM_5_BVALID,
    output wire                            M_AXIMM_5_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_5_ARADDR,
    output wire [7:0]                      M_AXIMM_5_ARLEN,
    output wire [2:0]                      M_AXIMM_5_ARSIZE,
    output wire [1:0]                      M_AXIMM_5_ARBURST,
    output wire [1:0]                      M_AXIMM_5_ARLOCK,
    output wire [3:0]                      M_AXIMM_5_ARCACHE,
    output wire [2:0]                      M_AXIMM_5_ARPROT,
    output wire [3:0]                      M_AXIMM_5_ARREGION,
    output wire [3:0]                      M_AXIMM_5_ARQOS,
    output wire                            M_AXIMM_5_ARVALID,
    input  wire                            M_AXIMM_5_ARREADY,
    input  wire [M_AXIMM_5_DATA_WIDTH-1:0]   M_AXIMM_5_RDATA,
    input  wire [1:0]                      M_AXIMM_5_RRESP,
    input  wire                            M_AXIMM_5_RLAST,
    input  wire                            M_AXIMM_5_RVALID,
    output wire                            M_AXIMM_5_RREADY,
    //AXI-MM pass-through interface 6
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_6_AWADDR,
    input wire [7:0]                      AP_AXIMM_6_AWLEN,
    input wire [2:0]                      AP_AXIMM_6_AWSIZE,
    input wire [1:0]                      AP_AXIMM_6_AWBURST,
    input wire [1:0]                      AP_AXIMM_6_AWLOCK,
    input wire [3:0]                      AP_AXIMM_6_AWCACHE,
    input wire [2:0]                      AP_AXIMM_6_AWPROT,
    input wire [3:0]                      AP_AXIMM_6_AWREGION,
    input wire [3:0]                      AP_AXIMM_6_AWQOS,
    input wire                            AP_AXIMM_6_AWVALID,
    output  wire                            AP_AXIMM_6_AWREADY,
    input wire [M_AXIMM_6_DATA_WIDTH-1:0]   AP_AXIMM_6_WDATA,
    input wire [M_AXIMM_6_DATA_WIDTH/8-1:0] AP_AXIMM_6_WSTRB,
    input wire                            AP_AXIMM_6_WLAST,
    input wire                            AP_AXIMM_6_WVALID,
    output  wire                            AP_AXIMM_6_WREADY,
    output  wire [1:0]                      AP_AXIMM_6_BRESP,
    output  wire                            AP_AXIMM_6_BVALID,
    input wire                            AP_AXIMM_6_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_6_ARADDR,
    input wire [7:0]                      AP_AXIMM_6_ARLEN,
    input wire [2:0]                      AP_AXIMM_6_ARSIZE,
    input wire [1:0]                      AP_AXIMM_6_ARBURST,
    input wire [1:0]                      AP_AXIMM_6_ARLOCK,
    input wire [3:0]                      AP_AXIMM_6_ARCACHE,
    input wire [2:0]                      AP_AXIMM_6_ARPROT,
    input wire [3:0]                      AP_AXIMM_6_ARREGION,
    input wire [3:0]                      AP_AXIMM_6_ARQOS,
    input wire                            AP_AXIMM_6_ARVALID,
    output  wire                            AP_AXIMM_6_ARREADY,
    output  wire [M_AXIMM_6_DATA_WIDTH-1:0]   AP_AXIMM_6_RDATA,
    output  wire [1:0]                      AP_AXIMM_6_RRESP,
    output  wire                            AP_AXIMM_6_RLAST,
    output  wire                            AP_AXIMM_6_RVALID,
    input  wire                            AP_AXIMM_6_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_6_AWADDR,
    output wire [7:0]                      M_AXIMM_6_AWLEN,
    output wire [2:0]                      M_AXIMM_6_AWSIZE,
    output wire [1:0]                      M_AXIMM_6_AWBURST,
    output wire [1:0]                      M_AXIMM_6_AWLOCK,
    output wire [3:0]                      M_AXIMM_6_AWCACHE,
    output wire [2:0]                      M_AXIMM_6_AWPROT,
    output wire [3:0]                      M_AXIMM_6_AWREGION,
    output wire [3:0]                      M_AXIMM_6_AWQOS,
    output wire                            M_AXIMM_6_AWVALID,
    input  wire                            M_AXIMM_6_AWREADY,
    output wire [M_AXIMM_6_DATA_WIDTH-1:0]   M_AXIMM_6_WDATA,
    output wire [M_AXIMM_6_DATA_WIDTH/8-1:0] M_AXIMM_6_WSTRB,
    output wire                            M_AXIMM_6_WLAST,
    output wire                            M_AXIMM_6_WVALID,
    input  wire                            M_AXIMM_6_WREADY,
    input  wire [1:0]                      M_AXIMM_6_BRESP,
    input  wire                            M_AXIMM_6_BVALID,
    output wire                            M_AXIMM_6_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_6_ARADDR,
    output wire [7:0]                      M_AXIMM_6_ARLEN,
    output wire [2:0]                      M_AXIMM_6_ARSIZE,
    output wire [1:0]                      M_AXIMM_6_ARBURST,
    output wire [1:0]                      M_AXIMM_6_ARLOCK,
    output wire [3:0]                      M_AXIMM_6_ARCACHE,
    output wire [2:0]                      M_AXIMM_6_ARPROT,
    output wire [3:0]                      M_AXIMM_6_ARREGION,
    output wire [3:0]                      M_AXIMM_6_ARQOS,
    output wire                            M_AXIMM_6_ARVALID,
    input  wire                            M_AXIMM_6_ARREADY,
    input  wire [M_AXIMM_6_DATA_WIDTH-1:0]   M_AXIMM_6_RDATA,
    input  wire [1:0]                      M_AXIMM_6_RRESP,
    input  wire                            M_AXIMM_6_RLAST,
    input  wire                            M_AXIMM_6_RVALID,
    output wire                            M_AXIMM_6_RREADY,
    //AXI-MM pass-through interface 7
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_7_AWADDR,
    input wire [7:0]                      AP_AXIMM_7_AWLEN,
    input wire [2:0]                      AP_AXIMM_7_AWSIZE,
    input wire [1:0]                      AP_AXIMM_7_AWBURST,
    input wire [1:0]                      AP_AXIMM_7_AWLOCK,
    input wire [3:0]                      AP_AXIMM_7_AWCACHE,
    input wire [2:0]                      AP_AXIMM_7_AWPROT,
    input wire [3:0]                      AP_AXIMM_7_AWREGION,
    input wire [3:0]                      AP_AXIMM_7_AWQOS,
    input wire                            AP_AXIMM_7_AWVALID,
    output  wire                            AP_AXIMM_7_AWREADY,
    input wire [M_AXIMM_7_DATA_WIDTH-1:0]   AP_AXIMM_7_WDATA,
    input wire [M_AXIMM_7_DATA_WIDTH/8-1:0] AP_AXIMM_7_WSTRB,
    input wire                            AP_AXIMM_7_WLAST,
    input wire                            AP_AXIMM_7_WVALID,
    output  wire                            AP_AXIMM_7_WREADY,
    output  wire [1:0]                      AP_AXIMM_7_BRESP,
    output  wire                            AP_AXIMM_7_BVALID,
    input wire                            AP_AXIMM_7_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_7_ARADDR,
    input wire [7:0]                      AP_AXIMM_7_ARLEN,
    input wire [2:0]                      AP_AXIMM_7_ARSIZE,
    input wire [1:0]                      AP_AXIMM_7_ARBURST,
    input wire [1:0]                      AP_AXIMM_7_ARLOCK,
    input wire [3:0]                      AP_AXIMM_7_ARCACHE,
    input wire [2:0]                      AP_AXIMM_7_ARPROT,
    input wire [3:0]                      AP_AXIMM_7_ARREGION,
    input wire [3:0]                      AP_AXIMM_7_ARQOS,
    input wire                            AP_AXIMM_7_ARVALID,
    output  wire                            AP_AXIMM_7_ARREADY,
    output  wire [M_AXIMM_7_DATA_WIDTH-1:0]   AP_AXIMM_7_RDATA,
    output  wire [1:0]                      AP_AXIMM_7_RRESP,
    output  wire                            AP_AXIMM_7_RLAST,
    output  wire                            AP_AXIMM_7_RVALID,
    input  wire                            AP_AXIMM_7_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_7_AWADDR,
    output wire [7:0]                      M_AXIMM_7_AWLEN,
    output wire [2:0]                      M_AXIMM_7_AWSIZE,
    output wire [1:0]                      M_AXIMM_7_AWBURST,
    output wire [1:0]                      M_AXIMM_7_AWLOCK,
    output wire [3:0]                      M_AXIMM_7_AWCACHE,
    output wire [2:0]                      M_AXIMM_7_AWPROT,
    output wire [3:0]                      M_AXIMM_7_AWREGION,
    output wire [3:0]                      M_AXIMM_7_AWQOS,
    output wire                            M_AXIMM_7_AWVALID,
    input  wire                            M_AXIMM_7_AWREADY,
    output wire [M_AXIMM_7_DATA_WIDTH-1:0]   M_AXIMM_7_WDATA,
    output wire [M_AXIMM_7_DATA_WIDTH/8-1:0] M_AXIMM_7_WSTRB,
    output wire                            M_AXIMM_7_WLAST,
    output wire                            M_AXIMM_7_WVALID,
    input  wire                            M_AXIMM_7_WREADY,
    input  wire [1:0]                      M_AXIMM_7_BRESP,
    input  wire                            M_AXIMM_7_BVALID,
    output wire                            M_AXIMM_7_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_7_ARADDR,
    output wire [7:0]                      M_AXIMM_7_ARLEN,
    output wire [2:0]                      M_AXIMM_7_ARSIZE,
    output wire [1:0]                      M_AXIMM_7_ARBURST,
    output wire [1:0]                      M_AXIMM_7_ARLOCK,
    output wire [3:0]                      M_AXIMM_7_ARCACHE,
    output wire [2:0]                      M_AXIMM_7_ARPROT,
    output wire [3:0]                      M_AXIMM_7_ARREGION,
    output wire [3:0]                      M_AXIMM_7_ARQOS,
    output wire                            M_AXIMM_7_ARVALID,
    input  wire                            M_AXIMM_7_ARREADY,
    input  wire [M_AXIMM_7_DATA_WIDTH-1:0]   M_AXIMM_7_RDATA,
    input  wire [1:0]                      M_AXIMM_7_RRESP,
    input  wire                            M_AXIMM_7_RLAST,
    input  wire                            M_AXIMM_7_RVALID,
    output wire                            M_AXIMM_7_RREADY,
    //AXI-MM pass-through interface 8
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_8_AWADDR,
    input wire [7:0]                      AP_AXIMM_8_AWLEN,
    input wire [2:0]                      AP_AXIMM_8_AWSIZE,
    input wire [1:0]                      AP_AXIMM_8_AWBURST,
    input wire [1:0]                      AP_AXIMM_8_AWLOCK,
    input wire [3:0]                      AP_AXIMM_8_AWCACHE,
    input wire [2:0]                      AP_AXIMM_8_AWPROT,
    input wire [3:0]                      AP_AXIMM_8_AWREGION,
    input wire [3:0]                      AP_AXIMM_8_AWQOS,
    input wire                            AP_AXIMM_8_AWVALID,
    output  wire                            AP_AXIMM_8_AWREADY,
    input wire [M_AXIMM_8_DATA_WIDTH-1:0]   AP_AXIMM_8_WDATA,
    input wire [M_AXIMM_8_DATA_WIDTH/8-1:0] AP_AXIMM_8_WSTRB,
    input wire                            AP_AXIMM_8_WLAST,
    input wire                            AP_AXIMM_8_WVALID,
    output  wire                            AP_AXIMM_8_WREADY,
    output  wire [1:0]                      AP_AXIMM_8_BRESP,
    output  wire                            AP_AXIMM_8_BVALID,
    input wire                            AP_AXIMM_8_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_8_ARADDR,
    input wire [7:0]                      AP_AXIMM_8_ARLEN,
    input wire [2:0]                      AP_AXIMM_8_ARSIZE,
    input wire [1:0]                      AP_AXIMM_8_ARBURST,
    input wire [1:0]                      AP_AXIMM_8_ARLOCK,
    input wire [3:0]                      AP_AXIMM_8_ARCACHE,
    input wire [2:0]                      AP_AXIMM_8_ARPROT,
    input wire [3:0]                      AP_AXIMM_8_ARREGION,
    input wire [3:0]                      AP_AXIMM_8_ARQOS,
    input wire                            AP_AXIMM_8_ARVALID,
    output  wire                            AP_AXIMM_8_ARREADY,
    output  wire [M_AXIMM_8_DATA_WIDTH-1:0]   AP_AXIMM_8_RDATA,
    output  wire [1:0]                      AP_AXIMM_8_RRESP,
    output  wire                            AP_AXIMM_8_RLAST,
    output  wire                            AP_AXIMM_8_RVALID,
    input  wire                            AP_AXIMM_8_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_8_AWADDR,
    output wire [7:0]                      M_AXIMM_8_AWLEN,
    output wire [2:0]                      M_AXIMM_8_AWSIZE,
    output wire [1:0]                      M_AXIMM_8_AWBURST,
    output wire [1:0]                      M_AXIMM_8_AWLOCK,
    output wire [3:0]                      M_AXIMM_8_AWCACHE,
    output wire [2:0]                      M_AXIMM_8_AWPROT,
    output wire [3:0]                      M_AXIMM_8_AWREGION,
    output wire [3:0]                      M_AXIMM_8_AWQOS,
    output wire                            M_AXIMM_8_AWVALID,
    input  wire                            M_AXIMM_8_AWREADY,
    output wire [M_AXIMM_8_DATA_WIDTH-1:0]   M_AXIMM_8_WDATA,
    output wire [M_AXIMM_8_DATA_WIDTH/8-1:0] M_AXIMM_8_WSTRB,
    output wire                            M_AXIMM_8_WLAST,
    output wire                            M_AXIMM_8_WVALID,
    input  wire                            M_AXIMM_8_WREADY,
    input  wire [1:0]                      M_AXIMM_8_BRESP,
    input  wire                            M_AXIMM_8_BVALID,
    output wire                            M_AXIMM_8_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_8_ARADDR,
    output wire [7:0]                      M_AXIMM_8_ARLEN,
    output wire [2:0]                      M_AXIMM_8_ARSIZE,
    output wire [1:0]                      M_AXIMM_8_ARBURST,
    output wire [1:0]                      M_AXIMM_8_ARLOCK,
    output wire [3:0]                      M_AXIMM_8_ARCACHE,
    output wire [2:0]                      M_AXIMM_8_ARPROT,
    output wire [3:0]                      M_AXIMM_8_ARREGION,
    output wire [3:0]                      M_AXIMM_8_ARQOS,
    output wire                            M_AXIMM_8_ARVALID,
    input  wire                            M_AXIMM_8_ARREADY,
    input  wire [M_AXIMM_8_DATA_WIDTH-1:0]   M_AXIMM_8_RDATA,
    input  wire [1:0]                      M_AXIMM_8_RRESP,
    input  wire                            M_AXIMM_8_RLAST,
    input  wire                            M_AXIMM_8_RVALID,
    output wire                            M_AXIMM_8_RREADY,
    //AXI-MM pass-through interface 9
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_9_AWADDR,
    input wire [7:0]                      AP_AXIMM_9_AWLEN,
    input wire [2:0]                      AP_AXIMM_9_AWSIZE,
    input wire [1:0]                      AP_AXIMM_9_AWBURST,
    input wire [1:0]                      AP_AXIMM_9_AWLOCK,
    input wire [3:0]                      AP_AXIMM_9_AWCACHE,
    input wire [2:0]                      AP_AXIMM_9_AWPROT,
    input wire [3:0]                      AP_AXIMM_9_AWREGION,
    input wire [3:0]                      AP_AXIMM_9_AWQOS,
    input wire                            AP_AXIMM_9_AWVALID,
    output  wire                            AP_AXIMM_9_AWREADY,
    input wire [M_AXIMM_9_DATA_WIDTH-1:0]   AP_AXIMM_9_WDATA,
    input wire [M_AXIMM_9_DATA_WIDTH/8-1:0] AP_AXIMM_9_WSTRB,
    input wire                            AP_AXIMM_9_WLAST,
    input wire                            AP_AXIMM_9_WVALID,
    output  wire                            AP_AXIMM_9_WREADY,
    output  wire [1:0]                      AP_AXIMM_9_BRESP,
    output  wire                            AP_AXIMM_9_BVALID,
    input wire                            AP_AXIMM_9_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_9_ARADDR,
    input wire [7:0]                      AP_AXIMM_9_ARLEN,
    input wire [2:0]                      AP_AXIMM_9_ARSIZE,
    input wire [1:0]                      AP_AXIMM_9_ARBURST,
    input wire [1:0]                      AP_AXIMM_9_ARLOCK,
    input wire [3:0]                      AP_AXIMM_9_ARCACHE,
    input wire [2:0]                      AP_AXIMM_9_ARPROT,
    input wire [3:0]                      AP_AXIMM_9_ARREGION,
    input wire [3:0]                      AP_AXIMM_9_ARQOS,
    input wire                            AP_AXIMM_9_ARVALID,
    output  wire                            AP_AXIMM_9_ARREADY,
    output  wire [M_AXIMM_9_DATA_WIDTH-1:0]   AP_AXIMM_9_RDATA,
    output  wire [1:0]                      AP_AXIMM_9_RRESP,
    output  wire                            AP_AXIMM_9_RLAST,
    output  wire                            AP_AXIMM_9_RVALID,
    input  wire                            AP_AXIMM_9_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_9_AWADDR,
    output wire [7:0]                      M_AXIMM_9_AWLEN,
    output wire [2:0]                      M_AXIMM_9_AWSIZE,
    output wire [1:0]                      M_AXIMM_9_AWBURST,
    output wire [1:0]                      M_AXIMM_9_AWLOCK,
    output wire [3:0]                      M_AXIMM_9_AWCACHE,
    output wire [2:0]                      M_AXIMM_9_AWPROT,
    output wire [3:0]                      M_AXIMM_9_AWREGION,
    output wire [3:0]                      M_AXIMM_9_AWQOS,
    output wire                            M_AXIMM_9_AWVALID,
    input  wire                            M_AXIMM_9_AWREADY,
    output wire [M_AXIMM_9_DATA_WIDTH-1:0]   M_AXIMM_9_WDATA,
    output wire [M_AXIMM_9_DATA_WIDTH/8-1:0] M_AXIMM_9_WSTRB,
    output wire                            M_AXIMM_9_WLAST,
    output wire                            M_AXIMM_9_WVALID,
    input  wire                            M_AXIMM_9_WREADY,
    input  wire [1:0]                      M_AXIMM_9_BRESP,
    input  wire                            M_AXIMM_9_BVALID,
    output wire                            M_AXIMM_9_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_9_ARADDR,
    output wire [7:0]                      M_AXIMM_9_ARLEN,
    output wire [2:0]                      M_AXIMM_9_ARSIZE,
    output wire [1:0]                      M_AXIMM_9_ARBURST,
    output wire [1:0]                      M_AXIMM_9_ARLOCK,
    output wire [3:0]                      M_AXIMM_9_ARCACHE,
    output wire [2:0]                      M_AXIMM_9_ARPROT,
    output wire [3:0]                      M_AXIMM_9_ARREGION,
    output wire [3:0]                      M_AXIMM_9_ARQOS,
    output wire                            M_AXIMM_9_ARVALID,
    input  wire                            M_AXIMM_9_ARREADY,
    input  wire [M_AXIMM_9_DATA_WIDTH-1:0]   M_AXIMM_9_RDATA,
    input  wire [1:0]                      M_AXIMM_9_RRESP,
    input  wire                            M_AXIMM_9_RLAST,
    input  wire                            M_AXIMM_9_RVALID,
    output wire                            M_AXIMM_9_RREADY,
    //AXI-MM pass-through interface 10
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_10_AWADDR,
    input wire [7:0]                      AP_AXIMM_10_AWLEN,
    input wire [2:0]                      AP_AXIMM_10_AWSIZE,
    input wire [1:0]                      AP_AXIMM_10_AWBURST,
    input wire [1:0]                      AP_AXIMM_10_AWLOCK,
    input wire [3:0]                      AP_AXIMM_10_AWCACHE,
    input wire [2:0]                      AP_AXIMM_10_AWPROT,
    input wire [3:0]                      AP_AXIMM_10_AWREGION,
    input wire [3:0]                      AP_AXIMM_10_AWQOS,
    input wire                            AP_AXIMM_10_AWVALID,
    output  wire                            AP_AXIMM_10_AWREADY,
    input wire [M_AXIMM_10_DATA_WIDTH-1:0]   AP_AXIMM_10_WDATA,
    input wire [M_AXIMM_10_DATA_WIDTH/8-1:0] AP_AXIMM_10_WSTRB,
    input wire                            AP_AXIMM_10_WLAST,
    input wire                            AP_AXIMM_10_WVALID,
    output  wire                            AP_AXIMM_10_WREADY,
    output  wire [1:0]                      AP_AXIMM_10_BRESP,
    output  wire                            AP_AXIMM_10_BVALID,
    input wire                            AP_AXIMM_10_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_10_ARADDR,
    input wire [7:0]                      AP_AXIMM_10_ARLEN,
    input wire [2:0]                      AP_AXIMM_10_ARSIZE,
    input wire [1:0]                      AP_AXIMM_10_ARBURST,
    input wire [1:0]                      AP_AXIMM_10_ARLOCK,
    input wire [3:0]                      AP_AXIMM_10_ARCACHE,
    input wire [2:0]                      AP_AXIMM_10_ARPROT,
    input wire [3:0]                      AP_AXIMM_10_ARREGION,
    input wire [3:0]                      AP_AXIMM_10_ARQOS,
    input wire                            AP_AXIMM_10_ARVALID,
    output  wire                            AP_AXIMM_10_ARREADY,
    output  wire [M_AXIMM_10_DATA_WIDTH-1:0]   AP_AXIMM_10_RDATA,
    output  wire [1:0]                      AP_AXIMM_10_RRESP,
    output  wire                            AP_AXIMM_10_RLAST,
    output  wire                            AP_AXIMM_10_RVALID,
    input  wire                            AP_AXIMM_10_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_10_AWADDR,
    output wire [7:0]                      M_AXIMM_10_AWLEN,
    output wire [2:0]                      M_AXIMM_10_AWSIZE,
    output wire [1:0]                      M_AXIMM_10_AWBURST,
    output wire [1:0]                      M_AXIMM_10_AWLOCK,
    output wire [3:0]                      M_AXIMM_10_AWCACHE,
    output wire [2:0]                      M_AXIMM_10_AWPROT,
    output wire [3:0]                      M_AXIMM_10_AWREGION,
    output wire [3:0]                      M_AXIMM_10_AWQOS,
    output wire                            M_AXIMM_10_AWVALID,
    input  wire                            M_AXIMM_10_AWREADY,
    output wire [M_AXIMM_10_DATA_WIDTH-1:0]   M_AXIMM_10_WDATA,
    output wire [M_AXIMM_10_DATA_WIDTH/8-1:0] M_AXIMM_10_WSTRB,
    output wire                            M_AXIMM_10_WLAST,
    output wire                            M_AXIMM_10_WVALID,
    input  wire                            M_AXIMM_10_WREADY,
    input  wire [1:0]                      M_AXIMM_10_BRESP,
    input  wire                            M_AXIMM_10_BVALID,
    output wire                            M_AXIMM_10_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_10_ARADDR,
    output wire [7:0]                      M_AXIMM_10_ARLEN,
    output wire [2:0]                      M_AXIMM_10_ARSIZE,
    output wire [1:0]                      M_AXIMM_10_ARBURST,
    output wire [1:0]                      M_AXIMM_10_ARLOCK,
    output wire [3:0]                      M_AXIMM_10_ARCACHE,
    output wire [2:0]                      M_AXIMM_10_ARPROT,
    output wire [3:0]                      M_AXIMM_10_ARREGION,
    output wire [3:0]                      M_AXIMM_10_ARQOS,
    output wire                            M_AXIMM_10_ARVALID,
    input  wire                            M_AXIMM_10_ARREADY,
    input  wire [M_AXIMM_10_DATA_WIDTH-1:0]   M_AXIMM_10_RDATA,
    input  wire [1:0]                      M_AXIMM_10_RRESP,
    input  wire                            M_AXIMM_10_RLAST,
    input  wire                            M_AXIMM_10_RVALID,
    output wire                            M_AXIMM_10_RREADY,
    //AXI-MM pass-through interface 11
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_11_AWADDR,
    input wire [7:0]                      AP_AXIMM_11_AWLEN,
    input wire [2:0]                      AP_AXIMM_11_AWSIZE,
    input wire [1:0]                      AP_AXIMM_11_AWBURST,
    input wire [1:0]                      AP_AXIMM_11_AWLOCK,
    input wire [3:0]                      AP_AXIMM_11_AWCACHE,
    input wire [2:0]                      AP_AXIMM_11_AWPROT,
    input wire [3:0]                      AP_AXIMM_11_AWREGION,
    input wire [3:0]                      AP_AXIMM_11_AWQOS,
    input wire                            AP_AXIMM_11_AWVALID,
    output  wire                            AP_AXIMM_11_AWREADY,
    input wire [M_AXIMM_11_DATA_WIDTH-1:0]   AP_AXIMM_11_WDATA,
    input wire [M_AXIMM_11_DATA_WIDTH/8-1:0] AP_AXIMM_11_WSTRB,
    input wire                            AP_AXIMM_11_WLAST,
    input wire                            AP_AXIMM_11_WVALID,
    output  wire                            AP_AXIMM_11_WREADY,
    output  wire [1:0]                      AP_AXIMM_11_BRESP,
    output  wire                            AP_AXIMM_11_BVALID,
    input wire                            AP_AXIMM_11_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_11_ARADDR,
    input wire [7:0]                      AP_AXIMM_11_ARLEN,
    input wire [2:0]                      AP_AXIMM_11_ARSIZE,
    input wire [1:0]                      AP_AXIMM_11_ARBURST,
    input wire [1:0]                      AP_AXIMM_11_ARLOCK,
    input wire [3:0]                      AP_AXIMM_11_ARCACHE,
    input wire [2:0]                      AP_AXIMM_11_ARPROT,
    input wire [3:0]                      AP_AXIMM_11_ARREGION,
    input wire [3:0]                      AP_AXIMM_11_ARQOS,
    input wire                            AP_AXIMM_11_ARVALID,
    output  wire                            AP_AXIMM_11_ARREADY,
    output  wire [M_AXIMM_11_DATA_WIDTH-1:0]   AP_AXIMM_11_RDATA,
    output  wire [1:0]                      AP_AXIMM_11_RRESP,
    output  wire                            AP_AXIMM_11_RLAST,
    output  wire                            AP_AXIMM_11_RVALID,
    input  wire                            AP_AXIMM_11_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_11_AWADDR,
    output wire [7:0]                      M_AXIMM_11_AWLEN,
    output wire [2:0]                      M_AXIMM_11_AWSIZE,
    output wire [1:0]                      M_AXIMM_11_AWBURST,
    output wire [1:0]                      M_AXIMM_11_AWLOCK,
    output wire [3:0]                      M_AXIMM_11_AWCACHE,
    output wire [2:0]                      M_AXIMM_11_AWPROT,
    output wire [3:0]                      M_AXIMM_11_AWREGION,
    output wire [3:0]                      M_AXIMM_11_AWQOS,
    output wire                            M_AXIMM_11_AWVALID,
    input  wire                            M_AXIMM_11_AWREADY,
    output wire [M_AXIMM_11_DATA_WIDTH-1:0]   M_AXIMM_11_WDATA,
    output wire [M_AXIMM_11_DATA_WIDTH/8-1:0] M_AXIMM_11_WSTRB,
    output wire                            M_AXIMM_11_WLAST,
    output wire                            M_AXIMM_11_WVALID,
    input  wire                            M_AXIMM_11_WREADY,
    input  wire [1:0]                      M_AXIMM_11_BRESP,
    input  wire                            M_AXIMM_11_BVALID,
    output wire                            M_AXIMM_11_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_11_ARADDR,
    output wire [7:0]                      M_AXIMM_11_ARLEN,
    output wire [2:0]                      M_AXIMM_11_ARSIZE,
    output wire [1:0]                      M_AXIMM_11_ARBURST,
    output wire [1:0]                      M_AXIMM_11_ARLOCK,
    output wire [3:0]                      M_AXIMM_11_ARCACHE,
    output wire [2:0]                      M_AXIMM_11_ARPROT,
    output wire [3:0]                      M_AXIMM_11_ARREGION,
    output wire [3:0]                      M_AXIMM_11_ARQOS,
    output wire                            M_AXIMM_11_ARVALID,
    input  wire                            M_AXIMM_11_ARREADY,
    input  wire [M_AXIMM_11_DATA_WIDTH-1:0]   M_AXIMM_11_RDATA,
    input  wire [1:0]                      M_AXIMM_11_RRESP,
    input  wire                            M_AXIMM_11_RLAST,
    input  wire                            M_AXIMM_11_RVALID,
    output wire                            M_AXIMM_11_RREADY,
    //AXI-MM pass-through interface 12
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_12_AWADDR,
    input wire [7:0]                      AP_AXIMM_12_AWLEN,
    input wire [2:0]                      AP_AXIMM_12_AWSIZE,
    input wire [1:0]                      AP_AXIMM_12_AWBURST,
    input wire [1:0]                      AP_AXIMM_12_AWLOCK,
    input wire [3:0]                      AP_AXIMM_12_AWCACHE,
    input wire [2:0]                      AP_AXIMM_12_AWPROT,
    input wire [3:0]                      AP_AXIMM_12_AWREGION,
    input wire [3:0]                      AP_AXIMM_12_AWQOS,
    input wire                            AP_AXIMM_12_AWVALID,
    output  wire                            AP_AXIMM_12_AWREADY,
    input wire [M_AXIMM_12_DATA_WIDTH-1:0]   AP_AXIMM_12_WDATA,
    input wire [M_AXIMM_12_DATA_WIDTH/8-1:0] AP_AXIMM_12_WSTRB,
    input wire                            AP_AXIMM_12_WLAST,
    input wire                            AP_AXIMM_12_WVALID,
    output  wire                            AP_AXIMM_12_WREADY,
    output  wire [1:0]                      AP_AXIMM_12_BRESP,
    output  wire                            AP_AXIMM_12_BVALID,
    input wire                            AP_AXIMM_12_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_12_ARADDR,
    input wire [7:0]                      AP_AXIMM_12_ARLEN,
    input wire [2:0]                      AP_AXIMM_12_ARSIZE,
    input wire [1:0]                      AP_AXIMM_12_ARBURST,
    input wire [1:0]                      AP_AXIMM_12_ARLOCK,
    input wire [3:0]                      AP_AXIMM_12_ARCACHE,
    input wire [2:0]                      AP_AXIMM_12_ARPROT,
    input wire [3:0]                      AP_AXIMM_12_ARREGION,
    input wire [3:0]                      AP_AXIMM_12_ARQOS,
    input wire                            AP_AXIMM_12_ARVALID,
    output  wire                            AP_AXIMM_12_ARREADY,
    output  wire [M_AXIMM_12_DATA_WIDTH-1:0]   AP_AXIMM_12_RDATA,
    output  wire [1:0]                      AP_AXIMM_12_RRESP,
    output  wire                            AP_AXIMM_12_RLAST,
    output  wire                            AP_AXIMM_12_RVALID,
    input  wire                            AP_AXIMM_12_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_12_AWADDR,
    output wire [7:0]                      M_AXIMM_12_AWLEN,
    output wire [2:0]                      M_AXIMM_12_AWSIZE,
    output wire [1:0]                      M_AXIMM_12_AWBURST,
    output wire [1:0]                      M_AXIMM_12_AWLOCK,
    output wire [3:0]                      M_AXIMM_12_AWCACHE,
    output wire [2:0]                      M_AXIMM_12_AWPROT,
    output wire [3:0]                      M_AXIMM_12_AWREGION,
    output wire [3:0]                      M_AXIMM_12_AWQOS,
    output wire                            M_AXIMM_12_AWVALID,
    input  wire                            M_AXIMM_12_AWREADY,
    output wire [M_AXIMM_12_DATA_WIDTH-1:0]   M_AXIMM_12_WDATA,
    output wire [M_AXIMM_12_DATA_WIDTH/8-1:0] M_AXIMM_12_WSTRB,
    output wire                            M_AXIMM_12_WLAST,
    output wire                            M_AXIMM_12_WVALID,
    input  wire                            M_AXIMM_12_WREADY,
    input  wire [1:0]                      M_AXIMM_12_BRESP,
    input  wire                            M_AXIMM_12_BVALID,
    output wire                            M_AXIMM_12_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_12_ARADDR,
    output wire [7:0]                      M_AXIMM_12_ARLEN,
    output wire [2:0]                      M_AXIMM_12_ARSIZE,
    output wire [1:0]                      M_AXIMM_12_ARBURST,
    output wire [1:0]                      M_AXIMM_12_ARLOCK,
    output wire [3:0]                      M_AXIMM_12_ARCACHE,
    output wire [2:0]                      M_AXIMM_12_ARPROT,
    output wire [3:0]                      M_AXIMM_12_ARREGION,
    output wire [3:0]                      M_AXIMM_12_ARQOS,
    output wire                            M_AXIMM_12_ARVALID,
    input  wire                            M_AXIMM_12_ARREADY,
    input  wire [M_AXIMM_12_DATA_WIDTH-1:0]   M_AXIMM_12_RDATA,
    input  wire [1:0]                      M_AXIMM_12_RRESP,
    input  wire                            M_AXIMM_12_RLAST,
    input  wire                            M_AXIMM_12_RVALID,
    output wire                            M_AXIMM_12_RREADY,
    //AXI-MM pass-through interface 13
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_13_AWADDR,
    input wire [7:0]                      AP_AXIMM_13_AWLEN,
    input wire [2:0]                      AP_AXIMM_13_AWSIZE,
    input wire [1:0]                      AP_AXIMM_13_AWBURST,
    input wire [1:0]                      AP_AXIMM_13_AWLOCK,
    input wire [3:0]                      AP_AXIMM_13_AWCACHE,
    input wire [2:0]                      AP_AXIMM_13_AWPROT,
    input wire [3:0]                      AP_AXIMM_13_AWREGION,
    input wire [3:0]                      AP_AXIMM_13_AWQOS,
    input wire                            AP_AXIMM_13_AWVALID,
    output  wire                            AP_AXIMM_13_AWREADY,
    input wire [M_AXIMM_13_DATA_WIDTH-1:0]   AP_AXIMM_13_WDATA,
    input wire [M_AXIMM_13_DATA_WIDTH/8-1:0] AP_AXIMM_13_WSTRB,
    input wire                            AP_AXIMM_13_WLAST,
    input wire                            AP_AXIMM_13_WVALID,
    output  wire                            AP_AXIMM_13_WREADY,
    output  wire [1:0]                      AP_AXIMM_13_BRESP,
    output  wire                            AP_AXIMM_13_BVALID,
    input wire                            AP_AXIMM_13_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_13_ARADDR,
    input wire [7:0]                      AP_AXIMM_13_ARLEN,
    input wire [2:0]                      AP_AXIMM_13_ARSIZE,
    input wire [1:0]                      AP_AXIMM_13_ARBURST,
    input wire [1:0]                      AP_AXIMM_13_ARLOCK,
    input wire [3:0]                      AP_AXIMM_13_ARCACHE,
    input wire [2:0]                      AP_AXIMM_13_ARPROT,
    input wire [3:0]                      AP_AXIMM_13_ARREGION,
    input wire [3:0]                      AP_AXIMM_13_ARQOS,
    input wire                            AP_AXIMM_13_ARVALID,
    output  wire                            AP_AXIMM_13_ARREADY,
    output  wire [M_AXIMM_13_DATA_WIDTH-1:0]   AP_AXIMM_13_RDATA,
    output  wire [1:0]                      AP_AXIMM_13_RRESP,
    output  wire                            AP_AXIMM_13_RLAST,
    output  wire                            AP_AXIMM_13_RVALID,
    input  wire                            AP_AXIMM_13_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_13_AWADDR,
    output wire [7:0]                      M_AXIMM_13_AWLEN,
    output wire [2:0]                      M_AXIMM_13_AWSIZE,
    output wire [1:0]                      M_AXIMM_13_AWBURST,
    output wire [1:0]                      M_AXIMM_13_AWLOCK,
    output wire [3:0]                      M_AXIMM_13_AWCACHE,
    output wire [2:0]                      M_AXIMM_13_AWPROT,
    output wire [3:0]                      M_AXIMM_13_AWREGION,
    output wire [3:0]                      M_AXIMM_13_AWQOS,
    output wire                            M_AXIMM_13_AWVALID,
    input  wire                            M_AXIMM_13_AWREADY,
    output wire [M_AXIMM_13_DATA_WIDTH-1:0]   M_AXIMM_13_WDATA,
    output wire [M_AXIMM_13_DATA_WIDTH/8-1:0] M_AXIMM_13_WSTRB,
    output wire                            M_AXIMM_13_WLAST,
    output wire                            M_AXIMM_13_WVALID,
    input  wire                            M_AXIMM_13_WREADY,
    input  wire [1:0]                      M_AXIMM_13_BRESP,
    input  wire                            M_AXIMM_13_BVALID,
    output wire                            M_AXIMM_13_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_13_ARADDR,
    output wire [7:0]                      M_AXIMM_13_ARLEN,
    output wire [2:0]                      M_AXIMM_13_ARSIZE,
    output wire [1:0]                      M_AXIMM_13_ARBURST,
    output wire [1:0]                      M_AXIMM_13_ARLOCK,
    output wire [3:0]                      M_AXIMM_13_ARCACHE,
    output wire [2:0]                      M_AXIMM_13_ARPROT,
    output wire [3:0]                      M_AXIMM_13_ARREGION,
    output wire [3:0]                      M_AXIMM_13_ARQOS,
    output wire                            M_AXIMM_13_ARVALID,
    input  wire                            M_AXIMM_13_ARREADY,
    input  wire [M_AXIMM_13_DATA_WIDTH-1:0]   M_AXIMM_13_RDATA,
    input  wire [1:0]                      M_AXIMM_13_RRESP,
    input  wire                            M_AXIMM_13_RLAST,
    input  wire                            M_AXIMM_13_RVALID,
    output wire                            M_AXIMM_13_RREADY,
    //AXI-MM pass-through interface 14
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_14_AWADDR,
    input wire [7:0]                      AP_AXIMM_14_AWLEN,
    input wire [2:0]                      AP_AXIMM_14_AWSIZE,
    input wire [1:0]                      AP_AXIMM_14_AWBURST,
    input wire [1:0]                      AP_AXIMM_14_AWLOCK,
    input wire [3:0]                      AP_AXIMM_14_AWCACHE,
    input wire [2:0]                      AP_AXIMM_14_AWPROT,
    input wire [3:0]                      AP_AXIMM_14_AWREGION,
    input wire [3:0]                      AP_AXIMM_14_AWQOS,
    input wire                            AP_AXIMM_14_AWVALID,
    output  wire                            AP_AXIMM_14_AWREADY,
    input wire [M_AXIMM_14_DATA_WIDTH-1:0]   AP_AXIMM_14_WDATA,
    input wire [M_AXIMM_14_DATA_WIDTH/8-1:0] AP_AXIMM_14_WSTRB,
    input wire                            AP_AXIMM_14_WLAST,
    input wire                            AP_AXIMM_14_WVALID,
    output  wire                            AP_AXIMM_14_WREADY,
    output  wire [1:0]                      AP_AXIMM_14_BRESP,
    output  wire                            AP_AXIMM_14_BVALID,
    input wire                            AP_AXIMM_14_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_14_ARADDR,
    input wire [7:0]                      AP_AXIMM_14_ARLEN,
    input wire [2:0]                      AP_AXIMM_14_ARSIZE,
    input wire [1:0]                      AP_AXIMM_14_ARBURST,
    input wire [1:0]                      AP_AXIMM_14_ARLOCK,
    input wire [3:0]                      AP_AXIMM_14_ARCACHE,
    input wire [2:0]                      AP_AXIMM_14_ARPROT,
    input wire [3:0]                      AP_AXIMM_14_ARREGION,
    input wire [3:0]                      AP_AXIMM_14_ARQOS,
    input wire                            AP_AXIMM_14_ARVALID,
    output  wire                            AP_AXIMM_14_ARREADY,
    output  wire [M_AXIMM_14_DATA_WIDTH-1:0]   AP_AXIMM_14_RDATA,
    output  wire [1:0]                      AP_AXIMM_14_RRESP,
    output  wire                            AP_AXIMM_14_RLAST,
    output  wire                            AP_AXIMM_14_RVALID,
    input  wire                            AP_AXIMM_14_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_14_AWADDR,
    output wire [7:0]                      M_AXIMM_14_AWLEN,
    output wire [2:0]                      M_AXIMM_14_AWSIZE,
    output wire [1:0]                      M_AXIMM_14_AWBURST,
    output wire [1:0]                      M_AXIMM_14_AWLOCK,
    output wire [3:0]                      M_AXIMM_14_AWCACHE,
    output wire [2:0]                      M_AXIMM_14_AWPROT,
    output wire [3:0]                      M_AXIMM_14_AWREGION,
    output wire [3:0]                      M_AXIMM_14_AWQOS,
    output wire                            M_AXIMM_14_AWVALID,
    input  wire                            M_AXIMM_14_AWREADY,
    output wire [M_AXIMM_14_DATA_WIDTH-1:0]   M_AXIMM_14_WDATA,
    output wire [M_AXIMM_14_DATA_WIDTH/8-1:0] M_AXIMM_14_WSTRB,
    output wire                            M_AXIMM_14_WLAST,
    output wire                            M_AXIMM_14_WVALID,
    input  wire                            M_AXIMM_14_WREADY,
    input  wire [1:0]                      M_AXIMM_14_BRESP,
    input  wire                            M_AXIMM_14_BVALID,
    output wire                            M_AXIMM_14_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_14_ARADDR,
    output wire [7:0]                      M_AXIMM_14_ARLEN,
    output wire [2:0]                      M_AXIMM_14_ARSIZE,
    output wire [1:0]                      M_AXIMM_14_ARBURST,
    output wire [1:0]                      M_AXIMM_14_ARLOCK,
    output wire [3:0]                      M_AXIMM_14_ARCACHE,
    output wire [2:0]                      M_AXIMM_14_ARPROT,
    output wire [3:0]                      M_AXIMM_14_ARREGION,
    output wire [3:0]                      M_AXIMM_14_ARQOS,
    output wire                            M_AXIMM_14_ARVALID,
    input  wire                            M_AXIMM_14_ARREADY,
    input  wire [M_AXIMM_14_DATA_WIDTH-1:0]   M_AXIMM_14_RDATA,
    input  wire [1:0]                      M_AXIMM_14_RRESP,
    input  wire                            M_AXIMM_14_RLAST,
    input  wire                            M_AXIMM_14_RVALID,
    output wire                            M_AXIMM_14_RREADY,
    //AXI-MM pass-through interface 15
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_15_AWADDR,
    input wire [7:0]                      AP_AXIMM_15_AWLEN,
    input wire [2:0]                      AP_AXIMM_15_AWSIZE,
    input wire [1:0]                      AP_AXIMM_15_AWBURST,
    input wire [1:0]                      AP_AXIMM_15_AWLOCK,
    input wire [3:0]                      AP_AXIMM_15_AWCACHE,
    input wire [2:0]                      AP_AXIMM_15_AWPROT,
    input wire [3:0]                      AP_AXIMM_15_AWREGION,
    input wire [3:0]                      AP_AXIMM_15_AWQOS,
    input wire                            AP_AXIMM_15_AWVALID,
    output  wire                            AP_AXIMM_15_AWREADY,
    input wire [M_AXIMM_15_DATA_WIDTH-1:0]   AP_AXIMM_15_WDATA,
    input wire [M_AXIMM_15_DATA_WIDTH/8-1:0] AP_AXIMM_15_WSTRB,
    input wire                            AP_AXIMM_15_WLAST,
    input wire                            AP_AXIMM_15_WVALID,
    output  wire                            AP_AXIMM_15_WREADY,
    output  wire [1:0]                      AP_AXIMM_15_BRESP,
    output  wire                            AP_AXIMM_15_BVALID,
    input wire                            AP_AXIMM_15_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_15_ARADDR,
    input wire [7:0]                      AP_AXIMM_15_ARLEN,
    input wire [2:0]                      AP_AXIMM_15_ARSIZE,
    input wire [1:0]                      AP_AXIMM_15_ARBURST,
    input wire [1:0]                      AP_AXIMM_15_ARLOCK,
    input wire [3:0]                      AP_AXIMM_15_ARCACHE,
    input wire [2:0]                      AP_AXIMM_15_ARPROT,
    input wire [3:0]                      AP_AXIMM_15_ARREGION,
    input wire [3:0]                      AP_AXIMM_15_ARQOS,
    input wire                            AP_AXIMM_15_ARVALID,
    output  wire                            AP_AXIMM_15_ARREADY,
    output  wire [M_AXIMM_15_DATA_WIDTH-1:0]   AP_AXIMM_15_RDATA,
    output  wire [1:0]                      AP_AXIMM_15_RRESP,
    output  wire                            AP_AXIMM_15_RLAST,
    output  wire                            AP_AXIMM_15_RVALID,
    input  wire                            AP_AXIMM_15_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_15_AWADDR,
    output wire [7:0]                      M_AXIMM_15_AWLEN,
    output wire [2:0]                      M_AXIMM_15_AWSIZE,
    output wire [1:0]                      M_AXIMM_15_AWBURST,
    output wire [1:0]                      M_AXIMM_15_AWLOCK,
    output wire [3:0]                      M_AXIMM_15_AWCACHE,
    output wire [2:0]                      M_AXIMM_15_AWPROT,
    output wire [3:0]                      M_AXIMM_15_AWREGION,
    output wire [3:0]                      M_AXIMM_15_AWQOS,
    output wire                            M_AXIMM_15_AWVALID,
    input  wire                            M_AXIMM_15_AWREADY,
    output wire [M_AXIMM_15_DATA_WIDTH-1:0]   M_AXIMM_15_WDATA,
    output wire [M_AXIMM_15_DATA_WIDTH/8-1:0] M_AXIMM_15_WSTRB,
    output wire                            M_AXIMM_15_WLAST,
    output wire                            M_AXIMM_15_WVALID,
    input  wire                            M_AXIMM_15_WREADY,
    input  wire [1:0]                      M_AXIMM_15_BRESP,
    input  wire                            M_AXIMM_15_BVALID,
    output wire                            M_AXIMM_15_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_15_ARADDR,
    output wire [7:0]                      M_AXIMM_15_ARLEN,
    output wire [2:0]                      M_AXIMM_15_ARSIZE,
    output wire [1:0]                      M_AXIMM_15_ARBURST,
    output wire [1:0]                      M_AXIMM_15_ARLOCK,
    output wire [3:0]                      M_AXIMM_15_ARCACHE,
    output wire [2:0]                      M_AXIMM_15_ARPROT,
    output wire [3:0]                      M_AXIMM_15_ARREGION,
    output wire [3:0]                      M_AXIMM_15_ARQOS,
    output wire                            M_AXIMM_15_ARVALID,
    input  wire                            M_AXIMM_15_ARREADY,
    input  wire [M_AXIMM_15_DATA_WIDTH-1:0]   M_AXIMM_15_RDATA,
    input  wire [1:0]                      M_AXIMM_15_RRESP,
    input  wire                            M_AXIMM_15_RLAST,
    input  wire                            M_AXIMM_15_RVALID,
    output wire                            M_AXIMM_15_RREADY,
    //AXI-MM pass-through interface 16
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_16_AWADDR,
    input wire [7:0]                      AP_AXIMM_16_AWLEN,
    input wire [2:0]                      AP_AXIMM_16_AWSIZE,
    input wire [1:0]                      AP_AXIMM_16_AWBURST,
    input wire [1:0]                      AP_AXIMM_16_AWLOCK,
    input wire [3:0]                      AP_AXIMM_16_AWCACHE,
    input wire [2:0]                      AP_AXIMM_16_AWPROT,
    input wire [3:0]                      AP_AXIMM_16_AWREGION,
    input wire [3:0]                      AP_AXIMM_16_AWQOS,
    input wire                            AP_AXIMM_16_AWVALID,
    output  wire                            AP_AXIMM_16_AWREADY,
    input wire [M_AXIMM_16_DATA_WIDTH-1:0]   AP_AXIMM_16_WDATA,
    input wire [M_AXIMM_16_DATA_WIDTH/8-1:0] AP_AXIMM_16_WSTRB,
    input wire                            AP_AXIMM_16_WLAST,
    input wire                            AP_AXIMM_16_WVALID,
    output  wire                            AP_AXIMM_16_WREADY,
    output  wire [1:0]                      AP_AXIMM_16_BRESP,
    output  wire                            AP_AXIMM_16_BVALID,
    input wire                            AP_AXIMM_16_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_16_ARADDR,
    input wire [7:0]                      AP_AXIMM_16_ARLEN,
    input wire [2:0]                      AP_AXIMM_16_ARSIZE,
    input wire [1:0]                      AP_AXIMM_16_ARBURST,
    input wire [1:0]                      AP_AXIMM_16_ARLOCK,
    input wire [3:0]                      AP_AXIMM_16_ARCACHE,
    input wire [2:0]                      AP_AXIMM_16_ARPROT,
    input wire [3:0]                      AP_AXIMM_16_ARREGION,
    input wire [3:0]                      AP_AXIMM_16_ARQOS,
    input wire                            AP_AXIMM_16_ARVALID,
    output  wire                            AP_AXIMM_16_ARREADY,
    output  wire [M_AXIMM_16_DATA_WIDTH-1:0]   AP_AXIMM_16_RDATA,
    output  wire [1:0]                      AP_AXIMM_16_RRESP,
    output  wire                            AP_AXIMM_16_RLAST,
    output  wire                            AP_AXIMM_16_RVALID,
    input  wire                            AP_AXIMM_16_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_16_AWADDR,
    output wire [7:0]                      M_AXIMM_16_AWLEN,
    output wire [2:0]                      M_AXIMM_16_AWSIZE,
    output wire [1:0]                      M_AXIMM_16_AWBURST,
    output wire [1:0]                      M_AXIMM_16_AWLOCK,
    output wire [3:0]                      M_AXIMM_16_AWCACHE,
    output wire [2:0]                      M_AXIMM_16_AWPROT,
    output wire [3:0]                      M_AXIMM_16_AWREGION,
    output wire [3:0]                      M_AXIMM_16_AWQOS,
    output wire                            M_AXIMM_16_AWVALID,
    input  wire                            M_AXIMM_16_AWREADY,
    output wire [M_AXIMM_16_DATA_WIDTH-1:0]   M_AXIMM_16_WDATA,
    output wire [M_AXIMM_16_DATA_WIDTH/8-1:0] M_AXIMM_16_WSTRB,
    output wire                            M_AXIMM_16_WLAST,
    output wire                            M_AXIMM_16_WVALID,
    input  wire                            M_AXIMM_16_WREADY,
    input  wire [1:0]                      M_AXIMM_16_BRESP,
    input  wire                            M_AXIMM_16_BVALID,
    output wire                            M_AXIMM_16_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_16_ARADDR,
    output wire [7:0]                      M_AXIMM_16_ARLEN,
    output wire [2:0]                      M_AXIMM_16_ARSIZE,
    output wire [1:0]                      M_AXIMM_16_ARBURST,
    output wire [1:0]                      M_AXIMM_16_ARLOCK,
    output wire [3:0]                      M_AXIMM_16_ARCACHE,
    output wire [2:0]                      M_AXIMM_16_ARPROT,
    output wire [3:0]                      M_AXIMM_16_ARREGION,
    output wire [3:0]                      M_AXIMM_16_ARQOS,
    output wire                            M_AXIMM_16_ARVALID,
    input  wire                            M_AXIMM_16_ARREADY,
    input  wire [M_AXIMM_16_DATA_WIDTH-1:0]   M_AXIMM_16_RDATA,
    input  wire [1:0]                      M_AXIMM_16_RRESP,
    input  wire                            M_AXIMM_16_RLAST,
    input  wire                            M_AXIMM_16_RVALID,
    output wire                            M_AXIMM_16_RREADY,
    //AXI-MM pass-through interface 17
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_17_AWADDR,
    input wire [7:0]                      AP_AXIMM_17_AWLEN,
    input wire [2:0]                      AP_AXIMM_17_AWSIZE,
    input wire [1:0]                      AP_AXIMM_17_AWBURST,
    input wire [1:0]                      AP_AXIMM_17_AWLOCK,
    input wire [3:0]                      AP_AXIMM_17_AWCACHE,
    input wire [2:0]                      AP_AXIMM_17_AWPROT,
    input wire [3:0]                      AP_AXIMM_17_AWREGION,
    input wire [3:0]                      AP_AXIMM_17_AWQOS,
    input wire                            AP_AXIMM_17_AWVALID,
    output  wire                            AP_AXIMM_17_AWREADY,
    input wire [M_AXIMM_17_DATA_WIDTH-1:0]   AP_AXIMM_17_WDATA,
    input wire [M_AXIMM_17_DATA_WIDTH/8-1:0] AP_AXIMM_17_WSTRB,
    input wire                            AP_AXIMM_17_WLAST,
    input wire                            AP_AXIMM_17_WVALID,
    output  wire                            AP_AXIMM_17_WREADY,
    output  wire [1:0]                      AP_AXIMM_17_BRESP,
    output  wire                            AP_AXIMM_17_BVALID,
    input wire                            AP_AXIMM_17_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_17_ARADDR,
    input wire [7:0]                      AP_AXIMM_17_ARLEN,
    input wire [2:0]                      AP_AXIMM_17_ARSIZE,
    input wire [1:0]                      AP_AXIMM_17_ARBURST,
    input wire [1:0]                      AP_AXIMM_17_ARLOCK,
    input wire [3:0]                      AP_AXIMM_17_ARCACHE,
    input wire [2:0]                      AP_AXIMM_17_ARPROT,
    input wire [3:0]                      AP_AXIMM_17_ARREGION,
    input wire [3:0]                      AP_AXIMM_17_ARQOS,
    input wire                            AP_AXIMM_17_ARVALID,
    output  wire                            AP_AXIMM_17_ARREADY,
    output  wire [M_AXIMM_17_DATA_WIDTH-1:0]   AP_AXIMM_17_RDATA,
    output  wire [1:0]                      AP_AXIMM_17_RRESP,
    output  wire                            AP_AXIMM_17_RLAST,
    output  wire                            AP_AXIMM_17_RVALID,
    input  wire                            AP_AXIMM_17_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_17_AWADDR,
    output wire [7:0]                      M_AXIMM_17_AWLEN,
    output wire [2:0]                      M_AXIMM_17_AWSIZE,
    output wire [1:0]                      M_AXIMM_17_AWBURST,
    output wire [1:0]                      M_AXIMM_17_AWLOCK,
    output wire [3:0]                      M_AXIMM_17_AWCACHE,
    output wire [2:0]                      M_AXIMM_17_AWPROT,
    output wire [3:0]                      M_AXIMM_17_AWREGION,
    output wire [3:0]                      M_AXIMM_17_AWQOS,
    output wire                            M_AXIMM_17_AWVALID,
    input  wire                            M_AXIMM_17_AWREADY,
    output wire [M_AXIMM_17_DATA_WIDTH-1:0]   M_AXIMM_17_WDATA,
    output wire [M_AXIMM_17_DATA_WIDTH/8-1:0] M_AXIMM_17_WSTRB,
    output wire                            M_AXIMM_17_WLAST,
    output wire                            M_AXIMM_17_WVALID,
    input  wire                            M_AXIMM_17_WREADY,
    input  wire [1:0]                      M_AXIMM_17_BRESP,
    input  wire                            M_AXIMM_17_BVALID,
    output wire                            M_AXIMM_17_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_17_ARADDR,
    output wire [7:0]                      M_AXIMM_17_ARLEN,
    output wire [2:0]                      M_AXIMM_17_ARSIZE,
    output wire [1:0]                      M_AXIMM_17_ARBURST,
    output wire [1:0]                      M_AXIMM_17_ARLOCK,
    output wire [3:0]                      M_AXIMM_17_ARCACHE,
    output wire [2:0]                      M_AXIMM_17_ARPROT,
    output wire [3:0]                      M_AXIMM_17_ARREGION,
    output wire [3:0]                      M_AXIMM_17_ARQOS,
    output wire                            M_AXIMM_17_ARVALID,
    input  wire                            M_AXIMM_17_ARREADY,
    input  wire [M_AXIMM_17_DATA_WIDTH-1:0]   M_AXIMM_17_RDATA,
    input  wire [1:0]                      M_AXIMM_17_RRESP,
    input  wire                            M_AXIMM_17_RLAST,
    input  wire                            M_AXIMM_17_RVALID,
    output wire                            M_AXIMM_17_RREADY,
    //AXI-MM pass-through interface 18
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_18_AWADDR,
    input wire [7:0]                      AP_AXIMM_18_AWLEN,
    input wire [2:0]                      AP_AXIMM_18_AWSIZE,
    input wire [1:0]                      AP_AXIMM_18_AWBURST,
    input wire [1:0]                      AP_AXIMM_18_AWLOCK,
    input wire [3:0]                      AP_AXIMM_18_AWCACHE,
    input wire [2:0]                      AP_AXIMM_18_AWPROT,
    input wire [3:0]                      AP_AXIMM_18_AWREGION,
    input wire [3:0]                      AP_AXIMM_18_AWQOS,
    input wire                            AP_AXIMM_18_AWVALID,
    output  wire                            AP_AXIMM_18_AWREADY,
    input wire [M_AXIMM_18_DATA_WIDTH-1:0]   AP_AXIMM_18_WDATA,
    input wire [M_AXIMM_18_DATA_WIDTH/8-1:0] AP_AXIMM_18_WSTRB,
    input wire                            AP_AXIMM_18_WLAST,
    input wire                            AP_AXIMM_18_WVALID,
    output  wire                            AP_AXIMM_18_WREADY,
    output  wire [1:0]                      AP_AXIMM_18_BRESP,
    output  wire                            AP_AXIMM_18_BVALID,
    input wire                            AP_AXIMM_18_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_18_ARADDR,
    input wire [7:0]                      AP_AXIMM_18_ARLEN,
    input wire [2:0]                      AP_AXIMM_18_ARSIZE,
    input wire [1:0]                      AP_AXIMM_18_ARBURST,
    input wire [1:0]                      AP_AXIMM_18_ARLOCK,
    input wire [3:0]                      AP_AXIMM_18_ARCACHE,
    input wire [2:0]                      AP_AXIMM_18_ARPROT,
    input wire [3:0]                      AP_AXIMM_18_ARREGION,
    input wire [3:0]                      AP_AXIMM_18_ARQOS,
    input wire                            AP_AXIMM_18_ARVALID,
    output  wire                            AP_AXIMM_18_ARREADY,
    output  wire [M_AXIMM_18_DATA_WIDTH-1:0]   AP_AXIMM_18_RDATA,
    output  wire [1:0]                      AP_AXIMM_18_RRESP,
    output  wire                            AP_AXIMM_18_RLAST,
    output  wire                            AP_AXIMM_18_RVALID,
    input  wire                            AP_AXIMM_18_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_18_AWADDR,
    output wire [7:0]                      M_AXIMM_18_AWLEN,
    output wire [2:0]                      M_AXIMM_18_AWSIZE,
    output wire [1:0]                      M_AXIMM_18_AWBURST,
    output wire [1:0]                      M_AXIMM_18_AWLOCK,
    output wire [3:0]                      M_AXIMM_18_AWCACHE,
    output wire [2:0]                      M_AXIMM_18_AWPROT,
    output wire [3:0]                      M_AXIMM_18_AWREGION,
    output wire [3:0]                      M_AXIMM_18_AWQOS,
    output wire                            M_AXIMM_18_AWVALID,
    input  wire                            M_AXIMM_18_AWREADY,
    output wire [M_AXIMM_18_DATA_WIDTH-1:0]   M_AXIMM_18_WDATA,
    output wire [M_AXIMM_18_DATA_WIDTH/8-1:0] M_AXIMM_18_WSTRB,
    output wire                            M_AXIMM_18_WLAST,
    output wire                            M_AXIMM_18_WVALID,
    input  wire                            M_AXIMM_18_WREADY,
    input  wire [1:0]                      M_AXIMM_18_BRESP,
    input  wire                            M_AXIMM_18_BVALID,
    output wire                            M_AXIMM_18_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_18_ARADDR,
    output wire [7:0]                      M_AXIMM_18_ARLEN,
    output wire [2:0]                      M_AXIMM_18_ARSIZE,
    output wire [1:0]                      M_AXIMM_18_ARBURST,
    output wire [1:0]                      M_AXIMM_18_ARLOCK,
    output wire [3:0]                      M_AXIMM_18_ARCACHE,
    output wire [2:0]                      M_AXIMM_18_ARPROT,
    output wire [3:0]                      M_AXIMM_18_ARREGION,
    output wire [3:0]                      M_AXIMM_18_ARQOS,
    output wire                            M_AXIMM_18_ARVALID,
    input  wire                            M_AXIMM_18_ARREADY,
    input  wire [M_AXIMM_18_DATA_WIDTH-1:0]   M_AXIMM_18_RDATA,
    input  wire [1:0]                      M_AXIMM_18_RRESP,
    input  wire                            M_AXIMM_18_RLAST,
    input  wire                            M_AXIMM_18_RVALID,
    output wire                            M_AXIMM_18_RREADY,
    //AXI-MM pass-through interface 19
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_19_AWADDR,
    input wire [7:0]                      AP_AXIMM_19_AWLEN,
    input wire [2:0]                      AP_AXIMM_19_AWSIZE,
    input wire [1:0]                      AP_AXIMM_19_AWBURST,
    input wire [1:0]                      AP_AXIMM_19_AWLOCK,
    input wire [3:0]                      AP_AXIMM_19_AWCACHE,
    input wire [2:0]                      AP_AXIMM_19_AWPROT,
    input wire [3:0]                      AP_AXIMM_19_AWREGION,
    input wire [3:0]                      AP_AXIMM_19_AWQOS,
    input wire                            AP_AXIMM_19_AWVALID,
    output  wire                            AP_AXIMM_19_AWREADY,
    input wire [M_AXIMM_19_DATA_WIDTH-1:0]   AP_AXIMM_19_WDATA,
    input wire [M_AXIMM_19_DATA_WIDTH/8-1:0] AP_AXIMM_19_WSTRB,
    input wire                            AP_AXIMM_19_WLAST,
    input wire                            AP_AXIMM_19_WVALID,
    output  wire                            AP_AXIMM_19_WREADY,
    output  wire [1:0]                      AP_AXIMM_19_BRESP,
    output  wire                            AP_AXIMM_19_BVALID,
    input wire                            AP_AXIMM_19_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_19_ARADDR,
    input wire [7:0]                      AP_AXIMM_19_ARLEN,
    input wire [2:0]                      AP_AXIMM_19_ARSIZE,
    input wire [1:0]                      AP_AXIMM_19_ARBURST,
    input wire [1:0]                      AP_AXIMM_19_ARLOCK,
    input wire [3:0]                      AP_AXIMM_19_ARCACHE,
    input wire [2:0]                      AP_AXIMM_19_ARPROT,
    input wire [3:0]                      AP_AXIMM_19_ARREGION,
    input wire [3:0]                      AP_AXIMM_19_ARQOS,
    input wire                            AP_AXIMM_19_ARVALID,
    output  wire                            AP_AXIMM_19_ARREADY,
    output  wire [M_AXIMM_19_DATA_WIDTH-1:0]   AP_AXIMM_19_RDATA,
    output  wire [1:0]                      AP_AXIMM_19_RRESP,
    output  wire                            AP_AXIMM_19_RLAST,
    output  wire                            AP_AXIMM_19_RVALID,
    input  wire                            AP_AXIMM_19_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_19_AWADDR,
    output wire [7:0]                      M_AXIMM_19_AWLEN,
    output wire [2:0]                      M_AXIMM_19_AWSIZE,
    output wire [1:0]                      M_AXIMM_19_AWBURST,
    output wire [1:0]                      M_AXIMM_19_AWLOCK,
    output wire [3:0]                      M_AXIMM_19_AWCACHE,
    output wire [2:0]                      M_AXIMM_19_AWPROT,
    output wire [3:0]                      M_AXIMM_19_AWREGION,
    output wire [3:0]                      M_AXIMM_19_AWQOS,
    output wire                            M_AXIMM_19_AWVALID,
    input  wire                            M_AXIMM_19_AWREADY,
    output wire [M_AXIMM_19_DATA_WIDTH-1:0]   M_AXIMM_19_WDATA,
    output wire [M_AXIMM_19_DATA_WIDTH/8-1:0] M_AXIMM_19_WSTRB,
    output wire                            M_AXIMM_19_WLAST,
    output wire                            M_AXIMM_19_WVALID,
    input  wire                            M_AXIMM_19_WREADY,
    input  wire [1:0]                      M_AXIMM_19_BRESP,
    input  wire                            M_AXIMM_19_BVALID,
    output wire                            M_AXIMM_19_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_19_ARADDR,
    output wire [7:0]                      M_AXIMM_19_ARLEN,
    output wire [2:0]                      M_AXIMM_19_ARSIZE,
    output wire [1:0]                      M_AXIMM_19_ARBURST,
    output wire [1:0]                      M_AXIMM_19_ARLOCK,
    output wire [3:0]                      M_AXIMM_19_ARCACHE,
    output wire [2:0]                      M_AXIMM_19_ARPROT,
    output wire [3:0]                      M_AXIMM_19_ARREGION,
    output wire [3:0]                      M_AXIMM_19_ARQOS,
    output wire                            M_AXIMM_19_ARVALID,
    input  wire                            M_AXIMM_19_ARREADY,
    input  wire [M_AXIMM_19_DATA_WIDTH-1:0]   M_AXIMM_19_RDATA,
    input  wire [1:0]                      M_AXIMM_19_RRESP,
    input  wire                            M_AXIMM_19_RLAST,
    input  wire                            M_AXIMM_19_RVALID,
    output wire                            M_AXIMM_19_RREADY,
    //AXI-MM pass-through interface 20
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_20_AWADDR,
    input wire [7:0]                      AP_AXIMM_20_AWLEN,
    input wire [2:0]                      AP_AXIMM_20_AWSIZE,
    input wire [1:0]                      AP_AXIMM_20_AWBURST,
    input wire [1:0]                      AP_AXIMM_20_AWLOCK,
    input wire [3:0]                      AP_AXIMM_20_AWCACHE,
    input wire [2:0]                      AP_AXIMM_20_AWPROT,
    input wire [3:0]                      AP_AXIMM_20_AWREGION,
    input wire [3:0]                      AP_AXIMM_20_AWQOS,
    input wire                            AP_AXIMM_20_AWVALID,
    output  wire                            AP_AXIMM_20_AWREADY,
    input wire [M_AXIMM_20_DATA_WIDTH-1:0]   AP_AXIMM_20_WDATA,
    input wire [M_AXIMM_20_DATA_WIDTH/8-1:0] AP_AXIMM_20_WSTRB,
    input wire                            AP_AXIMM_20_WLAST,
    input wire                            AP_AXIMM_20_WVALID,
    output  wire                            AP_AXIMM_20_WREADY,
    output  wire [1:0]                      AP_AXIMM_20_BRESP,
    output  wire                            AP_AXIMM_20_BVALID,
    input wire                            AP_AXIMM_20_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_20_ARADDR,
    input wire [7:0]                      AP_AXIMM_20_ARLEN,
    input wire [2:0]                      AP_AXIMM_20_ARSIZE,
    input wire [1:0]                      AP_AXIMM_20_ARBURST,
    input wire [1:0]                      AP_AXIMM_20_ARLOCK,
    input wire [3:0]                      AP_AXIMM_20_ARCACHE,
    input wire [2:0]                      AP_AXIMM_20_ARPROT,
    input wire [3:0]                      AP_AXIMM_20_ARREGION,
    input wire [3:0]                      AP_AXIMM_20_ARQOS,
    input wire                            AP_AXIMM_20_ARVALID,
    output  wire                            AP_AXIMM_20_ARREADY,
    output  wire [M_AXIMM_20_DATA_WIDTH-1:0]   AP_AXIMM_20_RDATA,
    output  wire [1:0]                      AP_AXIMM_20_RRESP,
    output  wire                            AP_AXIMM_20_RLAST,
    output  wire                            AP_AXIMM_20_RVALID,
    input  wire                            AP_AXIMM_20_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_20_AWADDR,
    output wire [7:0]                      M_AXIMM_20_AWLEN,
    output wire [2:0]                      M_AXIMM_20_AWSIZE,
    output wire [1:0]                      M_AXIMM_20_AWBURST,
    output wire [1:0]                      M_AXIMM_20_AWLOCK,
    output wire [3:0]                      M_AXIMM_20_AWCACHE,
    output wire [2:0]                      M_AXIMM_20_AWPROT,
    output wire [3:0]                      M_AXIMM_20_AWREGION,
    output wire [3:0]                      M_AXIMM_20_AWQOS,
    output wire                            M_AXIMM_20_AWVALID,
    input  wire                            M_AXIMM_20_AWREADY,
    output wire [M_AXIMM_20_DATA_WIDTH-1:0]   M_AXIMM_20_WDATA,
    output wire [M_AXIMM_20_DATA_WIDTH/8-1:0] M_AXIMM_20_WSTRB,
    output wire                            M_AXIMM_20_WLAST,
    output wire                            M_AXIMM_20_WVALID,
    input  wire                            M_AXIMM_20_WREADY,
    input  wire [1:0]                      M_AXIMM_20_BRESP,
    input  wire                            M_AXIMM_20_BVALID,
    output wire                            M_AXIMM_20_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_20_ARADDR,
    output wire [7:0]                      M_AXIMM_20_ARLEN,
    output wire [2:0]                      M_AXIMM_20_ARSIZE,
    output wire [1:0]                      M_AXIMM_20_ARBURST,
    output wire [1:0]                      M_AXIMM_20_ARLOCK,
    output wire [3:0]                      M_AXIMM_20_ARCACHE,
    output wire [2:0]                      M_AXIMM_20_ARPROT,
    output wire [3:0]                      M_AXIMM_20_ARREGION,
    output wire [3:0]                      M_AXIMM_20_ARQOS,
    output wire                            M_AXIMM_20_ARVALID,
    input  wire                            M_AXIMM_20_ARREADY,
    input  wire [M_AXIMM_20_DATA_WIDTH-1:0]   M_AXIMM_20_RDATA,
    input  wire [1:0]                      M_AXIMM_20_RRESP,
    input  wire                            M_AXIMM_20_RLAST,
    input  wire                            M_AXIMM_20_RVALID,
    output wire                            M_AXIMM_20_RREADY,
    //AXI-MM pass-through interface 21
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_21_AWADDR,
    input wire [7:0]                      AP_AXIMM_21_AWLEN,
    input wire [2:0]                      AP_AXIMM_21_AWSIZE,
    input wire [1:0]                      AP_AXIMM_21_AWBURST,
    input wire [1:0]                      AP_AXIMM_21_AWLOCK,
    input wire [3:0]                      AP_AXIMM_21_AWCACHE,
    input wire [2:0]                      AP_AXIMM_21_AWPROT,
    input wire [3:0]                      AP_AXIMM_21_AWREGION,
    input wire [3:0]                      AP_AXIMM_21_AWQOS,
    input wire                            AP_AXIMM_21_AWVALID,
    output  wire                            AP_AXIMM_21_AWREADY,
    input wire [M_AXIMM_21_DATA_WIDTH-1:0]   AP_AXIMM_21_WDATA,
    input wire [M_AXIMM_21_DATA_WIDTH/8-1:0] AP_AXIMM_21_WSTRB,
    input wire                            AP_AXIMM_21_WLAST,
    input wire                            AP_AXIMM_21_WVALID,
    output  wire                            AP_AXIMM_21_WREADY,
    output  wire [1:0]                      AP_AXIMM_21_BRESP,
    output  wire                            AP_AXIMM_21_BVALID,
    input wire                            AP_AXIMM_21_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_21_ARADDR,
    input wire [7:0]                      AP_AXIMM_21_ARLEN,
    input wire [2:0]                      AP_AXIMM_21_ARSIZE,
    input wire [1:0]                      AP_AXIMM_21_ARBURST,
    input wire [1:0]                      AP_AXIMM_21_ARLOCK,
    input wire [3:0]                      AP_AXIMM_21_ARCACHE,
    input wire [2:0]                      AP_AXIMM_21_ARPROT,
    input wire [3:0]                      AP_AXIMM_21_ARREGION,
    input wire [3:0]                      AP_AXIMM_21_ARQOS,
    input wire                            AP_AXIMM_21_ARVALID,
    output  wire                            AP_AXIMM_21_ARREADY,
    output  wire [M_AXIMM_21_DATA_WIDTH-1:0]   AP_AXIMM_21_RDATA,
    output  wire [1:0]                      AP_AXIMM_21_RRESP,
    output  wire                            AP_AXIMM_21_RLAST,
    output  wire                            AP_AXIMM_21_RVALID,
    input  wire                            AP_AXIMM_21_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_21_AWADDR,
    output wire [7:0]                      M_AXIMM_21_AWLEN,
    output wire [2:0]                      M_AXIMM_21_AWSIZE,
    output wire [1:0]                      M_AXIMM_21_AWBURST,
    output wire [1:0]                      M_AXIMM_21_AWLOCK,
    output wire [3:0]                      M_AXIMM_21_AWCACHE,
    output wire [2:0]                      M_AXIMM_21_AWPROT,
    output wire [3:0]                      M_AXIMM_21_AWREGION,
    output wire [3:0]                      M_AXIMM_21_AWQOS,
    output wire                            M_AXIMM_21_AWVALID,
    input  wire                            M_AXIMM_21_AWREADY,
    output wire [M_AXIMM_21_DATA_WIDTH-1:0]   M_AXIMM_21_WDATA,
    output wire [M_AXIMM_21_DATA_WIDTH/8-1:0] M_AXIMM_21_WSTRB,
    output wire                            M_AXIMM_21_WLAST,
    output wire                            M_AXIMM_21_WVALID,
    input  wire                            M_AXIMM_21_WREADY,
    input  wire [1:0]                      M_AXIMM_21_BRESP,
    input  wire                            M_AXIMM_21_BVALID,
    output wire                            M_AXIMM_21_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_21_ARADDR,
    output wire [7:0]                      M_AXIMM_21_ARLEN,
    output wire [2:0]                      M_AXIMM_21_ARSIZE,
    output wire [1:0]                      M_AXIMM_21_ARBURST,
    output wire [1:0]                      M_AXIMM_21_ARLOCK,
    output wire [3:0]                      M_AXIMM_21_ARCACHE,
    output wire [2:0]                      M_AXIMM_21_ARPROT,
    output wire [3:0]                      M_AXIMM_21_ARREGION,
    output wire [3:0]                      M_AXIMM_21_ARQOS,
    output wire                            M_AXIMM_21_ARVALID,
    input  wire                            M_AXIMM_21_ARREADY,
    input  wire [M_AXIMM_21_DATA_WIDTH-1:0]   M_AXIMM_21_RDATA,
    input  wire [1:0]                      M_AXIMM_21_RRESP,
    input  wire                            M_AXIMM_21_RLAST,
    input  wire                            M_AXIMM_21_RVALID,
    output wire                            M_AXIMM_21_RREADY,
    //AXI-MM pass-through interface 22
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_22_AWADDR,
    input wire [7:0]                      AP_AXIMM_22_AWLEN,
    input wire [2:0]                      AP_AXIMM_22_AWSIZE,
    input wire [1:0]                      AP_AXIMM_22_AWBURST,
    input wire [1:0]                      AP_AXIMM_22_AWLOCK,
    input wire [3:0]                      AP_AXIMM_22_AWCACHE,
    input wire [2:0]                      AP_AXIMM_22_AWPROT,
    input wire [3:0]                      AP_AXIMM_22_AWREGION,
    input wire [3:0]                      AP_AXIMM_22_AWQOS,
    input wire                            AP_AXIMM_22_AWVALID,
    output  wire                            AP_AXIMM_22_AWREADY,
    input wire [M_AXIMM_22_DATA_WIDTH-1:0]   AP_AXIMM_22_WDATA,
    input wire [M_AXIMM_22_DATA_WIDTH/8-1:0] AP_AXIMM_22_WSTRB,
    input wire                            AP_AXIMM_22_WLAST,
    input wire                            AP_AXIMM_22_WVALID,
    output  wire                            AP_AXIMM_22_WREADY,
    output  wire [1:0]                      AP_AXIMM_22_BRESP,
    output  wire                            AP_AXIMM_22_BVALID,
    input wire                            AP_AXIMM_22_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_22_ARADDR,
    input wire [7:0]                      AP_AXIMM_22_ARLEN,
    input wire [2:0]                      AP_AXIMM_22_ARSIZE,
    input wire [1:0]                      AP_AXIMM_22_ARBURST,
    input wire [1:0]                      AP_AXIMM_22_ARLOCK,
    input wire [3:0]                      AP_AXIMM_22_ARCACHE,
    input wire [2:0]                      AP_AXIMM_22_ARPROT,
    input wire [3:0]                      AP_AXIMM_22_ARREGION,
    input wire [3:0]                      AP_AXIMM_22_ARQOS,
    input wire                            AP_AXIMM_22_ARVALID,
    output  wire                            AP_AXIMM_22_ARREADY,
    output  wire [M_AXIMM_22_DATA_WIDTH-1:0]   AP_AXIMM_22_RDATA,
    output  wire [1:0]                      AP_AXIMM_22_RRESP,
    output  wire                            AP_AXIMM_22_RLAST,
    output  wire                            AP_AXIMM_22_RVALID,
    input  wire                            AP_AXIMM_22_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_22_AWADDR,
    output wire [7:0]                      M_AXIMM_22_AWLEN,
    output wire [2:0]                      M_AXIMM_22_AWSIZE,
    output wire [1:0]                      M_AXIMM_22_AWBURST,
    output wire [1:0]                      M_AXIMM_22_AWLOCK,
    output wire [3:0]                      M_AXIMM_22_AWCACHE,
    output wire [2:0]                      M_AXIMM_22_AWPROT,
    output wire [3:0]                      M_AXIMM_22_AWREGION,
    output wire [3:0]                      M_AXIMM_22_AWQOS,
    output wire                            M_AXIMM_22_AWVALID,
    input  wire                            M_AXIMM_22_AWREADY,
    output wire [M_AXIMM_22_DATA_WIDTH-1:0]   M_AXIMM_22_WDATA,
    output wire [M_AXIMM_22_DATA_WIDTH/8-1:0] M_AXIMM_22_WSTRB,
    output wire                            M_AXIMM_22_WLAST,
    output wire                            M_AXIMM_22_WVALID,
    input  wire                            M_AXIMM_22_WREADY,
    input  wire [1:0]                      M_AXIMM_22_BRESP,
    input  wire                            M_AXIMM_22_BVALID,
    output wire                            M_AXIMM_22_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_22_ARADDR,
    output wire [7:0]                      M_AXIMM_22_ARLEN,
    output wire [2:0]                      M_AXIMM_22_ARSIZE,
    output wire [1:0]                      M_AXIMM_22_ARBURST,
    output wire [1:0]                      M_AXIMM_22_ARLOCK,
    output wire [3:0]                      M_AXIMM_22_ARCACHE,
    output wire [2:0]                      M_AXIMM_22_ARPROT,
    output wire [3:0]                      M_AXIMM_22_ARREGION,
    output wire [3:0]                      M_AXIMM_22_ARQOS,
    output wire                            M_AXIMM_22_ARVALID,
    input  wire                            M_AXIMM_22_ARREADY,
    input  wire [M_AXIMM_22_DATA_WIDTH-1:0]   M_AXIMM_22_RDATA,
    input  wire [1:0]                      M_AXIMM_22_RRESP,
    input  wire                            M_AXIMM_22_RLAST,
    input  wire                            M_AXIMM_22_RVALID,
    output wire                            M_AXIMM_22_RREADY,
    //AXI-MM pass-through interface 23
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_23_AWADDR,
    input wire [7:0]                      AP_AXIMM_23_AWLEN,
    input wire [2:0]                      AP_AXIMM_23_AWSIZE,
    input wire [1:0]                      AP_AXIMM_23_AWBURST,
    input wire [1:0]                      AP_AXIMM_23_AWLOCK,
    input wire [3:0]                      AP_AXIMM_23_AWCACHE,
    input wire [2:0]                      AP_AXIMM_23_AWPROT,
    input wire [3:0]                      AP_AXIMM_23_AWREGION,
    input wire [3:0]                      AP_AXIMM_23_AWQOS,
    input wire                            AP_AXIMM_23_AWVALID,
    output  wire                            AP_AXIMM_23_AWREADY,
    input wire [M_AXIMM_23_DATA_WIDTH-1:0]   AP_AXIMM_23_WDATA,
    input wire [M_AXIMM_23_DATA_WIDTH/8-1:0] AP_AXIMM_23_WSTRB,
    input wire                            AP_AXIMM_23_WLAST,
    input wire                            AP_AXIMM_23_WVALID,
    output  wire                            AP_AXIMM_23_WREADY,
    output  wire [1:0]                      AP_AXIMM_23_BRESP,
    output  wire                            AP_AXIMM_23_BVALID,
    input wire                            AP_AXIMM_23_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_23_ARADDR,
    input wire [7:0]                      AP_AXIMM_23_ARLEN,
    input wire [2:0]                      AP_AXIMM_23_ARSIZE,
    input wire [1:0]                      AP_AXIMM_23_ARBURST,
    input wire [1:0]                      AP_AXIMM_23_ARLOCK,
    input wire [3:0]                      AP_AXIMM_23_ARCACHE,
    input wire [2:0]                      AP_AXIMM_23_ARPROT,
    input wire [3:0]                      AP_AXIMM_23_ARREGION,
    input wire [3:0]                      AP_AXIMM_23_ARQOS,
    input wire                            AP_AXIMM_23_ARVALID,
    output  wire                            AP_AXIMM_23_ARREADY,
    output  wire [M_AXIMM_23_DATA_WIDTH-1:0]   AP_AXIMM_23_RDATA,
    output  wire [1:0]                      AP_AXIMM_23_RRESP,
    output  wire                            AP_AXIMM_23_RLAST,
    output  wire                            AP_AXIMM_23_RVALID,
    input  wire                            AP_AXIMM_23_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_23_AWADDR,
    output wire [7:0]                      M_AXIMM_23_AWLEN,
    output wire [2:0]                      M_AXIMM_23_AWSIZE,
    output wire [1:0]                      M_AXIMM_23_AWBURST,
    output wire [1:0]                      M_AXIMM_23_AWLOCK,
    output wire [3:0]                      M_AXIMM_23_AWCACHE,
    output wire [2:0]                      M_AXIMM_23_AWPROT,
    output wire [3:0]                      M_AXIMM_23_AWREGION,
    output wire [3:0]                      M_AXIMM_23_AWQOS,
    output wire                            M_AXIMM_23_AWVALID,
    input  wire                            M_AXIMM_23_AWREADY,
    output wire [M_AXIMM_23_DATA_WIDTH-1:0]   M_AXIMM_23_WDATA,
    output wire [M_AXIMM_23_DATA_WIDTH/8-1:0] M_AXIMM_23_WSTRB,
    output wire                            M_AXIMM_23_WLAST,
    output wire                            M_AXIMM_23_WVALID,
    input  wire                            M_AXIMM_23_WREADY,
    input  wire [1:0]                      M_AXIMM_23_BRESP,
    input  wire                            M_AXIMM_23_BVALID,
    output wire                            M_AXIMM_23_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_23_ARADDR,
    output wire [7:0]                      M_AXIMM_23_ARLEN,
    output wire [2:0]                      M_AXIMM_23_ARSIZE,
    output wire [1:0]                      M_AXIMM_23_ARBURST,
    output wire [1:0]                      M_AXIMM_23_ARLOCK,
    output wire [3:0]                      M_AXIMM_23_ARCACHE,
    output wire [2:0]                      M_AXIMM_23_ARPROT,
    output wire [3:0]                      M_AXIMM_23_ARREGION,
    output wire [3:0]                      M_AXIMM_23_ARQOS,
    output wire                            M_AXIMM_23_ARVALID,
    input  wire                            M_AXIMM_23_ARREADY,
    input  wire [M_AXIMM_23_DATA_WIDTH-1:0]   M_AXIMM_23_RDATA,
    input  wire [1:0]                      M_AXIMM_23_RRESP,
    input  wire                            M_AXIMM_23_RLAST,
    input  wire                            M_AXIMM_23_RVALID,
    output wire                            M_AXIMM_23_RREADY,
    //AXI-MM pass-through interface 24
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_24_AWADDR,
    input wire [7:0]                      AP_AXIMM_24_AWLEN,
    input wire [2:0]                      AP_AXIMM_24_AWSIZE,
    input wire [1:0]                      AP_AXIMM_24_AWBURST,
    input wire [1:0]                      AP_AXIMM_24_AWLOCK,
    input wire [3:0]                      AP_AXIMM_24_AWCACHE,
    input wire [2:0]                      AP_AXIMM_24_AWPROT,
    input wire [3:0]                      AP_AXIMM_24_AWREGION,
    input wire [3:0]                      AP_AXIMM_24_AWQOS,
    input wire                            AP_AXIMM_24_AWVALID,
    output  wire                            AP_AXIMM_24_AWREADY,
    input wire [M_AXIMM_24_DATA_WIDTH-1:0]   AP_AXIMM_24_WDATA,
    input wire [M_AXIMM_24_DATA_WIDTH/8-1:0] AP_AXIMM_24_WSTRB,
    input wire                            AP_AXIMM_24_WLAST,
    input wire                            AP_AXIMM_24_WVALID,
    output  wire                            AP_AXIMM_24_WREADY,
    output  wire [1:0]                      AP_AXIMM_24_BRESP,
    output  wire                            AP_AXIMM_24_BVALID,
    input wire                            AP_AXIMM_24_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_24_ARADDR,
    input wire [7:0]                      AP_AXIMM_24_ARLEN,
    input wire [2:0]                      AP_AXIMM_24_ARSIZE,
    input wire [1:0]                      AP_AXIMM_24_ARBURST,
    input wire [1:0]                      AP_AXIMM_24_ARLOCK,
    input wire [3:0]                      AP_AXIMM_24_ARCACHE,
    input wire [2:0]                      AP_AXIMM_24_ARPROT,
    input wire [3:0]                      AP_AXIMM_24_ARREGION,
    input wire [3:0]                      AP_AXIMM_24_ARQOS,
    input wire                            AP_AXIMM_24_ARVALID,
    output  wire                            AP_AXIMM_24_ARREADY,
    output  wire [M_AXIMM_24_DATA_WIDTH-1:0]   AP_AXIMM_24_RDATA,
    output  wire [1:0]                      AP_AXIMM_24_RRESP,
    output  wire                            AP_AXIMM_24_RLAST,
    output  wire                            AP_AXIMM_24_RVALID,
    input  wire                            AP_AXIMM_24_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_24_AWADDR,
    output wire [7:0]                      M_AXIMM_24_AWLEN,
    output wire [2:0]                      M_AXIMM_24_AWSIZE,
    output wire [1:0]                      M_AXIMM_24_AWBURST,
    output wire [1:0]                      M_AXIMM_24_AWLOCK,
    output wire [3:0]                      M_AXIMM_24_AWCACHE,
    output wire [2:0]                      M_AXIMM_24_AWPROT,
    output wire [3:0]                      M_AXIMM_24_AWREGION,
    output wire [3:0]                      M_AXIMM_24_AWQOS,
    output wire                            M_AXIMM_24_AWVALID,
    input  wire                            M_AXIMM_24_AWREADY,
    output wire [M_AXIMM_24_DATA_WIDTH-1:0]   M_AXIMM_24_WDATA,
    output wire [M_AXIMM_24_DATA_WIDTH/8-1:0] M_AXIMM_24_WSTRB,
    output wire                            M_AXIMM_24_WLAST,
    output wire                            M_AXIMM_24_WVALID,
    input  wire                            M_AXIMM_24_WREADY,
    input  wire [1:0]                      M_AXIMM_24_BRESP,
    input  wire                            M_AXIMM_24_BVALID,
    output wire                            M_AXIMM_24_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_24_ARADDR,
    output wire [7:0]                      M_AXIMM_24_ARLEN,
    output wire [2:0]                      M_AXIMM_24_ARSIZE,
    output wire [1:0]                      M_AXIMM_24_ARBURST,
    output wire [1:0]                      M_AXIMM_24_ARLOCK,
    output wire [3:0]                      M_AXIMM_24_ARCACHE,
    output wire [2:0]                      M_AXIMM_24_ARPROT,
    output wire [3:0]                      M_AXIMM_24_ARREGION,
    output wire [3:0]                      M_AXIMM_24_ARQOS,
    output wire                            M_AXIMM_24_ARVALID,
    input  wire                            M_AXIMM_24_ARREADY,
    input  wire [M_AXIMM_24_DATA_WIDTH-1:0]   M_AXIMM_24_RDATA,
    input  wire [1:0]                      M_AXIMM_24_RRESP,
    input  wire                            M_AXIMM_24_RLAST,
    input  wire                            M_AXIMM_24_RVALID,
    output wire                            M_AXIMM_24_RREADY,
    //AXI-MM pass-through interface 25
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_25_AWADDR,
    input wire [7:0]                      AP_AXIMM_25_AWLEN,
    input wire [2:0]                      AP_AXIMM_25_AWSIZE,
    input wire [1:0]                      AP_AXIMM_25_AWBURST,
    input wire [1:0]                      AP_AXIMM_25_AWLOCK,
    input wire [3:0]                      AP_AXIMM_25_AWCACHE,
    input wire [2:0]                      AP_AXIMM_25_AWPROT,
    input wire [3:0]                      AP_AXIMM_25_AWREGION,
    input wire [3:0]                      AP_AXIMM_25_AWQOS,
    input wire                            AP_AXIMM_25_AWVALID,
    output  wire                            AP_AXIMM_25_AWREADY,
    input wire [M_AXIMM_25_DATA_WIDTH-1:0]   AP_AXIMM_25_WDATA,
    input wire [M_AXIMM_25_DATA_WIDTH/8-1:0] AP_AXIMM_25_WSTRB,
    input wire                            AP_AXIMM_25_WLAST,
    input wire                            AP_AXIMM_25_WVALID,
    output  wire                            AP_AXIMM_25_WREADY,
    output  wire [1:0]                      AP_AXIMM_25_BRESP,
    output  wire                            AP_AXIMM_25_BVALID,
    input wire                            AP_AXIMM_25_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_25_ARADDR,
    input wire [7:0]                      AP_AXIMM_25_ARLEN,
    input wire [2:0]                      AP_AXIMM_25_ARSIZE,
    input wire [1:0]                      AP_AXIMM_25_ARBURST,
    input wire [1:0]                      AP_AXIMM_25_ARLOCK,
    input wire [3:0]                      AP_AXIMM_25_ARCACHE,
    input wire [2:0]                      AP_AXIMM_25_ARPROT,
    input wire [3:0]                      AP_AXIMM_25_ARREGION,
    input wire [3:0]                      AP_AXIMM_25_ARQOS,
    input wire                            AP_AXIMM_25_ARVALID,
    output  wire                            AP_AXIMM_25_ARREADY,
    output  wire [M_AXIMM_25_DATA_WIDTH-1:0]   AP_AXIMM_25_RDATA,
    output  wire [1:0]                      AP_AXIMM_25_RRESP,
    output  wire                            AP_AXIMM_25_RLAST,
    output  wire                            AP_AXIMM_25_RVALID,
    input  wire                            AP_AXIMM_25_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_25_AWADDR,
    output wire [7:0]                      M_AXIMM_25_AWLEN,
    output wire [2:0]                      M_AXIMM_25_AWSIZE,
    output wire [1:0]                      M_AXIMM_25_AWBURST,
    output wire [1:0]                      M_AXIMM_25_AWLOCK,
    output wire [3:0]                      M_AXIMM_25_AWCACHE,
    output wire [2:0]                      M_AXIMM_25_AWPROT,
    output wire [3:0]                      M_AXIMM_25_AWREGION,
    output wire [3:0]                      M_AXIMM_25_AWQOS,
    output wire                            M_AXIMM_25_AWVALID,
    input  wire                            M_AXIMM_25_AWREADY,
    output wire [M_AXIMM_25_DATA_WIDTH-1:0]   M_AXIMM_25_WDATA,
    output wire [M_AXIMM_25_DATA_WIDTH/8-1:0] M_AXIMM_25_WSTRB,
    output wire                            M_AXIMM_25_WLAST,
    output wire                            M_AXIMM_25_WVALID,
    input  wire                            M_AXIMM_25_WREADY,
    input  wire [1:0]                      M_AXIMM_25_BRESP,
    input  wire                            M_AXIMM_25_BVALID,
    output wire                            M_AXIMM_25_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_25_ARADDR,
    output wire [7:0]                      M_AXIMM_25_ARLEN,
    output wire [2:0]                      M_AXIMM_25_ARSIZE,
    output wire [1:0]                      M_AXIMM_25_ARBURST,
    output wire [1:0]                      M_AXIMM_25_ARLOCK,
    output wire [3:0]                      M_AXIMM_25_ARCACHE,
    output wire [2:0]                      M_AXIMM_25_ARPROT,
    output wire [3:0]                      M_AXIMM_25_ARREGION,
    output wire [3:0]                      M_AXIMM_25_ARQOS,
    output wire                            M_AXIMM_25_ARVALID,
    input  wire                            M_AXIMM_25_ARREADY,
    input  wire [M_AXIMM_25_DATA_WIDTH-1:0]   M_AXIMM_25_RDATA,
    input  wire [1:0]                      M_AXIMM_25_RRESP,
    input  wire                            M_AXIMM_25_RLAST,
    input  wire                            M_AXIMM_25_RVALID,
    output wire                            M_AXIMM_25_RREADY,
    //AXI-MM pass-through interface 26
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_26_AWADDR,
    input wire [7:0]                      AP_AXIMM_26_AWLEN,
    input wire [2:0]                      AP_AXIMM_26_AWSIZE,
    input wire [1:0]                      AP_AXIMM_26_AWBURST,
    input wire [1:0]                      AP_AXIMM_26_AWLOCK,
    input wire [3:0]                      AP_AXIMM_26_AWCACHE,
    input wire [2:0]                      AP_AXIMM_26_AWPROT,
    input wire [3:0]                      AP_AXIMM_26_AWREGION,
    input wire [3:0]                      AP_AXIMM_26_AWQOS,
    input wire                            AP_AXIMM_26_AWVALID,
    output  wire                            AP_AXIMM_26_AWREADY,
    input wire [M_AXIMM_26_DATA_WIDTH-1:0]   AP_AXIMM_26_WDATA,
    input wire [M_AXIMM_26_DATA_WIDTH/8-1:0] AP_AXIMM_26_WSTRB,
    input wire                            AP_AXIMM_26_WLAST,
    input wire                            AP_AXIMM_26_WVALID,
    output  wire                            AP_AXIMM_26_WREADY,
    output  wire [1:0]                      AP_AXIMM_26_BRESP,
    output  wire                            AP_AXIMM_26_BVALID,
    input wire                            AP_AXIMM_26_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_26_ARADDR,
    input wire [7:0]                      AP_AXIMM_26_ARLEN,
    input wire [2:0]                      AP_AXIMM_26_ARSIZE,
    input wire [1:0]                      AP_AXIMM_26_ARBURST,
    input wire [1:0]                      AP_AXIMM_26_ARLOCK,
    input wire [3:0]                      AP_AXIMM_26_ARCACHE,
    input wire [2:0]                      AP_AXIMM_26_ARPROT,
    input wire [3:0]                      AP_AXIMM_26_ARREGION,
    input wire [3:0]                      AP_AXIMM_26_ARQOS,
    input wire                            AP_AXIMM_26_ARVALID,
    output  wire                            AP_AXIMM_26_ARREADY,
    output  wire [M_AXIMM_26_DATA_WIDTH-1:0]   AP_AXIMM_26_RDATA,
    output  wire [1:0]                      AP_AXIMM_26_RRESP,
    output  wire                            AP_AXIMM_26_RLAST,
    output  wire                            AP_AXIMM_26_RVALID,
    input  wire                            AP_AXIMM_26_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_26_AWADDR,
    output wire [7:0]                      M_AXIMM_26_AWLEN,
    output wire [2:0]                      M_AXIMM_26_AWSIZE,
    output wire [1:0]                      M_AXIMM_26_AWBURST,
    output wire [1:0]                      M_AXIMM_26_AWLOCK,
    output wire [3:0]                      M_AXIMM_26_AWCACHE,
    output wire [2:0]                      M_AXIMM_26_AWPROT,
    output wire [3:0]                      M_AXIMM_26_AWREGION,
    output wire [3:0]                      M_AXIMM_26_AWQOS,
    output wire                            M_AXIMM_26_AWVALID,
    input  wire                            M_AXIMM_26_AWREADY,
    output wire [M_AXIMM_26_DATA_WIDTH-1:0]   M_AXIMM_26_WDATA,
    output wire [M_AXIMM_26_DATA_WIDTH/8-1:0] M_AXIMM_26_WSTRB,
    output wire                            M_AXIMM_26_WLAST,
    output wire                            M_AXIMM_26_WVALID,
    input  wire                            M_AXIMM_26_WREADY,
    input  wire [1:0]                      M_AXIMM_26_BRESP,
    input  wire                            M_AXIMM_26_BVALID,
    output wire                            M_AXIMM_26_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_26_ARADDR,
    output wire [7:0]                      M_AXIMM_26_ARLEN,
    output wire [2:0]                      M_AXIMM_26_ARSIZE,
    output wire [1:0]                      M_AXIMM_26_ARBURST,
    output wire [1:0]                      M_AXIMM_26_ARLOCK,
    output wire [3:0]                      M_AXIMM_26_ARCACHE,
    output wire [2:0]                      M_AXIMM_26_ARPROT,
    output wire [3:0]                      M_AXIMM_26_ARREGION,
    output wire [3:0]                      M_AXIMM_26_ARQOS,
    output wire                            M_AXIMM_26_ARVALID,
    input  wire                            M_AXIMM_26_ARREADY,
    input  wire [M_AXIMM_26_DATA_WIDTH-1:0]   M_AXIMM_26_RDATA,
    input  wire [1:0]                      M_AXIMM_26_RRESP,
    input  wire                            M_AXIMM_26_RLAST,
    input  wire                            M_AXIMM_26_RVALID,
    output wire                            M_AXIMM_26_RREADY,
    //AXI-MM pass-through interface 27
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_27_AWADDR,
    input wire [7:0]                      AP_AXIMM_27_AWLEN,
    input wire [2:0]                      AP_AXIMM_27_AWSIZE,
    input wire [1:0]                      AP_AXIMM_27_AWBURST,
    input wire [1:0]                      AP_AXIMM_27_AWLOCK,
    input wire [3:0]                      AP_AXIMM_27_AWCACHE,
    input wire [2:0]                      AP_AXIMM_27_AWPROT,
    input wire [3:0]                      AP_AXIMM_27_AWREGION,
    input wire [3:0]                      AP_AXIMM_27_AWQOS,
    input wire                            AP_AXIMM_27_AWVALID,
    output  wire                            AP_AXIMM_27_AWREADY,
    input wire [M_AXIMM_27_DATA_WIDTH-1:0]   AP_AXIMM_27_WDATA,
    input wire [M_AXIMM_27_DATA_WIDTH/8-1:0] AP_AXIMM_27_WSTRB,
    input wire                            AP_AXIMM_27_WLAST,
    input wire                            AP_AXIMM_27_WVALID,
    output  wire                            AP_AXIMM_27_WREADY,
    output  wire [1:0]                      AP_AXIMM_27_BRESP,
    output  wire                            AP_AXIMM_27_BVALID,
    input wire                            AP_AXIMM_27_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_27_ARADDR,
    input wire [7:0]                      AP_AXIMM_27_ARLEN,
    input wire [2:0]                      AP_AXIMM_27_ARSIZE,
    input wire [1:0]                      AP_AXIMM_27_ARBURST,
    input wire [1:0]                      AP_AXIMM_27_ARLOCK,
    input wire [3:0]                      AP_AXIMM_27_ARCACHE,
    input wire [2:0]                      AP_AXIMM_27_ARPROT,
    input wire [3:0]                      AP_AXIMM_27_ARREGION,
    input wire [3:0]                      AP_AXIMM_27_ARQOS,
    input wire                            AP_AXIMM_27_ARVALID,
    output  wire                            AP_AXIMM_27_ARREADY,
    output  wire [M_AXIMM_27_DATA_WIDTH-1:0]   AP_AXIMM_27_RDATA,
    output  wire [1:0]                      AP_AXIMM_27_RRESP,
    output  wire                            AP_AXIMM_27_RLAST,
    output  wire                            AP_AXIMM_27_RVALID,
    input  wire                            AP_AXIMM_27_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_27_AWADDR,
    output wire [7:0]                      M_AXIMM_27_AWLEN,
    output wire [2:0]                      M_AXIMM_27_AWSIZE,
    output wire [1:0]                      M_AXIMM_27_AWBURST,
    output wire [1:0]                      M_AXIMM_27_AWLOCK,
    output wire [3:0]                      M_AXIMM_27_AWCACHE,
    output wire [2:0]                      M_AXIMM_27_AWPROT,
    output wire [3:0]                      M_AXIMM_27_AWREGION,
    output wire [3:0]                      M_AXIMM_27_AWQOS,
    output wire                            M_AXIMM_27_AWVALID,
    input  wire                            M_AXIMM_27_AWREADY,
    output wire [M_AXIMM_27_DATA_WIDTH-1:0]   M_AXIMM_27_WDATA,
    output wire [M_AXIMM_27_DATA_WIDTH/8-1:0] M_AXIMM_27_WSTRB,
    output wire                            M_AXIMM_27_WLAST,
    output wire                            M_AXIMM_27_WVALID,
    input  wire                            M_AXIMM_27_WREADY,
    input  wire [1:0]                      M_AXIMM_27_BRESP,
    input  wire                            M_AXIMM_27_BVALID,
    output wire                            M_AXIMM_27_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_27_ARADDR,
    output wire [7:0]                      M_AXIMM_27_ARLEN,
    output wire [2:0]                      M_AXIMM_27_ARSIZE,
    output wire [1:0]                      M_AXIMM_27_ARBURST,
    output wire [1:0]                      M_AXIMM_27_ARLOCK,
    output wire [3:0]                      M_AXIMM_27_ARCACHE,
    output wire [2:0]                      M_AXIMM_27_ARPROT,
    output wire [3:0]                      M_AXIMM_27_ARREGION,
    output wire [3:0]                      M_AXIMM_27_ARQOS,
    output wire                            M_AXIMM_27_ARVALID,
    input  wire                            M_AXIMM_27_ARREADY,
    input  wire [M_AXIMM_27_DATA_WIDTH-1:0]   M_AXIMM_27_RDATA,
    input  wire [1:0]                      M_AXIMM_27_RRESP,
    input  wire                            M_AXIMM_27_RLAST,
    input  wire                            M_AXIMM_27_RVALID,
    output wire                            M_AXIMM_27_RREADY,
    //AXI-MM pass-through interface 28
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_28_AWADDR,
    input wire [7:0]                      AP_AXIMM_28_AWLEN,
    input wire [2:0]                      AP_AXIMM_28_AWSIZE,
    input wire [1:0]                      AP_AXIMM_28_AWBURST,
    input wire [1:0]                      AP_AXIMM_28_AWLOCK,
    input wire [3:0]                      AP_AXIMM_28_AWCACHE,
    input wire [2:0]                      AP_AXIMM_28_AWPROT,
    input wire [3:0]                      AP_AXIMM_28_AWREGION,
    input wire [3:0]                      AP_AXIMM_28_AWQOS,
    input wire                            AP_AXIMM_28_AWVALID,
    output  wire                            AP_AXIMM_28_AWREADY,
    input wire [M_AXIMM_28_DATA_WIDTH-1:0]   AP_AXIMM_28_WDATA,
    input wire [M_AXIMM_28_DATA_WIDTH/8-1:0] AP_AXIMM_28_WSTRB,
    input wire                            AP_AXIMM_28_WLAST,
    input wire                            AP_AXIMM_28_WVALID,
    output  wire                            AP_AXIMM_28_WREADY,
    output  wire [1:0]                      AP_AXIMM_28_BRESP,
    output  wire                            AP_AXIMM_28_BVALID,
    input wire                            AP_AXIMM_28_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_28_ARADDR,
    input wire [7:0]                      AP_AXIMM_28_ARLEN,
    input wire [2:0]                      AP_AXIMM_28_ARSIZE,
    input wire [1:0]                      AP_AXIMM_28_ARBURST,
    input wire [1:0]                      AP_AXIMM_28_ARLOCK,
    input wire [3:0]                      AP_AXIMM_28_ARCACHE,
    input wire [2:0]                      AP_AXIMM_28_ARPROT,
    input wire [3:0]                      AP_AXIMM_28_ARREGION,
    input wire [3:0]                      AP_AXIMM_28_ARQOS,
    input wire                            AP_AXIMM_28_ARVALID,
    output  wire                            AP_AXIMM_28_ARREADY,
    output  wire [M_AXIMM_28_DATA_WIDTH-1:0]   AP_AXIMM_28_RDATA,
    output  wire [1:0]                      AP_AXIMM_28_RRESP,
    output  wire                            AP_AXIMM_28_RLAST,
    output  wire                            AP_AXIMM_28_RVALID,
    input  wire                            AP_AXIMM_28_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_28_AWADDR,
    output wire [7:0]                      M_AXIMM_28_AWLEN,
    output wire [2:0]                      M_AXIMM_28_AWSIZE,
    output wire [1:0]                      M_AXIMM_28_AWBURST,
    output wire [1:0]                      M_AXIMM_28_AWLOCK,
    output wire [3:0]                      M_AXIMM_28_AWCACHE,
    output wire [2:0]                      M_AXIMM_28_AWPROT,
    output wire [3:0]                      M_AXIMM_28_AWREGION,
    output wire [3:0]                      M_AXIMM_28_AWQOS,
    output wire                            M_AXIMM_28_AWVALID,
    input  wire                            M_AXIMM_28_AWREADY,
    output wire [M_AXIMM_28_DATA_WIDTH-1:0]   M_AXIMM_28_WDATA,
    output wire [M_AXIMM_28_DATA_WIDTH/8-1:0] M_AXIMM_28_WSTRB,
    output wire                            M_AXIMM_28_WLAST,
    output wire                            M_AXIMM_28_WVALID,
    input  wire                            M_AXIMM_28_WREADY,
    input  wire [1:0]                      M_AXIMM_28_BRESP,
    input  wire                            M_AXIMM_28_BVALID,
    output wire                            M_AXIMM_28_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_28_ARADDR,
    output wire [7:0]                      M_AXIMM_28_ARLEN,
    output wire [2:0]                      M_AXIMM_28_ARSIZE,
    output wire [1:0]                      M_AXIMM_28_ARBURST,
    output wire [1:0]                      M_AXIMM_28_ARLOCK,
    output wire [3:0]                      M_AXIMM_28_ARCACHE,
    output wire [2:0]                      M_AXIMM_28_ARPROT,
    output wire [3:0]                      M_AXIMM_28_ARREGION,
    output wire [3:0]                      M_AXIMM_28_ARQOS,
    output wire                            M_AXIMM_28_ARVALID,
    input  wire                            M_AXIMM_28_ARREADY,
    input  wire [M_AXIMM_28_DATA_WIDTH-1:0]   M_AXIMM_28_RDATA,
    input  wire [1:0]                      M_AXIMM_28_RRESP,
    input  wire                            M_AXIMM_28_RLAST,
    input  wire                            M_AXIMM_28_RVALID,
    output wire                            M_AXIMM_28_RREADY,
    //AXI-MM pass-through interface 29
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_29_AWADDR,
    input wire [7:0]                      AP_AXIMM_29_AWLEN,
    input wire [2:0]                      AP_AXIMM_29_AWSIZE,
    input wire [1:0]                      AP_AXIMM_29_AWBURST,
    input wire [1:0]                      AP_AXIMM_29_AWLOCK,
    input wire [3:0]                      AP_AXIMM_29_AWCACHE,
    input wire [2:0]                      AP_AXIMM_29_AWPROT,
    input wire [3:0]                      AP_AXIMM_29_AWREGION,
    input wire [3:0]                      AP_AXIMM_29_AWQOS,
    input wire                            AP_AXIMM_29_AWVALID,
    output  wire                            AP_AXIMM_29_AWREADY,
    input wire [M_AXIMM_29_DATA_WIDTH-1:0]   AP_AXIMM_29_WDATA,
    input wire [M_AXIMM_29_DATA_WIDTH/8-1:0] AP_AXIMM_29_WSTRB,
    input wire                            AP_AXIMM_29_WLAST,
    input wire                            AP_AXIMM_29_WVALID,
    output  wire                            AP_AXIMM_29_WREADY,
    output  wire [1:0]                      AP_AXIMM_29_BRESP,
    output  wire                            AP_AXIMM_29_BVALID,
    input wire                            AP_AXIMM_29_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_29_ARADDR,
    input wire [7:0]                      AP_AXIMM_29_ARLEN,
    input wire [2:0]                      AP_AXIMM_29_ARSIZE,
    input wire [1:0]                      AP_AXIMM_29_ARBURST,
    input wire [1:0]                      AP_AXIMM_29_ARLOCK,
    input wire [3:0]                      AP_AXIMM_29_ARCACHE,
    input wire [2:0]                      AP_AXIMM_29_ARPROT,
    input wire [3:0]                      AP_AXIMM_29_ARREGION,
    input wire [3:0]                      AP_AXIMM_29_ARQOS,
    input wire                            AP_AXIMM_29_ARVALID,
    output  wire                            AP_AXIMM_29_ARREADY,
    output  wire [M_AXIMM_29_DATA_WIDTH-1:0]   AP_AXIMM_29_RDATA,
    output  wire [1:0]                      AP_AXIMM_29_RRESP,
    output  wire                            AP_AXIMM_29_RLAST,
    output  wire                            AP_AXIMM_29_RVALID,
    input  wire                            AP_AXIMM_29_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_29_AWADDR,
    output wire [7:0]                      M_AXIMM_29_AWLEN,
    output wire [2:0]                      M_AXIMM_29_AWSIZE,
    output wire [1:0]                      M_AXIMM_29_AWBURST,
    output wire [1:0]                      M_AXIMM_29_AWLOCK,
    output wire [3:0]                      M_AXIMM_29_AWCACHE,
    output wire [2:0]                      M_AXIMM_29_AWPROT,
    output wire [3:0]                      M_AXIMM_29_AWREGION,
    output wire [3:0]                      M_AXIMM_29_AWQOS,
    output wire                            M_AXIMM_29_AWVALID,
    input  wire                            M_AXIMM_29_AWREADY,
    output wire [M_AXIMM_29_DATA_WIDTH-1:0]   M_AXIMM_29_WDATA,
    output wire [M_AXIMM_29_DATA_WIDTH/8-1:0] M_AXIMM_29_WSTRB,
    output wire                            M_AXIMM_29_WLAST,
    output wire                            M_AXIMM_29_WVALID,
    input  wire                            M_AXIMM_29_WREADY,
    input  wire [1:0]                      M_AXIMM_29_BRESP,
    input  wire                            M_AXIMM_29_BVALID,
    output wire                            M_AXIMM_29_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_29_ARADDR,
    output wire [7:0]                      M_AXIMM_29_ARLEN,
    output wire [2:0]                      M_AXIMM_29_ARSIZE,
    output wire [1:0]                      M_AXIMM_29_ARBURST,
    output wire [1:0]                      M_AXIMM_29_ARLOCK,
    output wire [3:0]                      M_AXIMM_29_ARCACHE,
    output wire [2:0]                      M_AXIMM_29_ARPROT,
    output wire [3:0]                      M_AXIMM_29_ARREGION,
    output wire [3:0]                      M_AXIMM_29_ARQOS,
    output wire                            M_AXIMM_29_ARVALID,
    input  wire                            M_AXIMM_29_ARREADY,
    input  wire [M_AXIMM_29_DATA_WIDTH-1:0]   M_AXIMM_29_RDATA,
    input  wire [1:0]                      M_AXIMM_29_RRESP,
    input  wire                            M_AXIMM_29_RLAST,
    input  wire                            M_AXIMM_29_RVALID,
    output wire                            M_AXIMM_29_RREADY,
    //AXI-MM pass-through interface 30
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_30_AWADDR,
    input wire [7:0]                      AP_AXIMM_30_AWLEN,
    input wire [2:0]                      AP_AXIMM_30_AWSIZE,
    input wire [1:0]                      AP_AXIMM_30_AWBURST,
    input wire [1:0]                      AP_AXIMM_30_AWLOCK,
    input wire [3:0]                      AP_AXIMM_30_AWCACHE,
    input wire [2:0]                      AP_AXIMM_30_AWPROT,
    input wire [3:0]                      AP_AXIMM_30_AWREGION,
    input wire [3:0]                      AP_AXIMM_30_AWQOS,
    input wire                            AP_AXIMM_30_AWVALID,
    output  wire                            AP_AXIMM_30_AWREADY,
    input wire [M_AXIMM_30_DATA_WIDTH-1:0]   AP_AXIMM_30_WDATA,
    input wire [M_AXIMM_30_DATA_WIDTH/8-1:0] AP_AXIMM_30_WSTRB,
    input wire                            AP_AXIMM_30_WLAST,
    input wire                            AP_AXIMM_30_WVALID,
    output  wire                            AP_AXIMM_30_WREADY,
    output  wire [1:0]                      AP_AXIMM_30_BRESP,
    output  wire                            AP_AXIMM_30_BVALID,
    input wire                            AP_AXIMM_30_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_30_ARADDR,
    input wire [7:0]                      AP_AXIMM_30_ARLEN,
    input wire [2:0]                      AP_AXIMM_30_ARSIZE,
    input wire [1:0]                      AP_AXIMM_30_ARBURST,
    input wire [1:0]                      AP_AXIMM_30_ARLOCK,
    input wire [3:0]                      AP_AXIMM_30_ARCACHE,
    input wire [2:0]                      AP_AXIMM_30_ARPROT,
    input wire [3:0]                      AP_AXIMM_30_ARREGION,
    input wire [3:0]                      AP_AXIMM_30_ARQOS,
    input wire                            AP_AXIMM_30_ARVALID,
    output  wire                            AP_AXIMM_30_ARREADY,
    output  wire [M_AXIMM_30_DATA_WIDTH-1:0]   AP_AXIMM_30_RDATA,
    output  wire [1:0]                      AP_AXIMM_30_RRESP,
    output  wire                            AP_AXIMM_30_RLAST,
    output  wire                            AP_AXIMM_30_RVALID,
    input  wire                            AP_AXIMM_30_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_30_AWADDR,
    output wire [7:0]                      M_AXIMM_30_AWLEN,
    output wire [2:0]                      M_AXIMM_30_AWSIZE,
    output wire [1:0]                      M_AXIMM_30_AWBURST,
    output wire [1:0]                      M_AXIMM_30_AWLOCK,
    output wire [3:0]                      M_AXIMM_30_AWCACHE,
    output wire [2:0]                      M_AXIMM_30_AWPROT,
    output wire [3:0]                      M_AXIMM_30_AWREGION,
    output wire [3:0]                      M_AXIMM_30_AWQOS,
    output wire                            M_AXIMM_30_AWVALID,
    input  wire                            M_AXIMM_30_AWREADY,
    output wire [M_AXIMM_30_DATA_WIDTH-1:0]   M_AXIMM_30_WDATA,
    output wire [M_AXIMM_30_DATA_WIDTH/8-1:0] M_AXIMM_30_WSTRB,
    output wire                            M_AXIMM_30_WLAST,
    output wire                            M_AXIMM_30_WVALID,
    input  wire                            M_AXIMM_30_WREADY,
    input  wire [1:0]                      M_AXIMM_30_BRESP,
    input  wire                            M_AXIMM_30_BVALID,
    output wire                            M_AXIMM_30_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_30_ARADDR,
    output wire [7:0]                      M_AXIMM_30_ARLEN,
    output wire [2:0]                      M_AXIMM_30_ARSIZE,
    output wire [1:0]                      M_AXIMM_30_ARBURST,
    output wire [1:0]                      M_AXIMM_30_ARLOCK,
    output wire [3:0]                      M_AXIMM_30_ARCACHE,
    output wire [2:0]                      M_AXIMM_30_ARPROT,
    output wire [3:0]                      M_AXIMM_30_ARREGION,
    output wire [3:0]                      M_AXIMM_30_ARQOS,
    output wire                            M_AXIMM_30_ARVALID,
    input  wire                            M_AXIMM_30_ARREADY,
    input  wire [M_AXIMM_30_DATA_WIDTH-1:0]   M_AXIMM_30_RDATA,
    input  wire [1:0]                      M_AXIMM_30_RRESP,
    input  wire                            M_AXIMM_30_RLAST,
    input  wire                            M_AXIMM_30_RVALID,
    output wire                            M_AXIMM_30_RREADY,
    //AXI-MM pass-through interface 31
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_31_AWADDR,
    input wire [7:0]                      AP_AXIMM_31_AWLEN,
    input wire [2:0]                      AP_AXIMM_31_AWSIZE,
    input wire [1:0]                      AP_AXIMM_31_AWBURST,
    input wire [1:0]                      AP_AXIMM_31_AWLOCK,
    input wire [3:0]                      AP_AXIMM_31_AWCACHE,
    input wire [2:0]                      AP_AXIMM_31_AWPROT,
    input wire [3:0]                      AP_AXIMM_31_AWREGION,
    input wire [3:0]                      AP_AXIMM_31_AWQOS,
    input wire                            AP_AXIMM_31_AWVALID,
    output  wire                            AP_AXIMM_31_AWREADY,
    input wire [M_AXIMM_31_DATA_WIDTH-1:0]   AP_AXIMM_31_WDATA,
    input wire [M_AXIMM_31_DATA_WIDTH/8-1:0] AP_AXIMM_31_WSTRB,
    input wire                            AP_AXIMM_31_WLAST,
    input wire                            AP_AXIMM_31_WVALID,
    output  wire                            AP_AXIMM_31_WREADY,
    output  wire [1:0]                      AP_AXIMM_31_BRESP,
    output  wire                            AP_AXIMM_31_BVALID,
    input wire                            AP_AXIMM_31_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_31_ARADDR,
    input wire [7:0]                      AP_AXIMM_31_ARLEN,
    input wire [2:0]                      AP_AXIMM_31_ARSIZE,
    input wire [1:0]                      AP_AXIMM_31_ARBURST,
    input wire [1:0]                      AP_AXIMM_31_ARLOCK,
    input wire [3:0]                      AP_AXIMM_31_ARCACHE,
    input wire [2:0]                      AP_AXIMM_31_ARPROT,
    input wire [3:0]                      AP_AXIMM_31_ARREGION,
    input wire [3:0]                      AP_AXIMM_31_ARQOS,
    input wire                            AP_AXIMM_31_ARVALID,
    output  wire                            AP_AXIMM_31_ARREADY,
    output  wire [M_AXIMM_31_DATA_WIDTH-1:0]   AP_AXIMM_31_RDATA,
    output  wire [1:0]                      AP_AXIMM_31_RRESP,
    output  wire                            AP_AXIMM_31_RLAST,
    output  wire                            AP_AXIMM_31_RVALID,
    input  wire                            AP_AXIMM_31_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_31_AWADDR,
    output wire [7:0]                      M_AXIMM_31_AWLEN,
    output wire [2:0]                      M_AXIMM_31_AWSIZE,
    output wire [1:0]                      M_AXIMM_31_AWBURST,
    output wire [1:0]                      M_AXIMM_31_AWLOCK,
    output wire [3:0]                      M_AXIMM_31_AWCACHE,
    output wire [2:0]                      M_AXIMM_31_AWPROT,
    output wire [3:0]                      M_AXIMM_31_AWREGION,
    output wire [3:0]                      M_AXIMM_31_AWQOS,
    output wire                            M_AXIMM_31_AWVALID,
    input  wire                            M_AXIMM_31_AWREADY,
    output wire [M_AXIMM_31_DATA_WIDTH-1:0]   M_AXIMM_31_WDATA,
    output wire [M_AXIMM_31_DATA_WIDTH/8-1:0] M_AXIMM_31_WSTRB,
    output wire                            M_AXIMM_31_WLAST,
    output wire                            M_AXIMM_31_WVALID,
    input  wire                            M_AXIMM_31_WREADY,
    input  wire [1:0]                      M_AXIMM_31_BRESP,
    input  wire                            M_AXIMM_31_BVALID,
    output wire                            M_AXIMM_31_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_31_ARADDR,
    output wire [7:0]                      M_AXIMM_31_ARLEN,
    output wire [2:0]                      M_AXIMM_31_ARSIZE,
    output wire [1:0]                      M_AXIMM_31_ARBURST,
    output wire [1:0]                      M_AXIMM_31_ARLOCK,
    output wire [3:0]                      M_AXIMM_31_ARCACHE,
    output wire [2:0]                      M_AXIMM_31_ARPROT,
    output wire [3:0]                      M_AXIMM_31_ARREGION,
    output wire [3:0]                      M_AXIMM_31_ARQOS,
    output wire                            M_AXIMM_31_ARVALID,
    input  wire                            M_AXIMM_31_ARREADY,
    input  wire [M_AXIMM_31_DATA_WIDTH-1:0]   M_AXIMM_31_RDATA,
    input  wire [1:0]                      M_AXIMM_31_RRESP,
    input  wire                            M_AXIMM_31_RLAST,
    input  wire                            M_AXIMM_31_RVALID,
    output wire                            M_AXIMM_31_RREADY,
    //AXI-MM pass-through interface 32
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_32_AWADDR,
    input wire [7:0]                      AP_AXIMM_32_AWLEN,
    input wire [2:0]                      AP_AXIMM_32_AWSIZE,
    input wire [1:0]                      AP_AXIMM_32_AWBURST,
    input wire [1:0]                      AP_AXIMM_32_AWLOCK,
    input wire [3:0]                      AP_AXIMM_32_AWCACHE,
    input wire [2:0]                      AP_AXIMM_32_AWPROT,
    input wire [3:0]                      AP_AXIMM_32_AWREGION,
    input wire [3:0]                      AP_AXIMM_32_AWQOS,
    input wire                            AP_AXIMM_32_AWVALID,
    output  wire                            AP_AXIMM_32_AWREADY,
    input wire [M_AXIMM_32_DATA_WIDTH-1:0]   AP_AXIMM_32_WDATA,
    input wire [M_AXIMM_32_DATA_WIDTH/8-1:0] AP_AXIMM_32_WSTRB,
    input wire                            AP_AXIMM_32_WLAST,
    input wire                            AP_AXIMM_32_WVALID,
    output  wire                            AP_AXIMM_32_WREADY,
    output  wire [1:0]                      AP_AXIMM_32_BRESP,
    output  wire                            AP_AXIMM_32_BVALID,
    input wire                            AP_AXIMM_32_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_32_ARADDR,
    input wire [7:0]                      AP_AXIMM_32_ARLEN,
    input wire [2:0]                      AP_AXIMM_32_ARSIZE,
    input wire [1:0]                      AP_AXIMM_32_ARBURST,
    input wire [1:0]                      AP_AXIMM_32_ARLOCK,
    input wire [3:0]                      AP_AXIMM_32_ARCACHE,
    input wire [2:0]                      AP_AXIMM_32_ARPROT,
    input wire [3:0]                      AP_AXIMM_32_ARREGION,
    input wire [3:0]                      AP_AXIMM_32_ARQOS,
    input wire                            AP_AXIMM_32_ARVALID,
    output  wire                            AP_AXIMM_32_ARREADY,
    output  wire [M_AXIMM_32_DATA_WIDTH-1:0]   AP_AXIMM_32_RDATA,
    output  wire [1:0]                      AP_AXIMM_32_RRESP,
    output  wire                            AP_AXIMM_32_RLAST,
    output  wire                            AP_AXIMM_32_RVALID,
    input  wire                            AP_AXIMM_32_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_32_AWADDR,
    output wire [7:0]                      M_AXIMM_32_AWLEN,
    output wire [2:0]                      M_AXIMM_32_AWSIZE,
    output wire [1:0]                      M_AXIMM_32_AWBURST,
    output wire [1:0]                      M_AXIMM_32_AWLOCK,
    output wire [3:0]                      M_AXIMM_32_AWCACHE,
    output wire [2:0]                      M_AXIMM_32_AWPROT,
    output wire [3:0]                      M_AXIMM_32_AWREGION,
    output wire [3:0]                      M_AXIMM_32_AWQOS,
    output wire                            M_AXIMM_32_AWVALID,
    input  wire                            M_AXIMM_32_AWREADY,
    output wire [M_AXIMM_32_DATA_WIDTH-1:0]   M_AXIMM_32_WDATA,
    output wire [M_AXIMM_32_DATA_WIDTH/8-1:0] M_AXIMM_32_WSTRB,
    output wire                            M_AXIMM_32_WLAST,
    output wire                            M_AXIMM_32_WVALID,
    input  wire                            M_AXIMM_32_WREADY,
    input  wire [1:0]                      M_AXIMM_32_BRESP,
    input  wire                            M_AXIMM_32_BVALID,
    output wire                            M_AXIMM_32_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_32_ARADDR,
    output wire [7:0]                      M_AXIMM_32_ARLEN,
    output wire [2:0]                      M_AXIMM_32_ARSIZE,
    output wire [1:0]                      M_AXIMM_32_ARBURST,
    output wire [1:0]                      M_AXIMM_32_ARLOCK,
    output wire [3:0]                      M_AXIMM_32_ARCACHE,
    output wire [2:0]                      M_AXIMM_32_ARPROT,
    output wire [3:0]                      M_AXIMM_32_ARREGION,
    output wire [3:0]                      M_AXIMM_32_ARQOS,
    output wire                            M_AXIMM_32_ARVALID,
    input  wire                            M_AXIMM_32_ARREADY,
    input  wire [M_AXIMM_32_DATA_WIDTH-1:0]   M_AXIMM_32_RDATA,
    input  wire [1:0]                      M_AXIMM_32_RRESP,
    input  wire                            M_AXIMM_32_RLAST,
    input  wire                            M_AXIMM_32_RVALID,
    output wire                            M_AXIMM_32_RREADY,
    //AXI-MM pass-through interface 33
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_33_AWADDR,
    input wire [7:0]                      AP_AXIMM_33_AWLEN,
    input wire [2:0]                      AP_AXIMM_33_AWSIZE,
    input wire [1:0]                      AP_AXIMM_33_AWBURST,
    input wire [1:0]                      AP_AXIMM_33_AWLOCK,
    input wire [3:0]                      AP_AXIMM_33_AWCACHE,
    input wire [2:0]                      AP_AXIMM_33_AWPROT,
    input wire [3:0]                      AP_AXIMM_33_AWREGION,
    input wire [3:0]                      AP_AXIMM_33_AWQOS,
    input wire                            AP_AXIMM_33_AWVALID,
    output  wire                            AP_AXIMM_33_AWREADY,
    input wire [M_AXIMM_33_DATA_WIDTH-1:0]   AP_AXIMM_33_WDATA,
    input wire [M_AXIMM_33_DATA_WIDTH/8-1:0] AP_AXIMM_33_WSTRB,
    input wire                            AP_AXIMM_33_WLAST,
    input wire                            AP_AXIMM_33_WVALID,
    output  wire                            AP_AXIMM_33_WREADY,
    output  wire [1:0]                      AP_AXIMM_33_BRESP,
    output  wire                            AP_AXIMM_33_BVALID,
    input wire                            AP_AXIMM_33_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_33_ARADDR,
    input wire [7:0]                      AP_AXIMM_33_ARLEN,
    input wire [2:0]                      AP_AXIMM_33_ARSIZE,
    input wire [1:0]                      AP_AXIMM_33_ARBURST,
    input wire [1:0]                      AP_AXIMM_33_ARLOCK,
    input wire [3:0]                      AP_AXIMM_33_ARCACHE,
    input wire [2:0]                      AP_AXIMM_33_ARPROT,
    input wire [3:0]                      AP_AXIMM_33_ARREGION,
    input wire [3:0]                      AP_AXIMM_33_ARQOS,
    input wire                            AP_AXIMM_33_ARVALID,
    output  wire                            AP_AXIMM_33_ARREADY,
    output  wire [M_AXIMM_33_DATA_WIDTH-1:0]   AP_AXIMM_33_RDATA,
    output  wire [1:0]                      AP_AXIMM_33_RRESP,
    output  wire                            AP_AXIMM_33_RLAST,
    output  wire                            AP_AXIMM_33_RVALID,
    input  wire                            AP_AXIMM_33_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_33_AWADDR,
    output wire [7:0]                      M_AXIMM_33_AWLEN,
    output wire [2:0]                      M_AXIMM_33_AWSIZE,
    output wire [1:0]                      M_AXIMM_33_AWBURST,
    output wire [1:0]                      M_AXIMM_33_AWLOCK,
    output wire [3:0]                      M_AXIMM_33_AWCACHE,
    output wire [2:0]                      M_AXIMM_33_AWPROT,
    output wire [3:0]                      M_AXIMM_33_AWREGION,
    output wire [3:0]                      M_AXIMM_33_AWQOS,
    output wire                            M_AXIMM_33_AWVALID,
    input  wire                            M_AXIMM_33_AWREADY,
    output wire [M_AXIMM_33_DATA_WIDTH-1:0]   M_AXIMM_33_WDATA,
    output wire [M_AXIMM_33_DATA_WIDTH/8-1:0] M_AXIMM_33_WSTRB,
    output wire                            M_AXIMM_33_WLAST,
    output wire                            M_AXIMM_33_WVALID,
    input  wire                            M_AXIMM_33_WREADY,
    input  wire [1:0]                      M_AXIMM_33_BRESP,
    input  wire                            M_AXIMM_33_BVALID,
    output wire                            M_AXIMM_33_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_33_ARADDR,
    output wire [7:0]                      M_AXIMM_33_ARLEN,
    output wire [2:0]                      M_AXIMM_33_ARSIZE,
    output wire [1:0]                      M_AXIMM_33_ARBURST,
    output wire [1:0]                      M_AXIMM_33_ARLOCK,
    output wire [3:0]                      M_AXIMM_33_ARCACHE,
    output wire [2:0]                      M_AXIMM_33_ARPROT,
    output wire [3:0]                      M_AXIMM_33_ARREGION,
    output wire [3:0]                      M_AXIMM_33_ARQOS,
    output wire                            M_AXIMM_33_ARVALID,
    input  wire                            M_AXIMM_33_ARREADY,
    input  wire [M_AXIMM_33_DATA_WIDTH-1:0]   M_AXIMM_33_RDATA,
    input  wire [1:0]                      M_AXIMM_33_RRESP,
    input  wire                            M_AXIMM_33_RLAST,
    input  wire                            M_AXIMM_33_RVALID,
    output wire                            M_AXIMM_33_RREADY,
    //AXI-MM pass-through interface 34
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_34_AWADDR,
    input wire [7:0]                      AP_AXIMM_34_AWLEN,
    input wire [2:0]                      AP_AXIMM_34_AWSIZE,
    input wire [1:0]                      AP_AXIMM_34_AWBURST,
    input wire [1:0]                      AP_AXIMM_34_AWLOCK,
    input wire [3:0]                      AP_AXIMM_34_AWCACHE,
    input wire [2:0]                      AP_AXIMM_34_AWPROT,
    input wire [3:0]                      AP_AXIMM_34_AWREGION,
    input wire [3:0]                      AP_AXIMM_34_AWQOS,
    input wire                            AP_AXIMM_34_AWVALID,
    output  wire                            AP_AXIMM_34_AWREADY,
    input wire [M_AXIMM_34_DATA_WIDTH-1:0]   AP_AXIMM_34_WDATA,
    input wire [M_AXIMM_34_DATA_WIDTH/8-1:0] AP_AXIMM_34_WSTRB,
    input wire                            AP_AXIMM_34_WLAST,
    input wire                            AP_AXIMM_34_WVALID,
    output  wire                            AP_AXIMM_34_WREADY,
    output  wire [1:0]                      AP_AXIMM_34_BRESP,
    output  wire                            AP_AXIMM_34_BVALID,
    input wire                            AP_AXIMM_34_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_34_ARADDR,
    input wire [7:0]                      AP_AXIMM_34_ARLEN,
    input wire [2:0]                      AP_AXIMM_34_ARSIZE,
    input wire [1:0]                      AP_AXIMM_34_ARBURST,
    input wire [1:0]                      AP_AXIMM_34_ARLOCK,
    input wire [3:0]                      AP_AXIMM_34_ARCACHE,
    input wire [2:0]                      AP_AXIMM_34_ARPROT,
    input wire [3:0]                      AP_AXIMM_34_ARREGION,
    input wire [3:0]                      AP_AXIMM_34_ARQOS,
    input wire                            AP_AXIMM_34_ARVALID,
    output  wire                            AP_AXIMM_34_ARREADY,
    output  wire [M_AXIMM_34_DATA_WIDTH-1:0]   AP_AXIMM_34_RDATA,
    output  wire [1:0]                      AP_AXIMM_34_RRESP,
    output  wire                            AP_AXIMM_34_RLAST,
    output  wire                            AP_AXIMM_34_RVALID,
    input  wire                            AP_AXIMM_34_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_34_AWADDR,
    output wire [7:0]                      M_AXIMM_34_AWLEN,
    output wire [2:0]                      M_AXIMM_34_AWSIZE,
    output wire [1:0]                      M_AXIMM_34_AWBURST,
    output wire [1:0]                      M_AXIMM_34_AWLOCK,
    output wire [3:0]                      M_AXIMM_34_AWCACHE,
    output wire [2:0]                      M_AXIMM_34_AWPROT,
    output wire [3:0]                      M_AXIMM_34_AWREGION,
    output wire [3:0]                      M_AXIMM_34_AWQOS,
    output wire                            M_AXIMM_34_AWVALID,
    input  wire                            M_AXIMM_34_AWREADY,
    output wire [M_AXIMM_34_DATA_WIDTH-1:0]   M_AXIMM_34_WDATA,
    output wire [M_AXIMM_34_DATA_WIDTH/8-1:0] M_AXIMM_34_WSTRB,
    output wire                            M_AXIMM_34_WLAST,
    output wire                            M_AXIMM_34_WVALID,
    input  wire                            M_AXIMM_34_WREADY,
    input  wire [1:0]                      M_AXIMM_34_BRESP,
    input  wire                            M_AXIMM_34_BVALID,
    output wire                            M_AXIMM_34_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_34_ARADDR,
    output wire [7:0]                      M_AXIMM_34_ARLEN,
    output wire [2:0]                      M_AXIMM_34_ARSIZE,
    output wire [1:0]                      M_AXIMM_34_ARBURST,
    output wire [1:0]                      M_AXIMM_34_ARLOCK,
    output wire [3:0]                      M_AXIMM_34_ARCACHE,
    output wire [2:0]                      M_AXIMM_34_ARPROT,
    output wire [3:0]                      M_AXIMM_34_ARREGION,
    output wire [3:0]                      M_AXIMM_34_ARQOS,
    output wire                            M_AXIMM_34_ARVALID,
    input  wire                            M_AXIMM_34_ARREADY,
    input  wire [M_AXIMM_34_DATA_WIDTH-1:0]   M_AXIMM_34_RDATA,
    input  wire [1:0]                      M_AXIMM_34_RRESP,
    input  wire                            M_AXIMM_34_RLAST,
    input  wire                            M_AXIMM_34_RVALID,
    output wire                            M_AXIMM_34_RREADY,
    //AXI-MM pass-through interface 35
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_35_AWADDR,
    input wire [7:0]                      AP_AXIMM_35_AWLEN,
    input wire [2:0]                      AP_AXIMM_35_AWSIZE,
    input wire [1:0]                      AP_AXIMM_35_AWBURST,
    input wire [1:0]                      AP_AXIMM_35_AWLOCK,
    input wire [3:0]                      AP_AXIMM_35_AWCACHE,
    input wire [2:0]                      AP_AXIMM_35_AWPROT,
    input wire [3:0]                      AP_AXIMM_35_AWREGION,
    input wire [3:0]                      AP_AXIMM_35_AWQOS,
    input wire                            AP_AXIMM_35_AWVALID,
    output  wire                            AP_AXIMM_35_AWREADY,
    input wire [M_AXIMM_35_DATA_WIDTH-1:0]   AP_AXIMM_35_WDATA,
    input wire [M_AXIMM_35_DATA_WIDTH/8-1:0] AP_AXIMM_35_WSTRB,
    input wire                            AP_AXIMM_35_WLAST,
    input wire                            AP_AXIMM_35_WVALID,
    output  wire                            AP_AXIMM_35_WREADY,
    output  wire [1:0]                      AP_AXIMM_35_BRESP,
    output  wire                            AP_AXIMM_35_BVALID,
    input wire                            AP_AXIMM_35_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_35_ARADDR,
    input wire [7:0]                      AP_AXIMM_35_ARLEN,
    input wire [2:0]                      AP_AXIMM_35_ARSIZE,
    input wire [1:0]                      AP_AXIMM_35_ARBURST,
    input wire [1:0]                      AP_AXIMM_35_ARLOCK,
    input wire [3:0]                      AP_AXIMM_35_ARCACHE,
    input wire [2:0]                      AP_AXIMM_35_ARPROT,
    input wire [3:0]                      AP_AXIMM_35_ARREGION,
    input wire [3:0]                      AP_AXIMM_35_ARQOS,
    input wire                            AP_AXIMM_35_ARVALID,
    output  wire                            AP_AXIMM_35_ARREADY,
    output  wire [M_AXIMM_35_DATA_WIDTH-1:0]   AP_AXIMM_35_RDATA,
    output  wire [1:0]                      AP_AXIMM_35_RRESP,
    output  wire                            AP_AXIMM_35_RLAST,
    output  wire                            AP_AXIMM_35_RVALID,
    input  wire                            AP_AXIMM_35_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_35_AWADDR,
    output wire [7:0]                      M_AXIMM_35_AWLEN,
    output wire [2:0]                      M_AXIMM_35_AWSIZE,
    output wire [1:0]                      M_AXIMM_35_AWBURST,
    output wire [1:0]                      M_AXIMM_35_AWLOCK,
    output wire [3:0]                      M_AXIMM_35_AWCACHE,
    output wire [2:0]                      M_AXIMM_35_AWPROT,
    output wire [3:0]                      M_AXIMM_35_AWREGION,
    output wire [3:0]                      M_AXIMM_35_AWQOS,
    output wire                            M_AXIMM_35_AWVALID,
    input  wire                            M_AXIMM_35_AWREADY,
    output wire [M_AXIMM_35_DATA_WIDTH-1:0]   M_AXIMM_35_WDATA,
    output wire [M_AXIMM_35_DATA_WIDTH/8-1:0] M_AXIMM_35_WSTRB,
    output wire                            M_AXIMM_35_WLAST,
    output wire                            M_AXIMM_35_WVALID,
    input  wire                            M_AXIMM_35_WREADY,
    input  wire [1:0]                      M_AXIMM_35_BRESP,
    input  wire                            M_AXIMM_35_BVALID,
    output wire                            M_AXIMM_35_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_35_ARADDR,
    output wire [7:0]                      M_AXIMM_35_ARLEN,
    output wire [2:0]                      M_AXIMM_35_ARSIZE,
    output wire [1:0]                      M_AXIMM_35_ARBURST,
    output wire [1:0]                      M_AXIMM_35_ARLOCK,
    output wire [3:0]                      M_AXIMM_35_ARCACHE,
    output wire [2:0]                      M_AXIMM_35_ARPROT,
    output wire [3:0]                      M_AXIMM_35_ARREGION,
    output wire [3:0]                      M_AXIMM_35_ARQOS,
    output wire                            M_AXIMM_35_ARVALID,
    input  wire                            M_AXIMM_35_ARREADY,
    input  wire [M_AXIMM_35_DATA_WIDTH-1:0]   M_AXIMM_35_RDATA,
    input  wire [1:0]                      M_AXIMM_35_RRESP,
    input  wire                            M_AXIMM_35_RLAST,
    input  wire                            M_AXIMM_35_RVALID,
    output wire                            M_AXIMM_35_RREADY,
    //AXI-MM pass-through interface 36
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_36_AWADDR,
    input wire [7:0]                      AP_AXIMM_36_AWLEN,
    input wire [2:0]                      AP_AXIMM_36_AWSIZE,
    input wire [1:0]                      AP_AXIMM_36_AWBURST,
    input wire [1:0]                      AP_AXIMM_36_AWLOCK,
    input wire [3:0]                      AP_AXIMM_36_AWCACHE,
    input wire [2:0]                      AP_AXIMM_36_AWPROT,
    input wire [3:0]                      AP_AXIMM_36_AWREGION,
    input wire [3:0]                      AP_AXIMM_36_AWQOS,
    input wire                            AP_AXIMM_36_AWVALID,
    output  wire                            AP_AXIMM_36_AWREADY,
    input wire [M_AXIMM_36_DATA_WIDTH-1:0]   AP_AXIMM_36_WDATA,
    input wire [M_AXIMM_36_DATA_WIDTH/8-1:0] AP_AXIMM_36_WSTRB,
    input wire                            AP_AXIMM_36_WLAST,
    input wire                            AP_AXIMM_36_WVALID,
    output  wire                            AP_AXIMM_36_WREADY,
    output  wire [1:0]                      AP_AXIMM_36_BRESP,
    output  wire                            AP_AXIMM_36_BVALID,
    input wire                            AP_AXIMM_36_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_36_ARADDR,
    input wire [7:0]                      AP_AXIMM_36_ARLEN,
    input wire [2:0]                      AP_AXIMM_36_ARSIZE,
    input wire [1:0]                      AP_AXIMM_36_ARBURST,
    input wire [1:0]                      AP_AXIMM_36_ARLOCK,
    input wire [3:0]                      AP_AXIMM_36_ARCACHE,
    input wire [2:0]                      AP_AXIMM_36_ARPROT,
    input wire [3:0]                      AP_AXIMM_36_ARREGION,
    input wire [3:0]                      AP_AXIMM_36_ARQOS,
    input wire                            AP_AXIMM_36_ARVALID,
    output  wire                            AP_AXIMM_36_ARREADY,
    output  wire [M_AXIMM_36_DATA_WIDTH-1:0]   AP_AXIMM_36_RDATA,
    output  wire [1:0]                      AP_AXIMM_36_RRESP,
    output  wire                            AP_AXIMM_36_RLAST,
    output  wire                            AP_AXIMM_36_RVALID,
    input  wire                            AP_AXIMM_36_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_36_AWADDR,
    output wire [7:0]                      M_AXIMM_36_AWLEN,
    output wire [2:0]                      M_AXIMM_36_AWSIZE,
    output wire [1:0]                      M_AXIMM_36_AWBURST,
    output wire [1:0]                      M_AXIMM_36_AWLOCK,
    output wire [3:0]                      M_AXIMM_36_AWCACHE,
    output wire [2:0]                      M_AXIMM_36_AWPROT,
    output wire [3:0]                      M_AXIMM_36_AWREGION,
    output wire [3:0]                      M_AXIMM_36_AWQOS,
    output wire                            M_AXIMM_36_AWVALID,
    input  wire                            M_AXIMM_36_AWREADY,
    output wire [M_AXIMM_36_DATA_WIDTH-1:0]   M_AXIMM_36_WDATA,
    output wire [M_AXIMM_36_DATA_WIDTH/8-1:0] M_AXIMM_36_WSTRB,
    output wire                            M_AXIMM_36_WLAST,
    output wire                            M_AXIMM_36_WVALID,
    input  wire                            M_AXIMM_36_WREADY,
    input  wire [1:0]                      M_AXIMM_36_BRESP,
    input  wire                            M_AXIMM_36_BVALID,
    output wire                            M_AXIMM_36_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_36_ARADDR,
    output wire [7:0]                      M_AXIMM_36_ARLEN,
    output wire [2:0]                      M_AXIMM_36_ARSIZE,
    output wire [1:0]                      M_AXIMM_36_ARBURST,
    output wire [1:0]                      M_AXIMM_36_ARLOCK,
    output wire [3:0]                      M_AXIMM_36_ARCACHE,
    output wire [2:0]                      M_AXIMM_36_ARPROT,
    output wire [3:0]                      M_AXIMM_36_ARREGION,
    output wire [3:0]                      M_AXIMM_36_ARQOS,
    output wire                            M_AXIMM_36_ARVALID,
    input  wire                            M_AXIMM_36_ARREADY,
    input  wire [M_AXIMM_36_DATA_WIDTH-1:0]   M_AXIMM_36_RDATA,
    input  wire [1:0]                      M_AXIMM_36_RRESP,
    input  wire                            M_AXIMM_36_RLAST,
    input  wire                            M_AXIMM_36_RVALID,
    output wire                            M_AXIMM_36_RREADY,
    //AXI-MM pass-through interface 37
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_37_AWADDR,
    input wire [7:0]                      AP_AXIMM_37_AWLEN,
    input wire [2:0]                      AP_AXIMM_37_AWSIZE,
    input wire [1:0]                      AP_AXIMM_37_AWBURST,
    input wire [1:0]                      AP_AXIMM_37_AWLOCK,
    input wire [3:0]                      AP_AXIMM_37_AWCACHE,
    input wire [2:0]                      AP_AXIMM_37_AWPROT,
    input wire [3:0]                      AP_AXIMM_37_AWREGION,
    input wire [3:0]                      AP_AXIMM_37_AWQOS,
    input wire                            AP_AXIMM_37_AWVALID,
    output  wire                            AP_AXIMM_37_AWREADY,
    input wire [M_AXIMM_37_DATA_WIDTH-1:0]   AP_AXIMM_37_WDATA,
    input wire [M_AXIMM_37_DATA_WIDTH/8-1:0] AP_AXIMM_37_WSTRB,
    input wire                            AP_AXIMM_37_WLAST,
    input wire                            AP_AXIMM_37_WVALID,
    output  wire                            AP_AXIMM_37_WREADY,
    output  wire [1:0]                      AP_AXIMM_37_BRESP,
    output  wire                            AP_AXIMM_37_BVALID,
    input wire                            AP_AXIMM_37_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_37_ARADDR,
    input wire [7:0]                      AP_AXIMM_37_ARLEN,
    input wire [2:0]                      AP_AXIMM_37_ARSIZE,
    input wire [1:0]                      AP_AXIMM_37_ARBURST,
    input wire [1:0]                      AP_AXIMM_37_ARLOCK,
    input wire [3:0]                      AP_AXIMM_37_ARCACHE,
    input wire [2:0]                      AP_AXIMM_37_ARPROT,
    input wire [3:0]                      AP_AXIMM_37_ARREGION,
    input wire [3:0]                      AP_AXIMM_37_ARQOS,
    input wire                            AP_AXIMM_37_ARVALID,
    output  wire                            AP_AXIMM_37_ARREADY,
    output  wire [M_AXIMM_37_DATA_WIDTH-1:0]   AP_AXIMM_37_RDATA,
    output  wire [1:0]                      AP_AXIMM_37_RRESP,
    output  wire                            AP_AXIMM_37_RLAST,
    output  wire                            AP_AXIMM_37_RVALID,
    input  wire                            AP_AXIMM_37_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_37_AWADDR,
    output wire [7:0]                      M_AXIMM_37_AWLEN,
    output wire [2:0]                      M_AXIMM_37_AWSIZE,
    output wire [1:0]                      M_AXIMM_37_AWBURST,
    output wire [1:0]                      M_AXIMM_37_AWLOCK,
    output wire [3:0]                      M_AXIMM_37_AWCACHE,
    output wire [2:0]                      M_AXIMM_37_AWPROT,
    output wire [3:0]                      M_AXIMM_37_AWREGION,
    output wire [3:0]                      M_AXIMM_37_AWQOS,
    output wire                            M_AXIMM_37_AWVALID,
    input  wire                            M_AXIMM_37_AWREADY,
    output wire [M_AXIMM_37_DATA_WIDTH-1:0]   M_AXIMM_37_WDATA,
    output wire [M_AXIMM_37_DATA_WIDTH/8-1:0] M_AXIMM_37_WSTRB,
    output wire                            M_AXIMM_37_WLAST,
    output wire                            M_AXIMM_37_WVALID,
    input  wire                            M_AXIMM_37_WREADY,
    input  wire [1:0]                      M_AXIMM_37_BRESP,
    input  wire                            M_AXIMM_37_BVALID,
    output wire                            M_AXIMM_37_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_37_ARADDR,
    output wire [7:0]                      M_AXIMM_37_ARLEN,
    output wire [2:0]                      M_AXIMM_37_ARSIZE,
    output wire [1:0]                      M_AXIMM_37_ARBURST,
    output wire [1:0]                      M_AXIMM_37_ARLOCK,
    output wire [3:0]                      M_AXIMM_37_ARCACHE,
    output wire [2:0]                      M_AXIMM_37_ARPROT,
    output wire [3:0]                      M_AXIMM_37_ARREGION,
    output wire [3:0]                      M_AXIMM_37_ARQOS,
    output wire                            M_AXIMM_37_ARVALID,
    input  wire                            M_AXIMM_37_ARREADY,
    input  wire [M_AXIMM_37_DATA_WIDTH-1:0]   M_AXIMM_37_RDATA,
    input  wire [1:0]                      M_AXIMM_37_RRESP,
    input  wire                            M_AXIMM_37_RLAST,
    input  wire                            M_AXIMM_37_RVALID,
    output wire                            M_AXIMM_37_RREADY,
    //AXI-MM pass-through interface 38
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_38_AWADDR,
    input wire [7:0]                      AP_AXIMM_38_AWLEN,
    input wire [2:0]                      AP_AXIMM_38_AWSIZE,
    input wire [1:0]                      AP_AXIMM_38_AWBURST,
    input wire [1:0]                      AP_AXIMM_38_AWLOCK,
    input wire [3:0]                      AP_AXIMM_38_AWCACHE,
    input wire [2:0]                      AP_AXIMM_38_AWPROT,
    input wire [3:0]                      AP_AXIMM_38_AWREGION,
    input wire [3:0]                      AP_AXIMM_38_AWQOS,
    input wire                            AP_AXIMM_38_AWVALID,
    output  wire                            AP_AXIMM_38_AWREADY,
    input wire [M_AXIMM_38_DATA_WIDTH-1:0]   AP_AXIMM_38_WDATA,
    input wire [M_AXIMM_38_DATA_WIDTH/8-1:0] AP_AXIMM_38_WSTRB,
    input wire                            AP_AXIMM_38_WLAST,
    input wire                            AP_AXIMM_38_WVALID,
    output  wire                            AP_AXIMM_38_WREADY,
    output  wire [1:0]                      AP_AXIMM_38_BRESP,
    output  wire                            AP_AXIMM_38_BVALID,
    input wire                            AP_AXIMM_38_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_38_ARADDR,
    input wire [7:0]                      AP_AXIMM_38_ARLEN,
    input wire [2:0]                      AP_AXIMM_38_ARSIZE,
    input wire [1:0]                      AP_AXIMM_38_ARBURST,
    input wire [1:0]                      AP_AXIMM_38_ARLOCK,
    input wire [3:0]                      AP_AXIMM_38_ARCACHE,
    input wire [2:0]                      AP_AXIMM_38_ARPROT,
    input wire [3:0]                      AP_AXIMM_38_ARREGION,
    input wire [3:0]                      AP_AXIMM_38_ARQOS,
    input wire                            AP_AXIMM_38_ARVALID,
    output  wire                            AP_AXIMM_38_ARREADY,
    output  wire [M_AXIMM_38_DATA_WIDTH-1:0]   AP_AXIMM_38_RDATA,
    output  wire [1:0]                      AP_AXIMM_38_RRESP,
    output  wire                            AP_AXIMM_38_RLAST,
    output  wire                            AP_AXIMM_38_RVALID,
    input  wire                            AP_AXIMM_38_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_38_AWADDR,
    output wire [7:0]                      M_AXIMM_38_AWLEN,
    output wire [2:0]                      M_AXIMM_38_AWSIZE,
    output wire [1:0]                      M_AXIMM_38_AWBURST,
    output wire [1:0]                      M_AXIMM_38_AWLOCK,
    output wire [3:0]                      M_AXIMM_38_AWCACHE,
    output wire [2:0]                      M_AXIMM_38_AWPROT,
    output wire [3:0]                      M_AXIMM_38_AWREGION,
    output wire [3:0]                      M_AXIMM_38_AWQOS,
    output wire                            M_AXIMM_38_AWVALID,
    input  wire                            M_AXIMM_38_AWREADY,
    output wire [M_AXIMM_38_DATA_WIDTH-1:0]   M_AXIMM_38_WDATA,
    output wire [M_AXIMM_38_DATA_WIDTH/8-1:0] M_AXIMM_38_WSTRB,
    output wire                            M_AXIMM_38_WLAST,
    output wire                            M_AXIMM_38_WVALID,
    input  wire                            M_AXIMM_38_WREADY,
    input  wire [1:0]                      M_AXIMM_38_BRESP,
    input  wire                            M_AXIMM_38_BVALID,
    output wire                            M_AXIMM_38_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_38_ARADDR,
    output wire [7:0]                      M_AXIMM_38_ARLEN,
    output wire [2:0]                      M_AXIMM_38_ARSIZE,
    output wire [1:0]                      M_AXIMM_38_ARBURST,
    output wire [1:0]                      M_AXIMM_38_ARLOCK,
    output wire [3:0]                      M_AXIMM_38_ARCACHE,
    output wire [2:0]                      M_AXIMM_38_ARPROT,
    output wire [3:0]                      M_AXIMM_38_ARREGION,
    output wire [3:0]                      M_AXIMM_38_ARQOS,
    output wire                            M_AXIMM_38_ARVALID,
    input  wire                            M_AXIMM_38_ARREADY,
    input  wire [M_AXIMM_38_DATA_WIDTH-1:0]   M_AXIMM_38_RDATA,
    input  wire [1:0]                      M_AXIMM_38_RRESP,
    input  wire                            M_AXIMM_38_RLAST,
    input  wire                            M_AXIMM_38_RVALID,
    output wire                            M_AXIMM_38_RREADY,
    //AXI-MM pass-through interface 39
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_39_AWADDR,
    input wire [7:0]                      AP_AXIMM_39_AWLEN,
    input wire [2:0]                      AP_AXIMM_39_AWSIZE,
    input wire [1:0]                      AP_AXIMM_39_AWBURST,
    input wire [1:0]                      AP_AXIMM_39_AWLOCK,
    input wire [3:0]                      AP_AXIMM_39_AWCACHE,
    input wire [2:0]                      AP_AXIMM_39_AWPROT,
    input wire [3:0]                      AP_AXIMM_39_AWREGION,
    input wire [3:0]                      AP_AXIMM_39_AWQOS,
    input wire                            AP_AXIMM_39_AWVALID,
    output  wire                            AP_AXIMM_39_AWREADY,
    input wire [M_AXIMM_39_DATA_WIDTH-1:0]   AP_AXIMM_39_WDATA,
    input wire [M_AXIMM_39_DATA_WIDTH/8-1:0] AP_AXIMM_39_WSTRB,
    input wire                            AP_AXIMM_39_WLAST,
    input wire                            AP_AXIMM_39_WVALID,
    output  wire                            AP_AXIMM_39_WREADY,
    output  wire [1:0]                      AP_AXIMM_39_BRESP,
    output  wire                            AP_AXIMM_39_BVALID,
    input wire                            AP_AXIMM_39_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_39_ARADDR,
    input wire [7:0]                      AP_AXIMM_39_ARLEN,
    input wire [2:0]                      AP_AXIMM_39_ARSIZE,
    input wire [1:0]                      AP_AXIMM_39_ARBURST,
    input wire [1:0]                      AP_AXIMM_39_ARLOCK,
    input wire [3:0]                      AP_AXIMM_39_ARCACHE,
    input wire [2:0]                      AP_AXIMM_39_ARPROT,
    input wire [3:0]                      AP_AXIMM_39_ARREGION,
    input wire [3:0]                      AP_AXIMM_39_ARQOS,
    input wire                            AP_AXIMM_39_ARVALID,
    output  wire                            AP_AXIMM_39_ARREADY,
    output  wire [M_AXIMM_39_DATA_WIDTH-1:0]   AP_AXIMM_39_RDATA,
    output  wire [1:0]                      AP_AXIMM_39_RRESP,
    output  wire                            AP_AXIMM_39_RLAST,
    output  wire                            AP_AXIMM_39_RVALID,
    input  wire                            AP_AXIMM_39_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_39_AWADDR,
    output wire [7:0]                      M_AXIMM_39_AWLEN,
    output wire [2:0]                      M_AXIMM_39_AWSIZE,
    output wire [1:0]                      M_AXIMM_39_AWBURST,
    output wire [1:0]                      M_AXIMM_39_AWLOCK,
    output wire [3:0]                      M_AXIMM_39_AWCACHE,
    output wire [2:0]                      M_AXIMM_39_AWPROT,
    output wire [3:0]                      M_AXIMM_39_AWREGION,
    output wire [3:0]                      M_AXIMM_39_AWQOS,
    output wire                            M_AXIMM_39_AWVALID,
    input  wire                            M_AXIMM_39_AWREADY,
    output wire [M_AXIMM_39_DATA_WIDTH-1:0]   M_AXIMM_39_WDATA,
    output wire [M_AXIMM_39_DATA_WIDTH/8-1:0] M_AXIMM_39_WSTRB,
    output wire                            M_AXIMM_39_WLAST,
    output wire                            M_AXIMM_39_WVALID,
    input  wire                            M_AXIMM_39_WREADY,
    input  wire [1:0]                      M_AXIMM_39_BRESP,
    input  wire                            M_AXIMM_39_BVALID,
    output wire                            M_AXIMM_39_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_39_ARADDR,
    output wire [7:0]                      M_AXIMM_39_ARLEN,
    output wire [2:0]                      M_AXIMM_39_ARSIZE,
    output wire [1:0]                      M_AXIMM_39_ARBURST,
    output wire [1:0]                      M_AXIMM_39_ARLOCK,
    output wire [3:0]                      M_AXIMM_39_ARCACHE,
    output wire [2:0]                      M_AXIMM_39_ARPROT,
    output wire [3:0]                      M_AXIMM_39_ARREGION,
    output wire [3:0]                      M_AXIMM_39_ARQOS,
    output wire                            M_AXIMM_39_ARVALID,
    input  wire                            M_AXIMM_39_ARREADY,
    input  wire [M_AXIMM_39_DATA_WIDTH-1:0]   M_AXIMM_39_RDATA,
    input  wire [1:0]                      M_AXIMM_39_RRESP,
    input  wire                            M_AXIMM_39_RLAST,
    input  wire                            M_AXIMM_39_RVALID,
    output wire                            M_AXIMM_39_RREADY,
    //AXI-MM pass-through interface 40
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_40_AWADDR,
    input wire [7:0]                      AP_AXIMM_40_AWLEN,
    input wire [2:0]                      AP_AXIMM_40_AWSIZE,
    input wire [1:0]                      AP_AXIMM_40_AWBURST,
    input wire [1:0]                      AP_AXIMM_40_AWLOCK,
    input wire [3:0]                      AP_AXIMM_40_AWCACHE,
    input wire [2:0]                      AP_AXIMM_40_AWPROT,
    input wire [3:0]                      AP_AXIMM_40_AWREGION,
    input wire [3:0]                      AP_AXIMM_40_AWQOS,
    input wire                            AP_AXIMM_40_AWVALID,
    output  wire                            AP_AXIMM_40_AWREADY,
    input wire [M_AXIMM_40_DATA_WIDTH-1:0]   AP_AXIMM_40_WDATA,
    input wire [M_AXIMM_40_DATA_WIDTH/8-1:0] AP_AXIMM_40_WSTRB,
    input wire                            AP_AXIMM_40_WLAST,
    input wire                            AP_AXIMM_40_WVALID,
    output  wire                            AP_AXIMM_40_WREADY,
    output  wire [1:0]                      AP_AXIMM_40_BRESP,
    output  wire                            AP_AXIMM_40_BVALID,
    input wire                            AP_AXIMM_40_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_40_ARADDR,
    input wire [7:0]                      AP_AXIMM_40_ARLEN,
    input wire [2:0]                      AP_AXIMM_40_ARSIZE,
    input wire [1:0]                      AP_AXIMM_40_ARBURST,
    input wire [1:0]                      AP_AXIMM_40_ARLOCK,
    input wire [3:0]                      AP_AXIMM_40_ARCACHE,
    input wire [2:0]                      AP_AXIMM_40_ARPROT,
    input wire [3:0]                      AP_AXIMM_40_ARREGION,
    input wire [3:0]                      AP_AXIMM_40_ARQOS,
    input wire                            AP_AXIMM_40_ARVALID,
    output  wire                            AP_AXIMM_40_ARREADY,
    output  wire [M_AXIMM_40_DATA_WIDTH-1:0]   AP_AXIMM_40_RDATA,
    output  wire [1:0]                      AP_AXIMM_40_RRESP,
    output  wire                            AP_AXIMM_40_RLAST,
    output  wire                            AP_AXIMM_40_RVALID,
    input  wire                            AP_AXIMM_40_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_40_AWADDR,
    output wire [7:0]                      M_AXIMM_40_AWLEN,
    output wire [2:0]                      M_AXIMM_40_AWSIZE,
    output wire [1:0]                      M_AXIMM_40_AWBURST,
    output wire [1:0]                      M_AXIMM_40_AWLOCK,
    output wire [3:0]                      M_AXIMM_40_AWCACHE,
    output wire [2:0]                      M_AXIMM_40_AWPROT,
    output wire [3:0]                      M_AXIMM_40_AWREGION,
    output wire [3:0]                      M_AXIMM_40_AWQOS,
    output wire                            M_AXIMM_40_AWVALID,
    input  wire                            M_AXIMM_40_AWREADY,
    output wire [M_AXIMM_40_DATA_WIDTH-1:0]   M_AXIMM_40_WDATA,
    output wire [M_AXIMM_40_DATA_WIDTH/8-1:0] M_AXIMM_40_WSTRB,
    output wire                            M_AXIMM_40_WLAST,
    output wire                            M_AXIMM_40_WVALID,
    input  wire                            M_AXIMM_40_WREADY,
    input  wire [1:0]                      M_AXIMM_40_BRESP,
    input  wire                            M_AXIMM_40_BVALID,
    output wire                            M_AXIMM_40_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_40_ARADDR,
    output wire [7:0]                      M_AXIMM_40_ARLEN,
    output wire [2:0]                      M_AXIMM_40_ARSIZE,
    output wire [1:0]                      M_AXIMM_40_ARBURST,
    output wire [1:0]                      M_AXIMM_40_ARLOCK,
    output wire [3:0]                      M_AXIMM_40_ARCACHE,
    output wire [2:0]                      M_AXIMM_40_ARPROT,
    output wire [3:0]                      M_AXIMM_40_ARREGION,
    output wire [3:0]                      M_AXIMM_40_ARQOS,
    output wire                            M_AXIMM_40_ARVALID,
    input  wire                            M_AXIMM_40_ARREADY,
    input  wire [M_AXIMM_40_DATA_WIDTH-1:0]   M_AXIMM_40_RDATA,
    input  wire [1:0]                      M_AXIMM_40_RRESP,
    input  wire                            M_AXIMM_40_RLAST,
    input  wire                            M_AXIMM_40_RVALID,
    output wire                            M_AXIMM_40_RREADY,
    //AXI-MM pass-through interface 41
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_41_AWADDR,
    input wire [7:0]                      AP_AXIMM_41_AWLEN,
    input wire [2:0]                      AP_AXIMM_41_AWSIZE,
    input wire [1:0]                      AP_AXIMM_41_AWBURST,
    input wire [1:0]                      AP_AXIMM_41_AWLOCK,
    input wire [3:0]                      AP_AXIMM_41_AWCACHE,
    input wire [2:0]                      AP_AXIMM_41_AWPROT,
    input wire [3:0]                      AP_AXIMM_41_AWREGION,
    input wire [3:0]                      AP_AXIMM_41_AWQOS,
    input wire                            AP_AXIMM_41_AWVALID,
    output  wire                            AP_AXIMM_41_AWREADY,
    input wire [M_AXIMM_41_DATA_WIDTH-1:0]   AP_AXIMM_41_WDATA,
    input wire [M_AXIMM_41_DATA_WIDTH/8-1:0] AP_AXIMM_41_WSTRB,
    input wire                            AP_AXIMM_41_WLAST,
    input wire                            AP_AXIMM_41_WVALID,
    output  wire                            AP_AXIMM_41_WREADY,
    output  wire [1:0]                      AP_AXIMM_41_BRESP,
    output  wire                            AP_AXIMM_41_BVALID,
    input wire                            AP_AXIMM_41_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_41_ARADDR,
    input wire [7:0]                      AP_AXIMM_41_ARLEN,
    input wire [2:0]                      AP_AXIMM_41_ARSIZE,
    input wire [1:0]                      AP_AXIMM_41_ARBURST,
    input wire [1:0]                      AP_AXIMM_41_ARLOCK,
    input wire [3:0]                      AP_AXIMM_41_ARCACHE,
    input wire [2:0]                      AP_AXIMM_41_ARPROT,
    input wire [3:0]                      AP_AXIMM_41_ARREGION,
    input wire [3:0]                      AP_AXIMM_41_ARQOS,
    input wire                            AP_AXIMM_41_ARVALID,
    output  wire                            AP_AXIMM_41_ARREADY,
    output  wire [M_AXIMM_41_DATA_WIDTH-1:0]   AP_AXIMM_41_RDATA,
    output  wire [1:0]                      AP_AXIMM_41_RRESP,
    output  wire                            AP_AXIMM_41_RLAST,
    output  wire                            AP_AXIMM_41_RVALID,
    input  wire                            AP_AXIMM_41_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_41_AWADDR,
    output wire [7:0]                      M_AXIMM_41_AWLEN,
    output wire [2:0]                      M_AXIMM_41_AWSIZE,
    output wire [1:0]                      M_AXIMM_41_AWBURST,
    output wire [1:0]                      M_AXIMM_41_AWLOCK,
    output wire [3:0]                      M_AXIMM_41_AWCACHE,
    output wire [2:0]                      M_AXIMM_41_AWPROT,
    output wire [3:0]                      M_AXIMM_41_AWREGION,
    output wire [3:0]                      M_AXIMM_41_AWQOS,
    output wire                            M_AXIMM_41_AWVALID,
    input  wire                            M_AXIMM_41_AWREADY,
    output wire [M_AXIMM_41_DATA_WIDTH-1:0]   M_AXIMM_41_WDATA,
    output wire [M_AXIMM_41_DATA_WIDTH/8-1:0] M_AXIMM_41_WSTRB,
    output wire                            M_AXIMM_41_WLAST,
    output wire                            M_AXIMM_41_WVALID,
    input  wire                            M_AXIMM_41_WREADY,
    input  wire [1:0]                      M_AXIMM_41_BRESP,
    input  wire                            M_AXIMM_41_BVALID,
    output wire                            M_AXIMM_41_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_41_ARADDR,
    output wire [7:0]                      M_AXIMM_41_ARLEN,
    output wire [2:0]                      M_AXIMM_41_ARSIZE,
    output wire [1:0]                      M_AXIMM_41_ARBURST,
    output wire [1:0]                      M_AXIMM_41_ARLOCK,
    output wire [3:0]                      M_AXIMM_41_ARCACHE,
    output wire [2:0]                      M_AXIMM_41_ARPROT,
    output wire [3:0]                      M_AXIMM_41_ARREGION,
    output wire [3:0]                      M_AXIMM_41_ARQOS,
    output wire                            M_AXIMM_41_ARVALID,
    input  wire                            M_AXIMM_41_ARREADY,
    input  wire [M_AXIMM_41_DATA_WIDTH-1:0]   M_AXIMM_41_RDATA,
    input  wire [1:0]                      M_AXIMM_41_RRESP,
    input  wire                            M_AXIMM_41_RLAST,
    input  wire                            M_AXIMM_41_RVALID,
    output wire                            M_AXIMM_41_RREADY,
    //AXI-MM pass-through interface 42
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_42_AWADDR,
    input wire [7:0]                      AP_AXIMM_42_AWLEN,
    input wire [2:0]                      AP_AXIMM_42_AWSIZE,
    input wire [1:0]                      AP_AXIMM_42_AWBURST,
    input wire [1:0]                      AP_AXIMM_42_AWLOCK,
    input wire [3:0]                      AP_AXIMM_42_AWCACHE,
    input wire [2:0]                      AP_AXIMM_42_AWPROT,
    input wire [3:0]                      AP_AXIMM_42_AWREGION,
    input wire [3:0]                      AP_AXIMM_42_AWQOS,
    input wire                            AP_AXIMM_42_AWVALID,
    output  wire                            AP_AXIMM_42_AWREADY,
    input wire [M_AXIMM_42_DATA_WIDTH-1:0]   AP_AXIMM_42_WDATA,
    input wire [M_AXIMM_42_DATA_WIDTH/8-1:0] AP_AXIMM_42_WSTRB,
    input wire                            AP_AXIMM_42_WLAST,
    input wire                            AP_AXIMM_42_WVALID,
    output  wire                            AP_AXIMM_42_WREADY,
    output  wire [1:0]                      AP_AXIMM_42_BRESP,
    output  wire                            AP_AXIMM_42_BVALID,
    input wire                            AP_AXIMM_42_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_42_ARADDR,
    input wire [7:0]                      AP_AXIMM_42_ARLEN,
    input wire [2:0]                      AP_AXIMM_42_ARSIZE,
    input wire [1:0]                      AP_AXIMM_42_ARBURST,
    input wire [1:0]                      AP_AXIMM_42_ARLOCK,
    input wire [3:0]                      AP_AXIMM_42_ARCACHE,
    input wire [2:0]                      AP_AXIMM_42_ARPROT,
    input wire [3:0]                      AP_AXIMM_42_ARREGION,
    input wire [3:0]                      AP_AXIMM_42_ARQOS,
    input wire                            AP_AXIMM_42_ARVALID,
    output  wire                            AP_AXIMM_42_ARREADY,
    output  wire [M_AXIMM_42_DATA_WIDTH-1:0]   AP_AXIMM_42_RDATA,
    output  wire [1:0]                      AP_AXIMM_42_RRESP,
    output  wire                            AP_AXIMM_42_RLAST,
    output  wire                            AP_AXIMM_42_RVALID,
    input  wire                            AP_AXIMM_42_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_42_AWADDR,
    output wire [7:0]                      M_AXIMM_42_AWLEN,
    output wire [2:0]                      M_AXIMM_42_AWSIZE,
    output wire [1:0]                      M_AXIMM_42_AWBURST,
    output wire [1:0]                      M_AXIMM_42_AWLOCK,
    output wire [3:0]                      M_AXIMM_42_AWCACHE,
    output wire [2:0]                      M_AXIMM_42_AWPROT,
    output wire [3:0]                      M_AXIMM_42_AWREGION,
    output wire [3:0]                      M_AXIMM_42_AWQOS,
    output wire                            M_AXIMM_42_AWVALID,
    input  wire                            M_AXIMM_42_AWREADY,
    output wire [M_AXIMM_42_DATA_WIDTH-1:0]   M_AXIMM_42_WDATA,
    output wire [M_AXIMM_42_DATA_WIDTH/8-1:0] M_AXIMM_42_WSTRB,
    output wire                            M_AXIMM_42_WLAST,
    output wire                            M_AXIMM_42_WVALID,
    input  wire                            M_AXIMM_42_WREADY,
    input  wire [1:0]                      M_AXIMM_42_BRESP,
    input  wire                            M_AXIMM_42_BVALID,
    output wire                            M_AXIMM_42_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_42_ARADDR,
    output wire [7:0]                      M_AXIMM_42_ARLEN,
    output wire [2:0]                      M_AXIMM_42_ARSIZE,
    output wire [1:0]                      M_AXIMM_42_ARBURST,
    output wire [1:0]                      M_AXIMM_42_ARLOCK,
    output wire [3:0]                      M_AXIMM_42_ARCACHE,
    output wire [2:0]                      M_AXIMM_42_ARPROT,
    output wire [3:0]                      M_AXIMM_42_ARREGION,
    output wire [3:0]                      M_AXIMM_42_ARQOS,
    output wire                            M_AXIMM_42_ARVALID,
    input  wire                            M_AXIMM_42_ARREADY,
    input  wire [M_AXIMM_42_DATA_WIDTH-1:0]   M_AXIMM_42_RDATA,
    input  wire [1:0]                      M_AXIMM_42_RRESP,
    input  wire                            M_AXIMM_42_RLAST,
    input  wire                            M_AXIMM_42_RVALID,
    output wire                            M_AXIMM_42_RREADY,
    //AXI-MM pass-through interface 43
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_43_AWADDR,
    input wire [7:0]                      AP_AXIMM_43_AWLEN,
    input wire [2:0]                      AP_AXIMM_43_AWSIZE,
    input wire [1:0]                      AP_AXIMM_43_AWBURST,
    input wire [1:0]                      AP_AXIMM_43_AWLOCK,
    input wire [3:0]                      AP_AXIMM_43_AWCACHE,
    input wire [2:0]                      AP_AXIMM_43_AWPROT,
    input wire [3:0]                      AP_AXIMM_43_AWREGION,
    input wire [3:0]                      AP_AXIMM_43_AWQOS,
    input wire                            AP_AXIMM_43_AWVALID,
    output  wire                            AP_AXIMM_43_AWREADY,
    input wire [M_AXIMM_43_DATA_WIDTH-1:0]   AP_AXIMM_43_WDATA,
    input wire [M_AXIMM_43_DATA_WIDTH/8-1:0] AP_AXIMM_43_WSTRB,
    input wire                            AP_AXIMM_43_WLAST,
    input wire                            AP_AXIMM_43_WVALID,
    output  wire                            AP_AXIMM_43_WREADY,
    output  wire [1:0]                      AP_AXIMM_43_BRESP,
    output  wire                            AP_AXIMM_43_BVALID,
    input wire                            AP_AXIMM_43_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_43_ARADDR,
    input wire [7:0]                      AP_AXIMM_43_ARLEN,
    input wire [2:0]                      AP_AXIMM_43_ARSIZE,
    input wire [1:0]                      AP_AXIMM_43_ARBURST,
    input wire [1:0]                      AP_AXIMM_43_ARLOCK,
    input wire [3:0]                      AP_AXIMM_43_ARCACHE,
    input wire [2:0]                      AP_AXIMM_43_ARPROT,
    input wire [3:0]                      AP_AXIMM_43_ARREGION,
    input wire [3:0]                      AP_AXIMM_43_ARQOS,
    input wire                            AP_AXIMM_43_ARVALID,
    output  wire                            AP_AXIMM_43_ARREADY,
    output  wire [M_AXIMM_43_DATA_WIDTH-1:0]   AP_AXIMM_43_RDATA,
    output  wire [1:0]                      AP_AXIMM_43_RRESP,
    output  wire                            AP_AXIMM_43_RLAST,
    output  wire                            AP_AXIMM_43_RVALID,
    input  wire                            AP_AXIMM_43_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_43_AWADDR,
    output wire [7:0]                      M_AXIMM_43_AWLEN,
    output wire [2:0]                      M_AXIMM_43_AWSIZE,
    output wire [1:0]                      M_AXIMM_43_AWBURST,
    output wire [1:0]                      M_AXIMM_43_AWLOCK,
    output wire [3:0]                      M_AXIMM_43_AWCACHE,
    output wire [2:0]                      M_AXIMM_43_AWPROT,
    output wire [3:0]                      M_AXIMM_43_AWREGION,
    output wire [3:0]                      M_AXIMM_43_AWQOS,
    output wire                            M_AXIMM_43_AWVALID,
    input  wire                            M_AXIMM_43_AWREADY,
    output wire [M_AXIMM_43_DATA_WIDTH-1:0]   M_AXIMM_43_WDATA,
    output wire [M_AXIMM_43_DATA_WIDTH/8-1:0] M_AXIMM_43_WSTRB,
    output wire                            M_AXIMM_43_WLAST,
    output wire                            M_AXIMM_43_WVALID,
    input  wire                            M_AXIMM_43_WREADY,
    input  wire [1:0]                      M_AXIMM_43_BRESP,
    input  wire                            M_AXIMM_43_BVALID,
    output wire                            M_AXIMM_43_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_43_ARADDR,
    output wire [7:0]                      M_AXIMM_43_ARLEN,
    output wire [2:0]                      M_AXIMM_43_ARSIZE,
    output wire [1:0]                      M_AXIMM_43_ARBURST,
    output wire [1:0]                      M_AXIMM_43_ARLOCK,
    output wire [3:0]                      M_AXIMM_43_ARCACHE,
    output wire [2:0]                      M_AXIMM_43_ARPROT,
    output wire [3:0]                      M_AXIMM_43_ARREGION,
    output wire [3:0]                      M_AXIMM_43_ARQOS,
    output wire                            M_AXIMM_43_ARVALID,
    input  wire                            M_AXIMM_43_ARREADY,
    input  wire [M_AXIMM_43_DATA_WIDTH-1:0]   M_AXIMM_43_RDATA,
    input  wire [1:0]                      M_AXIMM_43_RRESP,
    input  wire                            M_AXIMM_43_RLAST,
    input  wire                            M_AXIMM_43_RVALID,
    output wire                            M_AXIMM_43_RREADY,
    //AXI-MM pass-through interface 44
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_44_AWADDR,
    input wire [7:0]                      AP_AXIMM_44_AWLEN,
    input wire [2:0]                      AP_AXIMM_44_AWSIZE,
    input wire [1:0]                      AP_AXIMM_44_AWBURST,
    input wire [1:0]                      AP_AXIMM_44_AWLOCK,
    input wire [3:0]                      AP_AXIMM_44_AWCACHE,
    input wire [2:0]                      AP_AXIMM_44_AWPROT,
    input wire [3:0]                      AP_AXIMM_44_AWREGION,
    input wire [3:0]                      AP_AXIMM_44_AWQOS,
    input wire                            AP_AXIMM_44_AWVALID,
    output  wire                            AP_AXIMM_44_AWREADY,
    input wire [M_AXIMM_44_DATA_WIDTH-1:0]   AP_AXIMM_44_WDATA,
    input wire [M_AXIMM_44_DATA_WIDTH/8-1:0] AP_AXIMM_44_WSTRB,
    input wire                            AP_AXIMM_44_WLAST,
    input wire                            AP_AXIMM_44_WVALID,
    output  wire                            AP_AXIMM_44_WREADY,
    output  wire [1:0]                      AP_AXIMM_44_BRESP,
    output  wire                            AP_AXIMM_44_BVALID,
    input wire                            AP_AXIMM_44_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_44_ARADDR,
    input wire [7:0]                      AP_AXIMM_44_ARLEN,
    input wire [2:0]                      AP_AXIMM_44_ARSIZE,
    input wire [1:0]                      AP_AXIMM_44_ARBURST,
    input wire [1:0]                      AP_AXIMM_44_ARLOCK,
    input wire [3:0]                      AP_AXIMM_44_ARCACHE,
    input wire [2:0]                      AP_AXIMM_44_ARPROT,
    input wire [3:0]                      AP_AXIMM_44_ARREGION,
    input wire [3:0]                      AP_AXIMM_44_ARQOS,
    input wire                            AP_AXIMM_44_ARVALID,
    output  wire                            AP_AXIMM_44_ARREADY,
    output  wire [M_AXIMM_44_DATA_WIDTH-1:0]   AP_AXIMM_44_RDATA,
    output  wire [1:0]                      AP_AXIMM_44_RRESP,
    output  wire                            AP_AXIMM_44_RLAST,
    output  wire                            AP_AXIMM_44_RVALID,
    input  wire                            AP_AXIMM_44_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_44_AWADDR,
    output wire [7:0]                      M_AXIMM_44_AWLEN,
    output wire [2:0]                      M_AXIMM_44_AWSIZE,
    output wire [1:0]                      M_AXIMM_44_AWBURST,
    output wire [1:0]                      M_AXIMM_44_AWLOCK,
    output wire [3:0]                      M_AXIMM_44_AWCACHE,
    output wire [2:0]                      M_AXIMM_44_AWPROT,
    output wire [3:0]                      M_AXIMM_44_AWREGION,
    output wire [3:0]                      M_AXIMM_44_AWQOS,
    output wire                            M_AXIMM_44_AWVALID,
    input  wire                            M_AXIMM_44_AWREADY,
    output wire [M_AXIMM_44_DATA_WIDTH-1:0]   M_AXIMM_44_WDATA,
    output wire [M_AXIMM_44_DATA_WIDTH/8-1:0] M_AXIMM_44_WSTRB,
    output wire                            M_AXIMM_44_WLAST,
    output wire                            M_AXIMM_44_WVALID,
    input  wire                            M_AXIMM_44_WREADY,
    input  wire [1:0]                      M_AXIMM_44_BRESP,
    input  wire                            M_AXIMM_44_BVALID,
    output wire                            M_AXIMM_44_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_44_ARADDR,
    output wire [7:0]                      M_AXIMM_44_ARLEN,
    output wire [2:0]                      M_AXIMM_44_ARSIZE,
    output wire [1:0]                      M_AXIMM_44_ARBURST,
    output wire [1:0]                      M_AXIMM_44_ARLOCK,
    output wire [3:0]                      M_AXIMM_44_ARCACHE,
    output wire [2:0]                      M_AXIMM_44_ARPROT,
    output wire [3:0]                      M_AXIMM_44_ARREGION,
    output wire [3:0]                      M_AXIMM_44_ARQOS,
    output wire                            M_AXIMM_44_ARVALID,
    input  wire                            M_AXIMM_44_ARREADY,
    input  wire [M_AXIMM_44_DATA_WIDTH-1:0]   M_AXIMM_44_RDATA,
    input  wire [1:0]                      M_AXIMM_44_RRESP,
    input  wire                            M_AXIMM_44_RLAST,
    input  wire                            M_AXIMM_44_RVALID,
    output wire                            M_AXIMM_44_RREADY,
    //AXI-MM pass-through interface 45
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_45_AWADDR,
    input wire [7:0]                      AP_AXIMM_45_AWLEN,
    input wire [2:0]                      AP_AXIMM_45_AWSIZE,
    input wire [1:0]                      AP_AXIMM_45_AWBURST,
    input wire [1:0]                      AP_AXIMM_45_AWLOCK,
    input wire [3:0]                      AP_AXIMM_45_AWCACHE,
    input wire [2:0]                      AP_AXIMM_45_AWPROT,
    input wire [3:0]                      AP_AXIMM_45_AWREGION,
    input wire [3:0]                      AP_AXIMM_45_AWQOS,
    input wire                            AP_AXIMM_45_AWVALID,
    output  wire                            AP_AXIMM_45_AWREADY,
    input wire [M_AXIMM_45_DATA_WIDTH-1:0]   AP_AXIMM_45_WDATA,
    input wire [M_AXIMM_45_DATA_WIDTH/8-1:0] AP_AXIMM_45_WSTRB,
    input wire                            AP_AXIMM_45_WLAST,
    input wire                            AP_AXIMM_45_WVALID,
    output  wire                            AP_AXIMM_45_WREADY,
    output  wire [1:0]                      AP_AXIMM_45_BRESP,
    output  wire                            AP_AXIMM_45_BVALID,
    input wire                            AP_AXIMM_45_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_45_ARADDR,
    input wire [7:0]                      AP_AXIMM_45_ARLEN,
    input wire [2:0]                      AP_AXIMM_45_ARSIZE,
    input wire [1:0]                      AP_AXIMM_45_ARBURST,
    input wire [1:0]                      AP_AXIMM_45_ARLOCK,
    input wire [3:0]                      AP_AXIMM_45_ARCACHE,
    input wire [2:0]                      AP_AXIMM_45_ARPROT,
    input wire [3:0]                      AP_AXIMM_45_ARREGION,
    input wire [3:0]                      AP_AXIMM_45_ARQOS,
    input wire                            AP_AXIMM_45_ARVALID,
    output  wire                            AP_AXIMM_45_ARREADY,
    output  wire [M_AXIMM_45_DATA_WIDTH-1:0]   AP_AXIMM_45_RDATA,
    output  wire [1:0]                      AP_AXIMM_45_RRESP,
    output  wire                            AP_AXIMM_45_RLAST,
    output  wire                            AP_AXIMM_45_RVALID,
    input  wire                            AP_AXIMM_45_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_45_AWADDR,
    output wire [7:0]                      M_AXIMM_45_AWLEN,
    output wire [2:0]                      M_AXIMM_45_AWSIZE,
    output wire [1:0]                      M_AXIMM_45_AWBURST,
    output wire [1:0]                      M_AXIMM_45_AWLOCK,
    output wire [3:0]                      M_AXIMM_45_AWCACHE,
    output wire [2:0]                      M_AXIMM_45_AWPROT,
    output wire [3:0]                      M_AXIMM_45_AWREGION,
    output wire [3:0]                      M_AXIMM_45_AWQOS,
    output wire                            M_AXIMM_45_AWVALID,
    input  wire                            M_AXIMM_45_AWREADY,
    output wire [M_AXIMM_45_DATA_WIDTH-1:0]   M_AXIMM_45_WDATA,
    output wire [M_AXIMM_45_DATA_WIDTH/8-1:0] M_AXIMM_45_WSTRB,
    output wire                            M_AXIMM_45_WLAST,
    output wire                            M_AXIMM_45_WVALID,
    input  wire                            M_AXIMM_45_WREADY,
    input  wire [1:0]                      M_AXIMM_45_BRESP,
    input  wire                            M_AXIMM_45_BVALID,
    output wire                            M_AXIMM_45_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_45_ARADDR,
    output wire [7:0]                      M_AXIMM_45_ARLEN,
    output wire [2:0]                      M_AXIMM_45_ARSIZE,
    output wire [1:0]                      M_AXIMM_45_ARBURST,
    output wire [1:0]                      M_AXIMM_45_ARLOCK,
    output wire [3:0]                      M_AXIMM_45_ARCACHE,
    output wire [2:0]                      M_AXIMM_45_ARPROT,
    output wire [3:0]                      M_AXIMM_45_ARREGION,
    output wire [3:0]                      M_AXIMM_45_ARQOS,
    output wire                            M_AXIMM_45_ARVALID,
    input  wire                            M_AXIMM_45_ARREADY,
    input  wire [M_AXIMM_45_DATA_WIDTH-1:0]   M_AXIMM_45_RDATA,
    input  wire [1:0]                      M_AXIMM_45_RRESP,
    input  wire                            M_AXIMM_45_RLAST,
    input  wire                            M_AXIMM_45_RVALID,
    output wire                            M_AXIMM_45_RREADY,
    //AXI-MM pass-through interface 46
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_46_AWADDR,
    input wire [7:0]                      AP_AXIMM_46_AWLEN,
    input wire [2:0]                      AP_AXIMM_46_AWSIZE,
    input wire [1:0]                      AP_AXIMM_46_AWBURST,
    input wire [1:0]                      AP_AXIMM_46_AWLOCK,
    input wire [3:0]                      AP_AXIMM_46_AWCACHE,
    input wire [2:0]                      AP_AXIMM_46_AWPROT,
    input wire [3:0]                      AP_AXIMM_46_AWREGION,
    input wire [3:0]                      AP_AXIMM_46_AWQOS,
    input wire                            AP_AXIMM_46_AWVALID,
    output  wire                            AP_AXIMM_46_AWREADY,
    input wire [M_AXIMM_46_DATA_WIDTH-1:0]   AP_AXIMM_46_WDATA,
    input wire [M_AXIMM_46_DATA_WIDTH/8-1:0] AP_AXIMM_46_WSTRB,
    input wire                            AP_AXIMM_46_WLAST,
    input wire                            AP_AXIMM_46_WVALID,
    output  wire                            AP_AXIMM_46_WREADY,
    output  wire [1:0]                      AP_AXIMM_46_BRESP,
    output  wire                            AP_AXIMM_46_BVALID,
    input wire                            AP_AXIMM_46_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_46_ARADDR,
    input wire [7:0]                      AP_AXIMM_46_ARLEN,
    input wire [2:0]                      AP_AXIMM_46_ARSIZE,
    input wire [1:0]                      AP_AXIMM_46_ARBURST,
    input wire [1:0]                      AP_AXIMM_46_ARLOCK,
    input wire [3:0]                      AP_AXIMM_46_ARCACHE,
    input wire [2:0]                      AP_AXIMM_46_ARPROT,
    input wire [3:0]                      AP_AXIMM_46_ARREGION,
    input wire [3:0]                      AP_AXIMM_46_ARQOS,
    input wire                            AP_AXIMM_46_ARVALID,
    output  wire                            AP_AXIMM_46_ARREADY,
    output  wire [M_AXIMM_46_DATA_WIDTH-1:0]   AP_AXIMM_46_RDATA,
    output  wire [1:0]                      AP_AXIMM_46_RRESP,
    output  wire                            AP_AXIMM_46_RLAST,
    output  wire                            AP_AXIMM_46_RVALID,
    input  wire                            AP_AXIMM_46_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_46_AWADDR,
    output wire [7:0]                      M_AXIMM_46_AWLEN,
    output wire [2:0]                      M_AXIMM_46_AWSIZE,
    output wire [1:0]                      M_AXIMM_46_AWBURST,
    output wire [1:0]                      M_AXIMM_46_AWLOCK,
    output wire [3:0]                      M_AXIMM_46_AWCACHE,
    output wire [2:0]                      M_AXIMM_46_AWPROT,
    output wire [3:0]                      M_AXIMM_46_AWREGION,
    output wire [3:0]                      M_AXIMM_46_AWQOS,
    output wire                            M_AXIMM_46_AWVALID,
    input  wire                            M_AXIMM_46_AWREADY,
    output wire [M_AXIMM_46_DATA_WIDTH-1:0]   M_AXIMM_46_WDATA,
    output wire [M_AXIMM_46_DATA_WIDTH/8-1:0] M_AXIMM_46_WSTRB,
    output wire                            M_AXIMM_46_WLAST,
    output wire                            M_AXIMM_46_WVALID,
    input  wire                            M_AXIMM_46_WREADY,
    input  wire [1:0]                      M_AXIMM_46_BRESP,
    input  wire                            M_AXIMM_46_BVALID,
    output wire                            M_AXIMM_46_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_46_ARADDR,
    output wire [7:0]                      M_AXIMM_46_ARLEN,
    output wire [2:0]                      M_AXIMM_46_ARSIZE,
    output wire [1:0]                      M_AXIMM_46_ARBURST,
    output wire [1:0]                      M_AXIMM_46_ARLOCK,
    output wire [3:0]                      M_AXIMM_46_ARCACHE,
    output wire [2:0]                      M_AXIMM_46_ARPROT,
    output wire [3:0]                      M_AXIMM_46_ARREGION,
    output wire [3:0]                      M_AXIMM_46_ARQOS,
    output wire                            M_AXIMM_46_ARVALID,
    input  wire                            M_AXIMM_46_ARREADY,
    input  wire [M_AXIMM_46_DATA_WIDTH-1:0]   M_AXIMM_46_RDATA,
    input  wire [1:0]                      M_AXIMM_46_RRESP,
    input  wire                            M_AXIMM_46_RLAST,
    input  wire                            M_AXIMM_46_RVALID,
    output wire                            M_AXIMM_46_RREADY,
    //AXI-MM pass-through interface 47
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_47_AWADDR,
    input wire [7:0]                      AP_AXIMM_47_AWLEN,
    input wire [2:0]                      AP_AXIMM_47_AWSIZE,
    input wire [1:0]                      AP_AXIMM_47_AWBURST,
    input wire [1:0]                      AP_AXIMM_47_AWLOCK,
    input wire [3:0]                      AP_AXIMM_47_AWCACHE,
    input wire [2:0]                      AP_AXIMM_47_AWPROT,
    input wire [3:0]                      AP_AXIMM_47_AWREGION,
    input wire [3:0]                      AP_AXIMM_47_AWQOS,
    input wire                            AP_AXIMM_47_AWVALID,
    output  wire                            AP_AXIMM_47_AWREADY,
    input wire [M_AXIMM_47_DATA_WIDTH-1:0]   AP_AXIMM_47_WDATA,
    input wire [M_AXIMM_47_DATA_WIDTH/8-1:0] AP_AXIMM_47_WSTRB,
    input wire                            AP_AXIMM_47_WLAST,
    input wire                            AP_AXIMM_47_WVALID,
    output  wire                            AP_AXIMM_47_WREADY,
    output  wire [1:0]                      AP_AXIMM_47_BRESP,
    output  wire                            AP_AXIMM_47_BVALID,
    input wire                            AP_AXIMM_47_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_47_ARADDR,
    input wire [7:0]                      AP_AXIMM_47_ARLEN,
    input wire [2:0]                      AP_AXIMM_47_ARSIZE,
    input wire [1:0]                      AP_AXIMM_47_ARBURST,
    input wire [1:0]                      AP_AXIMM_47_ARLOCK,
    input wire [3:0]                      AP_AXIMM_47_ARCACHE,
    input wire [2:0]                      AP_AXIMM_47_ARPROT,
    input wire [3:0]                      AP_AXIMM_47_ARREGION,
    input wire [3:0]                      AP_AXIMM_47_ARQOS,
    input wire                            AP_AXIMM_47_ARVALID,
    output  wire                            AP_AXIMM_47_ARREADY,
    output  wire [M_AXIMM_47_DATA_WIDTH-1:0]   AP_AXIMM_47_RDATA,
    output  wire [1:0]                      AP_AXIMM_47_RRESP,
    output  wire                            AP_AXIMM_47_RLAST,
    output  wire                            AP_AXIMM_47_RVALID,
    input  wire                            AP_AXIMM_47_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_47_AWADDR,
    output wire [7:0]                      M_AXIMM_47_AWLEN,
    output wire [2:0]                      M_AXIMM_47_AWSIZE,
    output wire [1:0]                      M_AXIMM_47_AWBURST,
    output wire [1:0]                      M_AXIMM_47_AWLOCK,
    output wire [3:0]                      M_AXIMM_47_AWCACHE,
    output wire [2:0]                      M_AXIMM_47_AWPROT,
    output wire [3:0]                      M_AXIMM_47_AWREGION,
    output wire [3:0]                      M_AXIMM_47_AWQOS,
    output wire                            M_AXIMM_47_AWVALID,
    input  wire                            M_AXIMM_47_AWREADY,
    output wire [M_AXIMM_47_DATA_WIDTH-1:0]   M_AXIMM_47_WDATA,
    output wire [M_AXIMM_47_DATA_WIDTH/8-1:0] M_AXIMM_47_WSTRB,
    output wire                            M_AXIMM_47_WLAST,
    output wire                            M_AXIMM_47_WVALID,
    input  wire                            M_AXIMM_47_WREADY,
    input  wire [1:0]                      M_AXIMM_47_BRESP,
    input  wire                            M_AXIMM_47_BVALID,
    output wire                            M_AXIMM_47_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_47_ARADDR,
    output wire [7:0]                      M_AXIMM_47_ARLEN,
    output wire [2:0]                      M_AXIMM_47_ARSIZE,
    output wire [1:0]                      M_AXIMM_47_ARBURST,
    output wire [1:0]                      M_AXIMM_47_ARLOCK,
    output wire [3:0]                      M_AXIMM_47_ARCACHE,
    output wire [2:0]                      M_AXIMM_47_ARPROT,
    output wire [3:0]                      M_AXIMM_47_ARREGION,
    output wire [3:0]                      M_AXIMM_47_ARQOS,
    output wire                            M_AXIMM_47_ARVALID,
    input  wire                            M_AXIMM_47_ARREADY,
    input  wire [M_AXIMM_47_DATA_WIDTH-1:0]   M_AXIMM_47_RDATA,
    input  wire [1:0]                      M_AXIMM_47_RRESP,
    input  wire                            M_AXIMM_47_RLAST,
    input  wire                            M_AXIMM_47_RVALID,
    output wire                            M_AXIMM_47_RREADY,
    //AXI-MM pass-through interface 48
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_48_AWADDR,
    input wire [7:0]                      AP_AXIMM_48_AWLEN,
    input wire [2:0]                      AP_AXIMM_48_AWSIZE,
    input wire [1:0]                      AP_AXIMM_48_AWBURST,
    input wire [1:0]                      AP_AXIMM_48_AWLOCK,
    input wire [3:0]                      AP_AXIMM_48_AWCACHE,
    input wire [2:0]                      AP_AXIMM_48_AWPROT,
    input wire [3:0]                      AP_AXIMM_48_AWREGION,
    input wire [3:0]                      AP_AXIMM_48_AWQOS,
    input wire                            AP_AXIMM_48_AWVALID,
    output  wire                            AP_AXIMM_48_AWREADY,
    input wire [M_AXIMM_48_DATA_WIDTH-1:0]   AP_AXIMM_48_WDATA,
    input wire [M_AXIMM_48_DATA_WIDTH/8-1:0] AP_AXIMM_48_WSTRB,
    input wire                            AP_AXIMM_48_WLAST,
    input wire                            AP_AXIMM_48_WVALID,
    output  wire                            AP_AXIMM_48_WREADY,
    output  wire [1:0]                      AP_AXIMM_48_BRESP,
    output  wire                            AP_AXIMM_48_BVALID,
    input wire                            AP_AXIMM_48_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_48_ARADDR,
    input wire [7:0]                      AP_AXIMM_48_ARLEN,
    input wire [2:0]                      AP_AXIMM_48_ARSIZE,
    input wire [1:0]                      AP_AXIMM_48_ARBURST,
    input wire [1:0]                      AP_AXIMM_48_ARLOCK,
    input wire [3:0]                      AP_AXIMM_48_ARCACHE,
    input wire [2:0]                      AP_AXIMM_48_ARPROT,
    input wire [3:0]                      AP_AXIMM_48_ARREGION,
    input wire [3:0]                      AP_AXIMM_48_ARQOS,
    input wire                            AP_AXIMM_48_ARVALID,
    output  wire                            AP_AXIMM_48_ARREADY,
    output  wire [M_AXIMM_48_DATA_WIDTH-1:0]   AP_AXIMM_48_RDATA,
    output  wire [1:0]                      AP_AXIMM_48_RRESP,
    output  wire                            AP_AXIMM_48_RLAST,
    output  wire                            AP_AXIMM_48_RVALID,
    input  wire                            AP_AXIMM_48_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_48_AWADDR,
    output wire [7:0]                      M_AXIMM_48_AWLEN,
    output wire [2:0]                      M_AXIMM_48_AWSIZE,
    output wire [1:0]                      M_AXIMM_48_AWBURST,
    output wire [1:0]                      M_AXIMM_48_AWLOCK,
    output wire [3:0]                      M_AXIMM_48_AWCACHE,
    output wire [2:0]                      M_AXIMM_48_AWPROT,
    output wire [3:0]                      M_AXIMM_48_AWREGION,
    output wire [3:0]                      M_AXIMM_48_AWQOS,
    output wire                            M_AXIMM_48_AWVALID,
    input  wire                            M_AXIMM_48_AWREADY,
    output wire [M_AXIMM_48_DATA_WIDTH-1:0]   M_AXIMM_48_WDATA,
    output wire [M_AXIMM_48_DATA_WIDTH/8-1:0] M_AXIMM_48_WSTRB,
    output wire                            M_AXIMM_48_WLAST,
    output wire                            M_AXIMM_48_WVALID,
    input  wire                            M_AXIMM_48_WREADY,
    input  wire [1:0]                      M_AXIMM_48_BRESP,
    input  wire                            M_AXIMM_48_BVALID,
    output wire                            M_AXIMM_48_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_48_ARADDR,
    output wire [7:0]                      M_AXIMM_48_ARLEN,
    output wire [2:0]                      M_AXIMM_48_ARSIZE,
    output wire [1:0]                      M_AXIMM_48_ARBURST,
    output wire [1:0]                      M_AXIMM_48_ARLOCK,
    output wire [3:0]                      M_AXIMM_48_ARCACHE,
    output wire [2:0]                      M_AXIMM_48_ARPROT,
    output wire [3:0]                      M_AXIMM_48_ARREGION,
    output wire [3:0]                      M_AXIMM_48_ARQOS,
    output wire                            M_AXIMM_48_ARVALID,
    input  wire                            M_AXIMM_48_ARREADY,
    input  wire [M_AXIMM_48_DATA_WIDTH-1:0]   M_AXIMM_48_RDATA,
    input  wire [1:0]                      M_AXIMM_48_RRESP,
    input  wire                            M_AXIMM_48_RLAST,
    input  wire                            M_AXIMM_48_RVALID,
    output wire                            M_AXIMM_48_RREADY,
    //AXI-MM pass-through interface 49
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_49_AWADDR,
    input wire [7:0]                      AP_AXIMM_49_AWLEN,
    input wire [2:0]                      AP_AXIMM_49_AWSIZE,
    input wire [1:0]                      AP_AXIMM_49_AWBURST,
    input wire [1:0]                      AP_AXIMM_49_AWLOCK,
    input wire [3:0]                      AP_AXIMM_49_AWCACHE,
    input wire [2:0]                      AP_AXIMM_49_AWPROT,
    input wire [3:0]                      AP_AXIMM_49_AWREGION,
    input wire [3:0]                      AP_AXIMM_49_AWQOS,
    input wire                            AP_AXIMM_49_AWVALID,
    output  wire                            AP_AXIMM_49_AWREADY,
    input wire [M_AXIMM_49_DATA_WIDTH-1:0]   AP_AXIMM_49_WDATA,
    input wire [M_AXIMM_49_DATA_WIDTH/8-1:0] AP_AXIMM_49_WSTRB,
    input wire                            AP_AXIMM_49_WLAST,
    input wire                            AP_AXIMM_49_WVALID,
    output  wire                            AP_AXIMM_49_WREADY,
    output  wire [1:0]                      AP_AXIMM_49_BRESP,
    output  wire                            AP_AXIMM_49_BVALID,
    input wire                            AP_AXIMM_49_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_49_ARADDR,
    input wire [7:0]                      AP_AXIMM_49_ARLEN,
    input wire [2:0]                      AP_AXIMM_49_ARSIZE,
    input wire [1:0]                      AP_AXIMM_49_ARBURST,
    input wire [1:0]                      AP_AXIMM_49_ARLOCK,
    input wire [3:0]                      AP_AXIMM_49_ARCACHE,
    input wire [2:0]                      AP_AXIMM_49_ARPROT,
    input wire [3:0]                      AP_AXIMM_49_ARREGION,
    input wire [3:0]                      AP_AXIMM_49_ARQOS,
    input wire                            AP_AXIMM_49_ARVALID,
    output  wire                            AP_AXIMM_49_ARREADY,
    output  wire [M_AXIMM_49_DATA_WIDTH-1:0]   AP_AXIMM_49_RDATA,
    output  wire [1:0]                      AP_AXIMM_49_RRESP,
    output  wire                            AP_AXIMM_49_RLAST,
    output  wire                            AP_AXIMM_49_RVALID,
    input  wire                            AP_AXIMM_49_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_49_AWADDR,
    output wire [7:0]                      M_AXIMM_49_AWLEN,
    output wire [2:0]                      M_AXIMM_49_AWSIZE,
    output wire [1:0]                      M_AXIMM_49_AWBURST,
    output wire [1:0]                      M_AXIMM_49_AWLOCK,
    output wire [3:0]                      M_AXIMM_49_AWCACHE,
    output wire [2:0]                      M_AXIMM_49_AWPROT,
    output wire [3:0]                      M_AXIMM_49_AWREGION,
    output wire [3:0]                      M_AXIMM_49_AWQOS,
    output wire                            M_AXIMM_49_AWVALID,
    input  wire                            M_AXIMM_49_AWREADY,
    output wire [M_AXIMM_49_DATA_WIDTH-1:0]   M_AXIMM_49_WDATA,
    output wire [M_AXIMM_49_DATA_WIDTH/8-1:0] M_AXIMM_49_WSTRB,
    output wire                            M_AXIMM_49_WLAST,
    output wire                            M_AXIMM_49_WVALID,
    input  wire                            M_AXIMM_49_WREADY,
    input  wire [1:0]                      M_AXIMM_49_BRESP,
    input  wire                            M_AXIMM_49_BVALID,
    output wire                            M_AXIMM_49_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_49_ARADDR,
    output wire [7:0]                      M_AXIMM_49_ARLEN,
    output wire [2:0]                      M_AXIMM_49_ARSIZE,
    output wire [1:0]                      M_AXIMM_49_ARBURST,
    output wire [1:0]                      M_AXIMM_49_ARLOCK,
    output wire [3:0]                      M_AXIMM_49_ARCACHE,
    output wire [2:0]                      M_AXIMM_49_ARPROT,
    output wire [3:0]                      M_AXIMM_49_ARREGION,
    output wire [3:0]                      M_AXIMM_49_ARQOS,
    output wire                            M_AXIMM_49_ARVALID,
    input  wire                            M_AXIMM_49_ARREADY,
    input  wire [M_AXIMM_49_DATA_WIDTH-1:0]   M_AXIMM_49_RDATA,
    input  wire [1:0]                      M_AXIMM_49_RRESP,
    input  wire                            M_AXIMM_49_RLAST,
    input  wire                            M_AXIMM_49_RVALID,
    output wire                            M_AXIMM_49_RREADY,
    //AXI-MM pass-through interface 50
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_50_AWADDR,
    input wire [7:0]                      AP_AXIMM_50_AWLEN,
    input wire [2:0]                      AP_AXIMM_50_AWSIZE,
    input wire [1:0]                      AP_AXIMM_50_AWBURST,
    input wire [1:0]                      AP_AXIMM_50_AWLOCK,
    input wire [3:0]                      AP_AXIMM_50_AWCACHE,
    input wire [2:0]                      AP_AXIMM_50_AWPROT,
    input wire [3:0]                      AP_AXIMM_50_AWREGION,
    input wire [3:0]                      AP_AXIMM_50_AWQOS,
    input wire                            AP_AXIMM_50_AWVALID,
    output  wire                            AP_AXIMM_50_AWREADY,
    input wire [M_AXIMM_50_DATA_WIDTH-1:0]   AP_AXIMM_50_WDATA,
    input wire [M_AXIMM_50_DATA_WIDTH/8-1:0] AP_AXIMM_50_WSTRB,
    input wire                            AP_AXIMM_50_WLAST,
    input wire                            AP_AXIMM_50_WVALID,
    output  wire                            AP_AXIMM_50_WREADY,
    output  wire [1:0]                      AP_AXIMM_50_BRESP,
    output  wire                            AP_AXIMM_50_BVALID,
    input wire                            AP_AXIMM_50_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_50_ARADDR,
    input wire [7:0]                      AP_AXIMM_50_ARLEN,
    input wire [2:0]                      AP_AXIMM_50_ARSIZE,
    input wire [1:0]                      AP_AXIMM_50_ARBURST,
    input wire [1:0]                      AP_AXIMM_50_ARLOCK,
    input wire [3:0]                      AP_AXIMM_50_ARCACHE,
    input wire [2:0]                      AP_AXIMM_50_ARPROT,
    input wire [3:0]                      AP_AXIMM_50_ARREGION,
    input wire [3:0]                      AP_AXIMM_50_ARQOS,
    input wire                            AP_AXIMM_50_ARVALID,
    output  wire                            AP_AXIMM_50_ARREADY,
    output  wire [M_AXIMM_50_DATA_WIDTH-1:0]   AP_AXIMM_50_RDATA,
    output  wire [1:0]                      AP_AXIMM_50_RRESP,
    output  wire                            AP_AXIMM_50_RLAST,
    output  wire                            AP_AXIMM_50_RVALID,
    input  wire                            AP_AXIMM_50_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_50_AWADDR,
    output wire [7:0]                      M_AXIMM_50_AWLEN,
    output wire [2:0]                      M_AXIMM_50_AWSIZE,
    output wire [1:0]                      M_AXIMM_50_AWBURST,
    output wire [1:0]                      M_AXIMM_50_AWLOCK,
    output wire [3:0]                      M_AXIMM_50_AWCACHE,
    output wire [2:0]                      M_AXIMM_50_AWPROT,
    output wire [3:0]                      M_AXIMM_50_AWREGION,
    output wire [3:0]                      M_AXIMM_50_AWQOS,
    output wire                            M_AXIMM_50_AWVALID,
    input  wire                            M_AXIMM_50_AWREADY,
    output wire [M_AXIMM_50_DATA_WIDTH-1:0]   M_AXIMM_50_WDATA,
    output wire [M_AXIMM_50_DATA_WIDTH/8-1:0] M_AXIMM_50_WSTRB,
    output wire                            M_AXIMM_50_WLAST,
    output wire                            M_AXIMM_50_WVALID,
    input  wire                            M_AXIMM_50_WREADY,
    input  wire [1:0]                      M_AXIMM_50_BRESP,
    input  wire                            M_AXIMM_50_BVALID,
    output wire                            M_AXIMM_50_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_50_ARADDR,
    output wire [7:0]                      M_AXIMM_50_ARLEN,
    output wire [2:0]                      M_AXIMM_50_ARSIZE,
    output wire [1:0]                      M_AXIMM_50_ARBURST,
    output wire [1:0]                      M_AXIMM_50_ARLOCK,
    output wire [3:0]                      M_AXIMM_50_ARCACHE,
    output wire [2:0]                      M_AXIMM_50_ARPROT,
    output wire [3:0]                      M_AXIMM_50_ARREGION,
    output wire [3:0]                      M_AXIMM_50_ARQOS,
    output wire                            M_AXIMM_50_ARVALID,
    input  wire                            M_AXIMM_50_ARREADY,
    input  wire [M_AXIMM_50_DATA_WIDTH-1:0]   M_AXIMM_50_RDATA,
    input  wire [1:0]                      M_AXIMM_50_RRESP,
    input  wire                            M_AXIMM_50_RLAST,
    input  wire                            M_AXIMM_50_RVALID,
    output wire                            M_AXIMM_50_RREADY,
    //AXI-MM pass-through interface 51
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_51_AWADDR,
    input wire [7:0]                      AP_AXIMM_51_AWLEN,
    input wire [2:0]                      AP_AXIMM_51_AWSIZE,
    input wire [1:0]                      AP_AXIMM_51_AWBURST,
    input wire [1:0]                      AP_AXIMM_51_AWLOCK,
    input wire [3:0]                      AP_AXIMM_51_AWCACHE,
    input wire [2:0]                      AP_AXIMM_51_AWPROT,
    input wire [3:0]                      AP_AXIMM_51_AWREGION,
    input wire [3:0]                      AP_AXIMM_51_AWQOS,
    input wire                            AP_AXIMM_51_AWVALID,
    output  wire                            AP_AXIMM_51_AWREADY,
    input wire [M_AXIMM_51_DATA_WIDTH-1:0]   AP_AXIMM_51_WDATA,
    input wire [M_AXIMM_51_DATA_WIDTH/8-1:0] AP_AXIMM_51_WSTRB,
    input wire                            AP_AXIMM_51_WLAST,
    input wire                            AP_AXIMM_51_WVALID,
    output  wire                            AP_AXIMM_51_WREADY,
    output  wire [1:0]                      AP_AXIMM_51_BRESP,
    output  wire                            AP_AXIMM_51_BVALID,
    input wire                            AP_AXIMM_51_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_51_ARADDR,
    input wire [7:0]                      AP_AXIMM_51_ARLEN,
    input wire [2:0]                      AP_AXIMM_51_ARSIZE,
    input wire [1:0]                      AP_AXIMM_51_ARBURST,
    input wire [1:0]                      AP_AXIMM_51_ARLOCK,
    input wire [3:0]                      AP_AXIMM_51_ARCACHE,
    input wire [2:0]                      AP_AXIMM_51_ARPROT,
    input wire [3:0]                      AP_AXIMM_51_ARREGION,
    input wire [3:0]                      AP_AXIMM_51_ARQOS,
    input wire                            AP_AXIMM_51_ARVALID,
    output  wire                            AP_AXIMM_51_ARREADY,
    output  wire [M_AXIMM_51_DATA_WIDTH-1:0]   AP_AXIMM_51_RDATA,
    output  wire [1:0]                      AP_AXIMM_51_RRESP,
    output  wire                            AP_AXIMM_51_RLAST,
    output  wire                            AP_AXIMM_51_RVALID,
    input  wire                            AP_AXIMM_51_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_51_AWADDR,
    output wire [7:0]                      M_AXIMM_51_AWLEN,
    output wire [2:0]                      M_AXIMM_51_AWSIZE,
    output wire [1:0]                      M_AXIMM_51_AWBURST,
    output wire [1:0]                      M_AXIMM_51_AWLOCK,
    output wire [3:0]                      M_AXIMM_51_AWCACHE,
    output wire [2:0]                      M_AXIMM_51_AWPROT,
    output wire [3:0]                      M_AXIMM_51_AWREGION,
    output wire [3:0]                      M_AXIMM_51_AWQOS,
    output wire                            M_AXIMM_51_AWVALID,
    input  wire                            M_AXIMM_51_AWREADY,
    output wire [M_AXIMM_51_DATA_WIDTH-1:0]   M_AXIMM_51_WDATA,
    output wire [M_AXIMM_51_DATA_WIDTH/8-1:0] M_AXIMM_51_WSTRB,
    output wire                            M_AXIMM_51_WLAST,
    output wire                            M_AXIMM_51_WVALID,
    input  wire                            M_AXIMM_51_WREADY,
    input  wire [1:0]                      M_AXIMM_51_BRESP,
    input  wire                            M_AXIMM_51_BVALID,
    output wire                            M_AXIMM_51_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_51_ARADDR,
    output wire [7:0]                      M_AXIMM_51_ARLEN,
    output wire [2:0]                      M_AXIMM_51_ARSIZE,
    output wire [1:0]                      M_AXIMM_51_ARBURST,
    output wire [1:0]                      M_AXIMM_51_ARLOCK,
    output wire [3:0]                      M_AXIMM_51_ARCACHE,
    output wire [2:0]                      M_AXIMM_51_ARPROT,
    output wire [3:0]                      M_AXIMM_51_ARREGION,
    output wire [3:0]                      M_AXIMM_51_ARQOS,
    output wire                            M_AXIMM_51_ARVALID,
    input  wire                            M_AXIMM_51_ARREADY,
    input  wire [M_AXIMM_51_DATA_WIDTH-1:0]   M_AXIMM_51_RDATA,
    input  wire [1:0]                      M_AXIMM_51_RRESP,
    input  wire                            M_AXIMM_51_RLAST,
    input  wire                            M_AXIMM_51_RVALID,
    output wire                            M_AXIMM_51_RREADY,
    //AXI-MM pass-through interface 52
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_52_AWADDR,
    input wire [7:0]                      AP_AXIMM_52_AWLEN,
    input wire [2:0]                      AP_AXIMM_52_AWSIZE,
    input wire [1:0]                      AP_AXIMM_52_AWBURST,
    input wire [1:0]                      AP_AXIMM_52_AWLOCK,
    input wire [3:0]                      AP_AXIMM_52_AWCACHE,
    input wire [2:0]                      AP_AXIMM_52_AWPROT,
    input wire [3:0]                      AP_AXIMM_52_AWREGION,
    input wire [3:0]                      AP_AXIMM_52_AWQOS,
    input wire                            AP_AXIMM_52_AWVALID,
    output  wire                            AP_AXIMM_52_AWREADY,
    input wire [M_AXIMM_52_DATA_WIDTH-1:0]   AP_AXIMM_52_WDATA,
    input wire [M_AXIMM_52_DATA_WIDTH/8-1:0] AP_AXIMM_52_WSTRB,
    input wire                            AP_AXIMM_52_WLAST,
    input wire                            AP_AXIMM_52_WVALID,
    output  wire                            AP_AXIMM_52_WREADY,
    output  wire [1:0]                      AP_AXIMM_52_BRESP,
    output  wire                            AP_AXIMM_52_BVALID,
    input wire                            AP_AXIMM_52_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_52_ARADDR,
    input wire [7:0]                      AP_AXIMM_52_ARLEN,
    input wire [2:0]                      AP_AXIMM_52_ARSIZE,
    input wire [1:0]                      AP_AXIMM_52_ARBURST,
    input wire [1:0]                      AP_AXIMM_52_ARLOCK,
    input wire [3:0]                      AP_AXIMM_52_ARCACHE,
    input wire [2:0]                      AP_AXIMM_52_ARPROT,
    input wire [3:0]                      AP_AXIMM_52_ARREGION,
    input wire [3:0]                      AP_AXIMM_52_ARQOS,
    input wire                            AP_AXIMM_52_ARVALID,
    output  wire                            AP_AXIMM_52_ARREADY,
    output  wire [M_AXIMM_52_DATA_WIDTH-1:0]   AP_AXIMM_52_RDATA,
    output  wire [1:0]                      AP_AXIMM_52_RRESP,
    output  wire                            AP_AXIMM_52_RLAST,
    output  wire                            AP_AXIMM_52_RVALID,
    input  wire                            AP_AXIMM_52_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_52_AWADDR,
    output wire [7:0]                      M_AXIMM_52_AWLEN,
    output wire [2:0]                      M_AXIMM_52_AWSIZE,
    output wire [1:0]                      M_AXIMM_52_AWBURST,
    output wire [1:0]                      M_AXIMM_52_AWLOCK,
    output wire [3:0]                      M_AXIMM_52_AWCACHE,
    output wire [2:0]                      M_AXIMM_52_AWPROT,
    output wire [3:0]                      M_AXIMM_52_AWREGION,
    output wire [3:0]                      M_AXIMM_52_AWQOS,
    output wire                            M_AXIMM_52_AWVALID,
    input  wire                            M_AXIMM_52_AWREADY,
    output wire [M_AXIMM_52_DATA_WIDTH-1:0]   M_AXIMM_52_WDATA,
    output wire [M_AXIMM_52_DATA_WIDTH/8-1:0] M_AXIMM_52_WSTRB,
    output wire                            M_AXIMM_52_WLAST,
    output wire                            M_AXIMM_52_WVALID,
    input  wire                            M_AXIMM_52_WREADY,
    input  wire [1:0]                      M_AXIMM_52_BRESP,
    input  wire                            M_AXIMM_52_BVALID,
    output wire                            M_AXIMM_52_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_52_ARADDR,
    output wire [7:0]                      M_AXIMM_52_ARLEN,
    output wire [2:0]                      M_AXIMM_52_ARSIZE,
    output wire [1:0]                      M_AXIMM_52_ARBURST,
    output wire [1:0]                      M_AXIMM_52_ARLOCK,
    output wire [3:0]                      M_AXIMM_52_ARCACHE,
    output wire [2:0]                      M_AXIMM_52_ARPROT,
    output wire [3:0]                      M_AXIMM_52_ARREGION,
    output wire [3:0]                      M_AXIMM_52_ARQOS,
    output wire                            M_AXIMM_52_ARVALID,
    input  wire                            M_AXIMM_52_ARREADY,
    input  wire [M_AXIMM_52_DATA_WIDTH-1:0]   M_AXIMM_52_RDATA,
    input  wire [1:0]                      M_AXIMM_52_RRESP,
    input  wire                            M_AXIMM_52_RLAST,
    input  wire                            M_AXIMM_52_RVALID,
    output wire                            M_AXIMM_52_RREADY,
    //AXI-MM pass-through interface 53
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_53_AWADDR,
    input wire [7:0]                      AP_AXIMM_53_AWLEN,
    input wire [2:0]                      AP_AXIMM_53_AWSIZE,
    input wire [1:0]                      AP_AXIMM_53_AWBURST,
    input wire [1:0]                      AP_AXIMM_53_AWLOCK,
    input wire [3:0]                      AP_AXIMM_53_AWCACHE,
    input wire [2:0]                      AP_AXIMM_53_AWPROT,
    input wire [3:0]                      AP_AXIMM_53_AWREGION,
    input wire [3:0]                      AP_AXIMM_53_AWQOS,
    input wire                            AP_AXIMM_53_AWVALID,
    output  wire                            AP_AXIMM_53_AWREADY,
    input wire [M_AXIMM_53_DATA_WIDTH-1:0]   AP_AXIMM_53_WDATA,
    input wire [M_AXIMM_53_DATA_WIDTH/8-1:0] AP_AXIMM_53_WSTRB,
    input wire                            AP_AXIMM_53_WLAST,
    input wire                            AP_AXIMM_53_WVALID,
    output  wire                            AP_AXIMM_53_WREADY,
    output  wire [1:0]                      AP_AXIMM_53_BRESP,
    output  wire                            AP_AXIMM_53_BVALID,
    input wire                            AP_AXIMM_53_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_53_ARADDR,
    input wire [7:0]                      AP_AXIMM_53_ARLEN,
    input wire [2:0]                      AP_AXIMM_53_ARSIZE,
    input wire [1:0]                      AP_AXIMM_53_ARBURST,
    input wire [1:0]                      AP_AXIMM_53_ARLOCK,
    input wire [3:0]                      AP_AXIMM_53_ARCACHE,
    input wire [2:0]                      AP_AXIMM_53_ARPROT,
    input wire [3:0]                      AP_AXIMM_53_ARREGION,
    input wire [3:0]                      AP_AXIMM_53_ARQOS,
    input wire                            AP_AXIMM_53_ARVALID,
    output  wire                            AP_AXIMM_53_ARREADY,
    output  wire [M_AXIMM_53_DATA_WIDTH-1:0]   AP_AXIMM_53_RDATA,
    output  wire [1:0]                      AP_AXIMM_53_RRESP,
    output  wire                            AP_AXIMM_53_RLAST,
    output  wire                            AP_AXIMM_53_RVALID,
    input  wire                            AP_AXIMM_53_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_53_AWADDR,
    output wire [7:0]                      M_AXIMM_53_AWLEN,
    output wire [2:0]                      M_AXIMM_53_AWSIZE,
    output wire [1:0]                      M_AXIMM_53_AWBURST,
    output wire [1:0]                      M_AXIMM_53_AWLOCK,
    output wire [3:0]                      M_AXIMM_53_AWCACHE,
    output wire [2:0]                      M_AXIMM_53_AWPROT,
    output wire [3:0]                      M_AXIMM_53_AWREGION,
    output wire [3:0]                      M_AXIMM_53_AWQOS,
    output wire                            M_AXIMM_53_AWVALID,
    input  wire                            M_AXIMM_53_AWREADY,
    output wire [M_AXIMM_53_DATA_WIDTH-1:0]   M_AXIMM_53_WDATA,
    output wire [M_AXIMM_53_DATA_WIDTH/8-1:0] M_AXIMM_53_WSTRB,
    output wire                            M_AXIMM_53_WLAST,
    output wire                            M_AXIMM_53_WVALID,
    input  wire                            M_AXIMM_53_WREADY,
    input  wire [1:0]                      M_AXIMM_53_BRESP,
    input  wire                            M_AXIMM_53_BVALID,
    output wire                            M_AXIMM_53_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_53_ARADDR,
    output wire [7:0]                      M_AXIMM_53_ARLEN,
    output wire [2:0]                      M_AXIMM_53_ARSIZE,
    output wire [1:0]                      M_AXIMM_53_ARBURST,
    output wire [1:0]                      M_AXIMM_53_ARLOCK,
    output wire [3:0]                      M_AXIMM_53_ARCACHE,
    output wire [2:0]                      M_AXIMM_53_ARPROT,
    output wire [3:0]                      M_AXIMM_53_ARREGION,
    output wire [3:0]                      M_AXIMM_53_ARQOS,
    output wire                            M_AXIMM_53_ARVALID,
    input  wire                            M_AXIMM_53_ARREADY,
    input  wire [M_AXIMM_53_DATA_WIDTH-1:0]   M_AXIMM_53_RDATA,
    input  wire [1:0]                      M_AXIMM_53_RRESP,
    input  wire                            M_AXIMM_53_RLAST,
    input  wire                            M_AXIMM_53_RVALID,
    output wire                            M_AXIMM_53_RREADY,
    //AXI-MM pass-through interface 54
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_54_AWADDR,
    input wire [7:0]                      AP_AXIMM_54_AWLEN,
    input wire [2:0]                      AP_AXIMM_54_AWSIZE,
    input wire [1:0]                      AP_AXIMM_54_AWBURST,
    input wire [1:0]                      AP_AXIMM_54_AWLOCK,
    input wire [3:0]                      AP_AXIMM_54_AWCACHE,
    input wire [2:0]                      AP_AXIMM_54_AWPROT,
    input wire [3:0]                      AP_AXIMM_54_AWREGION,
    input wire [3:0]                      AP_AXIMM_54_AWQOS,
    input wire                            AP_AXIMM_54_AWVALID,
    output  wire                            AP_AXIMM_54_AWREADY,
    input wire [M_AXIMM_54_DATA_WIDTH-1:0]   AP_AXIMM_54_WDATA,
    input wire [M_AXIMM_54_DATA_WIDTH/8-1:0] AP_AXIMM_54_WSTRB,
    input wire                            AP_AXIMM_54_WLAST,
    input wire                            AP_AXIMM_54_WVALID,
    output  wire                            AP_AXIMM_54_WREADY,
    output  wire [1:0]                      AP_AXIMM_54_BRESP,
    output  wire                            AP_AXIMM_54_BVALID,
    input wire                            AP_AXIMM_54_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_54_ARADDR,
    input wire [7:0]                      AP_AXIMM_54_ARLEN,
    input wire [2:0]                      AP_AXIMM_54_ARSIZE,
    input wire [1:0]                      AP_AXIMM_54_ARBURST,
    input wire [1:0]                      AP_AXIMM_54_ARLOCK,
    input wire [3:0]                      AP_AXIMM_54_ARCACHE,
    input wire [2:0]                      AP_AXIMM_54_ARPROT,
    input wire [3:0]                      AP_AXIMM_54_ARREGION,
    input wire [3:0]                      AP_AXIMM_54_ARQOS,
    input wire                            AP_AXIMM_54_ARVALID,
    output  wire                            AP_AXIMM_54_ARREADY,
    output  wire [M_AXIMM_54_DATA_WIDTH-1:0]   AP_AXIMM_54_RDATA,
    output  wire [1:0]                      AP_AXIMM_54_RRESP,
    output  wire                            AP_AXIMM_54_RLAST,
    output  wire                            AP_AXIMM_54_RVALID,
    input  wire                            AP_AXIMM_54_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_54_AWADDR,
    output wire [7:0]                      M_AXIMM_54_AWLEN,
    output wire [2:0]                      M_AXIMM_54_AWSIZE,
    output wire [1:0]                      M_AXIMM_54_AWBURST,
    output wire [1:0]                      M_AXIMM_54_AWLOCK,
    output wire [3:0]                      M_AXIMM_54_AWCACHE,
    output wire [2:0]                      M_AXIMM_54_AWPROT,
    output wire [3:0]                      M_AXIMM_54_AWREGION,
    output wire [3:0]                      M_AXIMM_54_AWQOS,
    output wire                            M_AXIMM_54_AWVALID,
    input  wire                            M_AXIMM_54_AWREADY,
    output wire [M_AXIMM_54_DATA_WIDTH-1:0]   M_AXIMM_54_WDATA,
    output wire [M_AXIMM_54_DATA_WIDTH/8-1:0] M_AXIMM_54_WSTRB,
    output wire                            M_AXIMM_54_WLAST,
    output wire                            M_AXIMM_54_WVALID,
    input  wire                            M_AXIMM_54_WREADY,
    input  wire [1:0]                      M_AXIMM_54_BRESP,
    input  wire                            M_AXIMM_54_BVALID,
    output wire                            M_AXIMM_54_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_54_ARADDR,
    output wire [7:0]                      M_AXIMM_54_ARLEN,
    output wire [2:0]                      M_AXIMM_54_ARSIZE,
    output wire [1:0]                      M_AXIMM_54_ARBURST,
    output wire [1:0]                      M_AXIMM_54_ARLOCK,
    output wire [3:0]                      M_AXIMM_54_ARCACHE,
    output wire [2:0]                      M_AXIMM_54_ARPROT,
    output wire [3:0]                      M_AXIMM_54_ARREGION,
    output wire [3:0]                      M_AXIMM_54_ARQOS,
    output wire                            M_AXIMM_54_ARVALID,
    input  wire                            M_AXIMM_54_ARREADY,
    input  wire [M_AXIMM_54_DATA_WIDTH-1:0]   M_AXIMM_54_RDATA,
    input  wire [1:0]                      M_AXIMM_54_RRESP,
    input  wire                            M_AXIMM_54_RLAST,
    input  wire                            M_AXIMM_54_RVALID,
    output wire                            M_AXIMM_54_RREADY,
    //AXI-MM pass-through interface 55
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_55_AWADDR,
    input wire [7:0]                      AP_AXIMM_55_AWLEN,
    input wire [2:0]                      AP_AXIMM_55_AWSIZE,
    input wire [1:0]                      AP_AXIMM_55_AWBURST,
    input wire [1:0]                      AP_AXIMM_55_AWLOCK,
    input wire [3:0]                      AP_AXIMM_55_AWCACHE,
    input wire [2:0]                      AP_AXIMM_55_AWPROT,
    input wire [3:0]                      AP_AXIMM_55_AWREGION,
    input wire [3:0]                      AP_AXIMM_55_AWQOS,
    input wire                            AP_AXIMM_55_AWVALID,
    output  wire                            AP_AXIMM_55_AWREADY,
    input wire [M_AXIMM_55_DATA_WIDTH-1:0]   AP_AXIMM_55_WDATA,
    input wire [M_AXIMM_55_DATA_WIDTH/8-1:0] AP_AXIMM_55_WSTRB,
    input wire                            AP_AXIMM_55_WLAST,
    input wire                            AP_AXIMM_55_WVALID,
    output  wire                            AP_AXIMM_55_WREADY,
    output  wire [1:0]                      AP_AXIMM_55_BRESP,
    output  wire                            AP_AXIMM_55_BVALID,
    input wire                            AP_AXIMM_55_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_55_ARADDR,
    input wire [7:0]                      AP_AXIMM_55_ARLEN,
    input wire [2:0]                      AP_AXIMM_55_ARSIZE,
    input wire [1:0]                      AP_AXIMM_55_ARBURST,
    input wire [1:0]                      AP_AXIMM_55_ARLOCK,
    input wire [3:0]                      AP_AXIMM_55_ARCACHE,
    input wire [2:0]                      AP_AXIMM_55_ARPROT,
    input wire [3:0]                      AP_AXIMM_55_ARREGION,
    input wire [3:0]                      AP_AXIMM_55_ARQOS,
    input wire                            AP_AXIMM_55_ARVALID,
    output  wire                            AP_AXIMM_55_ARREADY,
    output  wire [M_AXIMM_55_DATA_WIDTH-1:0]   AP_AXIMM_55_RDATA,
    output  wire [1:0]                      AP_AXIMM_55_RRESP,
    output  wire                            AP_AXIMM_55_RLAST,
    output  wire                            AP_AXIMM_55_RVALID,
    input  wire                            AP_AXIMM_55_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_55_AWADDR,
    output wire [7:0]                      M_AXIMM_55_AWLEN,
    output wire [2:0]                      M_AXIMM_55_AWSIZE,
    output wire [1:0]                      M_AXIMM_55_AWBURST,
    output wire [1:0]                      M_AXIMM_55_AWLOCK,
    output wire [3:0]                      M_AXIMM_55_AWCACHE,
    output wire [2:0]                      M_AXIMM_55_AWPROT,
    output wire [3:0]                      M_AXIMM_55_AWREGION,
    output wire [3:0]                      M_AXIMM_55_AWQOS,
    output wire                            M_AXIMM_55_AWVALID,
    input  wire                            M_AXIMM_55_AWREADY,
    output wire [M_AXIMM_55_DATA_WIDTH-1:0]   M_AXIMM_55_WDATA,
    output wire [M_AXIMM_55_DATA_WIDTH/8-1:0] M_AXIMM_55_WSTRB,
    output wire                            M_AXIMM_55_WLAST,
    output wire                            M_AXIMM_55_WVALID,
    input  wire                            M_AXIMM_55_WREADY,
    input  wire [1:0]                      M_AXIMM_55_BRESP,
    input  wire                            M_AXIMM_55_BVALID,
    output wire                            M_AXIMM_55_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_55_ARADDR,
    output wire [7:0]                      M_AXIMM_55_ARLEN,
    output wire [2:0]                      M_AXIMM_55_ARSIZE,
    output wire [1:0]                      M_AXIMM_55_ARBURST,
    output wire [1:0]                      M_AXIMM_55_ARLOCK,
    output wire [3:0]                      M_AXIMM_55_ARCACHE,
    output wire [2:0]                      M_AXIMM_55_ARPROT,
    output wire [3:0]                      M_AXIMM_55_ARREGION,
    output wire [3:0]                      M_AXIMM_55_ARQOS,
    output wire                            M_AXIMM_55_ARVALID,
    input  wire                            M_AXIMM_55_ARREADY,
    input  wire [M_AXIMM_55_DATA_WIDTH-1:0]   M_AXIMM_55_RDATA,
    input  wire [1:0]                      M_AXIMM_55_RRESP,
    input  wire                            M_AXIMM_55_RLAST,
    input  wire                            M_AXIMM_55_RVALID,
    output wire                            M_AXIMM_55_RREADY,
    //AXI-MM pass-through interface 56
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_56_AWADDR,
    input wire [7:0]                      AP_AXIMM_56_AWLEN,
    input wire [2:0]                      AP_AXIMM_56_AWSIZE,
    input wire [1:0]                      AP_AXIMM_56_AWBURST,
    input wire [1:0]                      AP_AXIMM_56_AWLOCK,
    input wire [3:0]                      AP_AXIMM_56_AWCACHE,
    input wire [2:0]                      AP_AXIMM_56_AWPROT,
    input wire [3:0]                      AP_AXIMM_56_AWREGION,
    input wire [3:0]                      AP_AXIMM_56_AWQOS,
    input wire                            AP_AXIMM_56_AWVALID,
    output  wire                            AP_AXIMM_56_AWREADY,
    input wire [M_AXIMM_56_DATA_WIDTH-1:0]   AP_AXIMM_56_WDATA,
    input wire [M_AXIMM_56_DATA_WIDTH/8-1:0] AP_AXIMM_56_WSTRB,
    input wire                            AP_AXIMM_56_WLAST,
    input wire                            AP_AXIMM_56_WVALID,
    output  wire                            AP_AXIMM_56_WREADY,
    output  wire [1:0]                      AP_AXIMM_56_BRESP,
    output  wire                            AP_AXIMM_56_BVALID,
    input wire                            AP_AXIMM_56_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_56_ARADDR,
    input wire [7:0]                      AP_AXIMM_56_ARLEN,
    input wire [2:0]                      AP_AXIMM_56_ARSIZE,
    input wire [1:0]                      AP_AXIMM_56_ARBURST,
    input wire [1:0]                      AP_AXIMM_56_ARLOCK,
    input wire [3:0]                      AP_AXIMM_56_ARCACHE,
    input wire [2:0]                      AP_AXIMM_56_ARPROT,
    input wire [3:0]                      AP_AXIMM_56_ARREGION,
    input wire [3:0]                      AP_AXIMM_56_ARQOS,
    input wire                            AP_AXIMM_56_ARVALID,
    output  wire                            AP_AXIMM_56_ARREADY,
    output  wire [M_AXIMM_56_DATA_WIDTH-1:0]   AP_AXIMM_56_RDATA,
    output  wire [1:0]                      AP_AXIMM_56_RRESP,
    output  wire                            AP_AXIMM_56_RLAST,
    output  wire                            AP_AXIMM_56_RVALID,
    input  wire                            AP_AXIMM_56_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_56_AWADDR,
    output wire [7:0]                      M_AXIMM_56_AWLEN,
    output wire [2:0]                      M_AXIMM_56_AWSIZE,
    output wire [1:0]                      M_AXIMM_56_AWBURST,
    output wire [1:0]                      M_AXIMM_56_AWLOCK,
    output wire [3:0]                      M_AXIMM_56_AWCACHE,
    output wire [2:0]                      M_AXIMM_56_AWPROT,
    output wire [3:0]                      M_AXIMM_56_AWREGION,
    output wire [3:0]                      M_AXIMM_56_AWQOS,
    output wire                            M_AXIMM_56_AWVALID,
    input  wire                            M_AXIMM_56_AWREADY,
    output wire [M_AXIMM_56_DATA_WIDTH-1:0]   M_AXIMM_56_WDATA,
    output wire [M_AXIMM_56_DATA_WIDTH/8-1:0] M_AXIMM_56_WSTRB,
    output wire                            M_AXIMM_56_WLAST,
    output wire                            M_AXIMM_56_WVALID,
    input  wire                            M_AXIMM_56_WREADY,
    input  wire [1:0]                      M_AXIMM_56_BRESP,
    input  wire                            M_AXIMM_56_BVALID,
    output wire                            M_AXIMM_56_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_56_ARADDR,
    output wire [7:0]                      M_AXIMM_56_ARLEN,
    output wire [2:0]                      M_AXIMM_56_ARSIZE,
    output wire [1:0]                      M_AXIMM_56_ARBURST,
    output wire [1:0]                      M_AXIMM_56_ARLOCK,
    output wire [3:0]                      M_AXIMM_56_ARCACHE,
    output wire [2:0]                      M_AXIMM_56_ARPROT,
    output wire [3:0]                      M_AXIMM_56_ARREGION,
    output wire [3:0]                      M_AXIMM_56_ARQOS,
    output wire                            M_AXIMM_56_ARVALID,
    input  wire                            M_AXIMM_56_ARREADY,
    input  wire [M_AXIMM_56_DATA_WIDTH-1:0]   M_AXIMM_56_RDATA,
    input  wire [1:0]                      M_AXIMM_56_RRESP,
    input  wire                            M_AXIMM_56_RLAST,
    input  wire                            M_AXIMM_56_RVALID,
    output wire                            M_AXIMM_56_RREADY,
    //AXI-MM pass-through interface 57
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_57_AWADDR,
    input wire [7:0]                      AP_AXIMM_57_AWLEN,
    input wire [2:0]                      AP_AXIMM_57_AWSIZE,
    input wire [1:0]                      AP_AXIMM_57_AWBURST,
    input wire [1:0]                      AP_AXIMM_57_AWLOCK,
    input wire [3:0]                      AP_AXIMM_57_AWCACHE,
    input wire [2:0]                      AP_AXIMM_57_AWPROT,
    input wire [3:0]                      AP_AXIMM_57_AWREGION,
    input wire [3:0]                      AP_AXIMM_57_AWQOS,
    input wire                            AP_AXIMM_57_AWVALID,
    output  wire                            AP_AXIMM_57_AWREADY,
    input wire [M_AXIMM_57_DATA_WIDTH-1:0]   AP_AXIMM_57_WDATA,
    input wire [M_AXIMM_57_DATA_WIDTH/8-1:0] AP_AXIMM_57_WSTRB,
    input wire                            AP_AXIMM_57_WLAST,
    input wire                            AP_AXIMM_57_WVALID,
    output  wire                            AP_AXIMM_57_WREADY,
    output  wire [1:0]                      AP_AXIMM_57_BRESP,
    output  wire                            AP_AXIMM_57_BVALID,
    input wire                            AP_AXIMM_57_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_57_ARADDR,
    input wire [7:0]                      AP_AXIMM_57_ARLEN,
    input wire [2:0]                      AP_AXIMM_57_ARSIZE,
    input wire [1:0]                      AP_AXIMM_57_ARBURST,
    input wire [1:0]                      AP_AXIMM_57_ARLOCK,
    input wire [3:0]                      AP_AXIMM_57_ARCACHE,
    input wire [2:0]                      AP_AXIMM_57_ARPROT,
    input wire [3:0]                      AP_AXIMM_57_ARREGION,
    input wire [3:0]                      AP_AXIMM_57_ARQOS,
    input wire                            AP_AXIMM_57_ARVALID,
    output  wire                            AP_AXIMM_57_ARREADY,
    output  wire [M_AXIMM_57_DATA_WIDTH-1:0]   AP_AXIMM_57_RDATA,
    output  wire [1:0]                      AP_AXIMM_57_RRESP,
    output  wire                            AP_AXIMM_57_RLAST,
    output  wire                            AP_AXIMM_57_RVALID,
    input  wire                            AP_AXIMM_57_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_57_AWADDR,
    output wire [7:0]                      M_AXIMM_57_AWLEN,
    output wire [2:0]                      M_AXIMM_57_AWSIZE,
    output wire [1:0]                      M_AXIMM_57_AWBURST,
    output wire [1:0]                      M_AXIMM_57_AWLOCK,
    output wire [3:0]                      M_AXIMM_57_AWCACHE,
    output wire [2:0]                      M_AXIMM_57_AWPROT,
    output wire [3:0]                      M_AXIMM_57_AWREGION,
    output wire [3:0]                      M_AXIMM_57_AWQOS,
    output wire                            M_AXIMM_57_AWVALID,
    input  wire                            M_AXIMM_57_AWREADY,
    output wire [M_AXIMM_57_DATA_WIDTH-1:0]   M_AXIMM_57_WDATA,
    output wire [M_AXIMM_57_DATA_WIDTH/8-1:0] M_AXIMM_57_WSTRB,
    output wire                            M_AXIMM_57_WLAST,
    output wire                            M_AXIMM_57_WVALID,
    input  wire                            M_AXIMM_57_WREADY,
    input  wire [1:0]                      M_AXIMM_57_BRESP,
    input  wire                            M_AXIMM_57_BVALID,
    output wire                            M_AXIMM_57_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_57_ARADDR,
    output wire [7:0]                      M_AXIMM_57_ARLEN,
    output wire [2:0]                      M_AXIMM_57_ARSIZE,
    output wire [1:0]                      M_AXIMM_57_ARBURST,
    output wire [1:0]                      M_AXIMM_57_ARLOCK,
    output wire [3:0]                      M_AXIMM_57_ARCACHE,
    output wire [2:0]                      M_AXIMM_57_ARPROT,
    output wire [3:0]                      M_AXIMM_57_ARREGION,
    output wire [3:0]                      M_AXIMM_57_ARQOS,
    output wire                            M_AXIMM_57_ARVALID,
    input  wire                            M_AXIMM_57_ARREADY,
    input  wire [M_AXIMM_57_DATA_WIDTH-1:0]   M_AXIMM_57_RDATA,
    input  wire [1:0]                      M_AXIMM_57_RRESP,
    input  wire                            M_AXIMM_57_RLAST,
    input  wire                            M_AXIMM_57_RVALID,
    output wire                            M_AXIMM_57_RREADY,
    //AXI-MM pass-through interface 58
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_58_AWADDR,
    input wire [7:0]                      AP_AXIMM_58_AWLEN,
    input wire [2:0]                      AP_AXIMM_58_AWSIZE,
    input wire [1:0]                      AP_AXIMM_58_AWBURST,
    input wire [1:0]                      AP_AXIMM_58_AWLOCK,
    input wire [3:0]                      AP_AXIMM_58_AWCACHE,
    input wire [2:0]                      AP_AXIMM_58_AWPROT,
    input wire [3:0]                      AP_AXIMM_58_AWREGION,
    input wire [3:0]                      AP_AXIMM_58_AWQOS,
    input wire                            AP_AXIMM_58_AWVALID,
    output  wire                            AP_AXIMM_58_AWREADY,
    input wire [M_AXIMM_58_DATA_WIDTH-1:0]   AP_AXIMM_58_WDATA,
    input wire [M_AXIMM_58_DATA_WIDTH/8-1:0] AP_AXIMM_58_WSTRB,
    input wire                            AP_AXIMM_58_WLAST,
    input wire                            AP_AXIMM_58_WVALID,
    output  wire                            AP_AXIMM_58_WREADY,
    output  wire [1:0]                      AP_AXIMM_58_BRESP,
    output  wire                            AP_AXIMM_58_BVALID,
    input wire                            AP_AXIMM_58_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_58_ARADDR,
    input wire [7:0]                      AP_AXIMM_58_ARLEN,
    input wire [2:0]                      AP_AXIMM_58_ARSIZE,
    input wire [1:0]                      AP_AXIMM_58_ARBURST,
    input wire [1:0]                      AP_AXIMM_58_ARLOCK,
    input wire [3:0]                      AP_AXIMM_58_ARCACHE,
    input wire [2:0]                      AP_AXIMM_58_ARPROT,
    input wire [3:0]                      AP_AXIMM_58_ARREGION,
    input wire [3:0]                      AP_AXIMM_58_ARQOS,
    input wire                            AP_AXIMM_58_ARVALID,
    output  wire                            AP_AXIMM_58_ARREADY,
    output  wire [M_AXIMM_58_DATA_WIDTH-1:0]   AP_AXIMM_58_RDATA,
    output  wire [1:0]                      AP_AXIMM_58_RRESP,
    output  wire                            AP_AXIMM_58_RLAST,
    output  wire                            AP_AXIMM_58_RVALID,
    input  wire                            AP_AXIMM_58_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_58_AWADDR,
    output wire [7:0]                      M_AXIMM_58_AWLEN,
    output wire [2:0]                      M_AXIMM_58_AWSIZE,
    output wire [1:0]                      M_AXIMM_58_AWBURST,
    output wire [1:0]                      M_AXIMM_58_AWLOCK,
    output wire [3:0]                      M_AXIMM_58_AWCACHE,
    output wire [2:0]                      M_AXIMM_58_AWPROT,
    output wire [3:0]                      M_AXIMM_58_AWREGION,
    output wire [3:0]                      M_AXIMM_58_AWQOS,
    output wire                            M_AXIMM_58_AWVALID,
    input  wire                            M_AXIMM_58_AWREADY,
    output wire [M_AXIMM_58_DATA_WIDTH-1:0]   M_AXIMM_58_WDATA,
    output wire [M_AXIMM_58_DATA_WIDTH/8-1:0] M_AXIMM_58_WSTRB,
    output wire                            M_AXIMM_58_WLAST,
    output wire                            M_AXIMM_58_WVALID,
    input  wire                            M_AXIMM_58_WREADY,
    input  wire [1:0]                      M_AXIMM_58_BRESP,
    input  wire                            M_AXIMM_58_BVALID,
    output wire                            M_AXIMM_58_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_58_ARADDR,
    output wire [7:0]                      M_AXIMM_58_ARLEN,
    output wire [2:0]                      M_AXIMM_58_ARSIZE,
    output wire [1:0]                      M_AXIMM_58_ARBURST,
    output wire [1:0]                      M_AXIMM_58_ARLOCK,
    output wire [3:0]                      M_AXIMM_58_ARCACHE,
    output wire [2:0]                      M_AXIMM_58_ARPROT,
    output wire [3:0]                      M_AXIMM_58_ARREGION,
    output wire [3:0]                      M_AXIMM_58_ARQOS,
    output wire                            M_AXIMM_58_ARVALID,
    input  wire                            M_AXIMM_58_ARREADY,
    input  wire [M_AXIMM_58_DATA_WIDTH-1:0]   M_AXIMM_58_RDATA,
    input  wire [1:0]                      M_AXIMM_58_RRESP,
    input  wire                            M_AXIMM_58_RLAST,
    input  wire                            M_AXIMM_58_RVALID,
    output wire                            M_AXIMM_58_RREADY,
    //AXI-MM pass-through interface 59
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_59_AWADDR,
    input wire [7:0]                      AP_AXIMM_59_AWLEN,
    input wire [2:0]                      AP_AXIMM_59_AWSIZE,
    input wire [1:0]                      AP_AXIMM_59_AWBURST,
    input wire [1:0]                      AP_AXIMM_59_AWLOCK,
    input wire [3:0]                      AP_AXIMM_59_AWCACHE,
    input wire [2:0]                      AP_AXIMM_59_AWPROT,
    input wire [3:0]                      AP_AXIMM_59_AWREGION,
    input wire [3:0]                      AP_AXIMM_59_AWQOS,
    input wire                            AP_AXIMM_59_AWVALID,
    output  wire                            AP_AXIMM_59_AWREADY,
    input wire [M_AXIMM_59_DATA_WIDTH-1:0]   AP_AXIMM_59_WDATA,
    input wire [M_AXIMM_59_DATA_WIDTH/8-1:0] AP_AXIMM_59_WSTRB,
    input wire                            AP_AXIMM_59_WLAST,
    input wire                            AP_AXIMM_59_WVALID,
    output  wire                            AP_AXIMM_59_WREADY,
    output  wire [1:0]                      AP_AXIMM_59_BRESP,
    output  wire                            AP_AXIMM_59_BVALID,
    input wire                            AP_AXIMM_59_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_59_ARADDR,
    input wire [7:0]                      AP_AXIMM_59_ARLEN,
    input wire [2:0]                      AP_AXIMM_59_ARSIZE,
    input wire [1:0]                      AP_AXIMM_59_ARBURST,
    input wire [1:0]                      AP_AXIMM_59_ARLOCK,
    input wire [3:0]                      AP_AXIMM_59_ARCACHE,
    input wire [2:0]                      AP_AXIMM_59_ARPROT,
    input wire [3:0]                      AP_AXIMM_59_ARREGION,
    input wire [3:0]                      AP_AXIMM_59_ARQOS,
    input wire                            AP_AXIMM_59_ARVALID,
    output  wire                            AP_AXIMM_59_ARREADY,
    output  wire [M_AXIMM_59_DATA_WIDTH-1:0]   AP_AXIMM_59_RDATA,
    output  wire [1:0]                      AP_AXIMM_59_RRESP,
    output  wire                            AP_AXIMM_59_RLAST,
    output  wire                            AP_AXIMM_59_RVALID,
    input  wire                            AP_AXIMM_59_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_59_AWADDR,
    output wire [7:0]                      M_AXIMM_59_AWLEN,
    output wire [2:0]                      M_AXIMM_59_AWSIZE,
    output wire [1:0]                      M_AXIMM_59_AWBURST,
    output wire [1:0]                      M_AXIMM_59_AWLOCK,
    output wire [3:0]                      M_AXIMM_59_AWCACHE,
    output wire [2:0]                      M_AXIMM_59_AWPROT,
    output wire [3:0]                      M_AXIMM_59_AWREGION,
    output wire [3:0]                      M_AXIMM_59_AWQOS,
    output wire                            M_AXIMM_59_AWVALID,
    input  wire                            M_AXIMM_59_AWREADY,
    output wire [M_AXIMM_59_DATA_WIDTH-1:0]   M_AXIMM_59_WDATA,
    output wire [M_AXIMM_59_DATA_WIDTH/8-1:0] M_AXIMM_59_WSTRB,
    output wire                            M_AXIMM_59_WLAST,
    output wire                            M_AXIMM_59_WVALID,
    input  wire                            M_AXIMM_59_WREADY,
    input  wire [1:0]                      M_AXIMM_59_BRESP,
    input  wire                            M_AXIMM_59_BVALID,
    output wire                            M_AXIMM_59_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_59_ARADDR,
    output wire [7:0]                      M_AXIMM_59_ARLEN,
    output wire [2:0]                      M_AXIMM_59_ARSIZE,
    output wire [1:0]                      M_AXIMM_59_ARBURST,
    output wire [1:0]                      M_AXIMM_59_ARLOCK,
    output wire [3:0]                      M_AXIMM_59_ARCACHE,
    output wire [2:0]                      M_AXIMM_59_ARPROT,
    output wire [3:0]                      M_AXIMM_59_ARREGION,
    output wire [3:0]                      M_AXIMM_59_ARQOS,
    output wire                            M_AXIMM_59_ARVALID,
    input  wire                            M_AXIMM_59_ARREADY,
    input  wire [M_AXIMM_59_DATA_WIDTH-1:0]   M_AXIMM_59_RDATA,
    input  wire [1:0]                      M_AXIMM_59_RRESP,
    input  wire                            M_AXIMM_59_RLAST,
    input  wire                            M_AXIMM_59_RVALID,
    output wire                            M_AXIMM_59_RREADY,
    //AXI-MM pass-through interface 60
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_60_AWADDR,
    input wire [7:0]                      AP_AXIMM_60_AWLEN,
    input wire [2:0]                      AP_AXIMM_60_AWSIZE,
    input wire [1:0]                      AP_AXIMM_60_AWBURST,
    input wire [1:0]                      AP_AXIMM_60_AWLOCK,
    input wire [3:0]                      AP_AXIMM_60_AWCACHE,
    input wire [2:0]                      AP_AXIMM_60_AWPROT,
    input wire [3:0]                      AP_AXIMM_60_AWREGION,
    input wire [3:0]                      AP_AXIMM_60_AWQOS,
    input wire                            AP_AXIMM_60_AWVALID,
    output  wire                            AP_AXIMM_60_AWREADY,
    input wire [M_AXIMM_60_DATA_WIDTH-1:0]   AP_AXIMM_60_WDATA,
    input wire [M_AXIMM_60_DATA_WIDTH/8-1:0] AP_AXIMM_60_WSTRB,
    input wire                            AP_AXIMM_60_WLAST,
    input wire                            AP_AXIMM_60_WVALID,
    output  wire                            AP_AXIMM_60_WREADY,
    output  wire [1:0]                      AP_AXIMM_60_BRESP,
    output  wire                            AP_AXIMM_60_BVALID,
    input wire                            AP_AXIMM_60_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_60_ARADDR,
    input wire [7:0]                      AP_AXIMM_60_ARLEN,
    input wire [2:0]                      AP_AXIMM_60_ARSIZE,
    input wire [1:0]                      AP_AXIMM_60_ARBURST,
    input wire [1:0]                      AP_AXIMM_60_ARLOCK,
    input wire [3:0]                      AP_AXIMM_60_ARCACHE,
    input wire [2:0]                      AP_AXIMM_60_ARPROT,
    input wire [3:0]                      AP_AXIMM_60_ARREGION,
    input wire [3:0]                      AP_AXIMM_60_ARQOS,
    input wire                            AP_AXIMM_60_ARVALID,
    output  wire                            AP_AXIMM_60_ARREADY,
    output  wire [M_AXIMM_60_DATA_WIDTH-1:0]   AP_AXIMM_60_RDATA,
    output  wire [1:0]                      AP_AXIMM_60_RRESP,
    output  wire                            AP_AXIMM_60_RLAST,
    output  wire                            AP_AXIMM_60_RVALID,
    input  wire                            AP_AXIMM_60_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_60_AWADDR,
    output wire [7:0]                      M_AXIMM_60_AWLEN,
    output wire [2:0]                      M_AXIMM_60_AWSIZE,
    output wire [1:0]                      M_AXIMM_60_AWBURST,
    output wire [1:0]                      M_AXIMM_60_AWLOCK,
    output wire [3:0]                      M_AXIMM_60_AWCACHE,
    output wire [2:0]                      M_AXIMM_60_AWPROT,
    output wire [3:0]                      M_AXIMM_60_AWREGION,
    output wire [3:0]                      M_AXIMM_60_AWQOS,
    output wire                            M_AXIMM_60_AWVALID,
    input  wire                            M_AXIMM_60_AWREADY,
    output wire [M_AXIMM_60_DATA_WIDTH-1:0]   M_AXIMM_60_WDATA,
    output wire [M_AXIMM_60_DATA_WIDTH/8-1:0] M_AXIMM_60_WSTRB,
    output wire                            M_AXIMM_60_WLAST,
    output wire                            M_AXIMM_60_WVALID,
    input  wire                            M_AXIMM_60_WREADY,
    input  wire [1:0]                      M_AXIMM_60_BRESP,
    input  wire                            M_AXIMM_60_BVALID,
    output wire                            M_AXIMM_60_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_60_ARADDR,
    output wire [7:0]                      M_AXIMM_60_ARLEN,
    output wire [2:0]                      M_AXIMM_60_ARSIZE,
    output wire [1:0]                      M_AXIMM_60_ARBURST,
    output wire [1:0]                      M_AXIMM_60_ARLOCK,
    output wire [3:0]                      M_AXIMM_60_ARCACHE,
    output wire [2:0]                      M_AXIMM_60_ARPROT,
    output wire [3:0]                      M_AXIMM_60_ARREGION,
    output wire [3:0]                      M_AXIMM_60_ARQOS,
    output wire                            M_AXIMM_60_ARVALID,
    input  wire                            M_AXIMM_60_ARREADY,
    input  wire [M_AXIMM_60_DATA_WIDTH-1:0]   M_AXIMM_60_RDATA,
    input  wire [1:0]                      M_AXIMM_60_RRESP,
    input  wire                            M_AXIMM_60_RLAST,
    input  wire                            M_AXIMM_60_RVALID,
    output wire                            M_AXIMM_60_RREADY,
    //AXI-MM pass-through interface 61
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_61_AWADDR,
    input wire [7:0]                      AP_AXIMM_61_AWLEN,
    input wire [2:0]                      AP_AXIMM_61_AWSIZE,
    input wire [1:0]                      AP_AXIMM_61_AWBURST,
    input wire [1:0]                      AP_AXIMM_61_AWLOCK,
    input wire [3:0]                      AP_AXIMM_61_AWCACHE,
    input wire [2:0]                      AP_AXIMM_61_AWPROT,
    input wire [3:0]                      AP_AXIMM_61_AWREGION,
    input wire [3:0]                      AP_AXIMM_61_AWQOS,
    input wire                            AP_AXIMM_61_AWVALID,
    output  wire                            AP_AXIMM_61_AWREADY,
    input wire [M_AXIMM_61_DATA_WIDTH-1:0]   AP_AXIMM_61_WDATA,
    input wire [M_AXIMM_61_DATA_WIDTH/8-1:0] AP_AXIMM_61_WSTRB,
    input wire                            AP_AXIMM_61_WLAST,
    input wire                            AP_AXIMM_61_WVALID,
    output  wire                            AP_AXIMM_61_WREADY,
    output  wire [1:0]                      AP_AXIMM_61_BRESP,
    output  wire                            AP_AXIMM_61_BVALID,
    input wire                            AP_AXIMM_61_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_61_ARADDR,
    input wire [7:0]                      AP_AXIMM_61_ARLEN,
    input wire [2:0]                      AP_AXIMM_61_ARSIZE,
    input wire [1:0]                      AP_AXIMM_61_ARBURST,
    input wire [1:0]                      AP_AXIMM_61_ARLOCK,
    input wire [3:0]                      AP_AXIMM_61_ARCACHE,
    input wire [2:0]                      AP_AXIMM_61_ARPROT,
    input wire [3:0]                      AP_AXIMM_61_ARREGION,
    input wire [3:0]                      AP_AXIMM_61_ARQOS,
    input wire                            AP_AXIMM_61_ARVALID,
    output  wire                            AP_AXIMM_61_ARREADY,
    output  wire [M_AXIMM_61_DATA_WIDTH-1:0]   AP_AXIMM_61_RDATA,
    output  wire [1:0]                      AP_AXIMM_61_RRESP,
    output  wire                            AP_AXIMM_61_RLAST,
    output  wire                            AP_AXIMM_61_RVALID,
    input  wire                            AP_AXIMM_61_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_61_AWADDR,
    output wire [7:0]                      M_AXIMM_61_AWLEN,
    output wire [2:0]                      M_AXIMM_61_AWSIZE,
    output wire [1:0]                      M_AXIMM_61_AWBURST,
    output wire [1:0]                      M_AXIMM_61_AWLOCK,
    output wire [3:0]                      M_AXIMM_61_AWCACHE,
    output wire [2:0]                      M_AXIMM_61_AWPROT,
    output wire [3:0]                      M_AXIMM_61_AWREGION,
    output wire [3:0]                      M_AXIMM_61_AWQOS,
    output wire                            M_AXIMM_61_AWVALID,
    input  wire                            M_AXIMM_61_AWREADY,
    output wire [M_AXIMM_61_DATA_WIDTH-1:0]   M_AXIMM_61_WDATA,
    output wire [M_AXIMM_61_DATA_WIDTH/8-1:0] M_AXIMM_61_WSTRB,
    output wire                            M_AXIMM_61_WLAST,
    output wire                            M_AXIMM_61_WVALID,
    input  wire                            M_AXIMM_61_WREADY,
    input  wire [1:0]                      M_AXIMM_61_BRESP,
    input  wire                            M_AXIMM_61_BVALID,
    output wire                            M_AXIMM_61_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_61_ARADDR,
    output wire [7:0]                      M_AXIMM_61_ARLEN,
    output wire [2:0]                      M_AXIMM_61_ARSIZE,
    output wire [1:0]                      M_AXIMM_61_ARBURST,
    output wire [1:0]                      M_AXIMM_61_ARLOCK,
    output wire [3:0]                      M_AXIMM_61_ARCACHE,
    output wire [2:0]                      M_AXIMM_61_ARPROT,
    output wire [3:0]                      M_AXIMM_61_ARREGION,
    output wire [3:0]                      M_AXIMM_61_ARQOS,
    output wire                            M_AXIMM_61_ARVALID,
    input  wire                            M_AXIMM_61_ARREADY,
    input  wire [M_AXIMM_61_DATA_WIDTH-1:0]   M_AXIMM_61_RDATA,
    input  wire [1:0]                      M_AXIMM_61_RRESP,
    input  wire                            M_AXIMM_61_RLAST,
    input  wire                            M_AXIMM_61_RVALID,
    output wire                            M_AXIMM_61_RREADY,
    //AXI-MM pass-through interface 62
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_62_AWADDR,
    input wire [7:0]                      AP_AXIMM_62_AWLEN,
    input wire [2:0]                      AP_AXIMM_62_AWSIZE,
    input wire [1:0]                      AP_AXIMM_62_AWBURST,
    input wire [1:0]                      AP_AXIMM_62_AWLOCK,
    input wire [3:0]                      AP_AXIMM_62_AWCACHE,
    input wire [2:0]                      AP_AXIMM_62_AWPROT,
    input wire [3:0]                      AP_AXIMM_62_AWREGION,
    input wire [3:0]                      AP_AXIMM_62_AWQOS,
    input wire                            AP_AXIMM_62_AWVALID,
    output  wire                            AP_AXIMM_62_AWREADY,
    input wire [M_AXIMM_62_DATA_WIDTH-1:0]   AP_AXIMM_62_WDATA,
    input wire [M_AXIMM_62_DATA_WIDTH/8-1:0] AP_AXIMM_62_WSTRB,
    input wire                            AP_AXIMM_62_WLAST,
    input wire                            AP_AXIMM_62_WVALID,
    output  wire                            AP_AXIMM_62_WREADY,
    output  wire [1:0]                      AP_AXIMM_62_BRESP,
    output  wire                            AP_AXIMM_62_BVALID,
    input wire                            AP_AXIMM_62_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_62_ARADDR,
    input wire [7:0]                      AP_AXIMM_62_ARLEN,
    input wire [2:0]                      AP_AXIMM_62_ARSIZE,
    input wire [1:0]                      AP_AXIMM_62_ARBURST,
    input wire [1:0]                      AP_AXIMM_62_ARLOCK,
    input wire [3:0]                      AP_AXIMM_62_ARCACHE,
    input wire [2:0]                      AP_AXIMM_62_ARPROT,
    input wire [3:0]                      AP_AXIMM_62_ARREGION,
    input wire [3:0]                      AP_AXIMM_62_ARQOS,
    input wire                            AP_AXIMM_62_ARVALID,
    output  wire                            AP_AXIMM_62_ARREADY,
    output  wire [M_AXIMM_62_DATA_WIDTH-1:0]   AP_AXIMM_62_RDATA,
    output  wire [1:0]                      AP_AXIMM_62_RRESP,
    output  wire                            AP_AXIMM_62_RLAST,
    output  wire                            AP_AXIMM_62_RVALID,
    input  wire                            AP_AXIMM_62_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_62_AWADDR,
    output wire [7:0]                      M_AXIMM_62_AWLEN,
    output wire [2:0]                      M_AXIMM_62_AWSIZE,
    output wire [1:0]                      M_AXIMM_62_AWBURST,
    output wire [1:0]                      M_AXIMM_62_AWLOCK,
    output wire [3:0]                      M_AXIMM_62_AWCACHE,
    output wire [2:0]                      M_AXIMM_62_AWPROT,
    output wire [3:0]                      M_AXIMM_62_AWREGION,
    output wire [3:0]                      M_AXIMM_62_AWQOS,
    output wire                            M_AXIMM_62_AWVALID,
    input  wire                            M_AXIMM_62_AWREADY,
    output wire [M_AXIMM_62_DATA_WIDTH-1:0]   M_AXIMM_62_WDATA,
    output wire [M_AXIMM_62_DATA_WIDTH/8-1:0] M_AXIMM_62_WSTRB,
    output wire                            M_AXIMM_62_WLAST,
    output wire                            M_AXIMM_62_WVALID,
    input  wire                            M_AXIMM_62_WREADY,
    input  wire [1:0]                      M_AXIMM_62_BRESP,
    input  wire                            M_AXIMM_62_BVALID,
    output wire                            M_AXIMM_62_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_62_ARADDR,
    output wire [7:0]                      M_AXIMM_62_ARLEN,
    output wire [2:0]                      M_AXIMM_62_ARSIZE,
    output wire [1:0]                      M_AXIMM_62_ARBURST,
    output wire [1:0]                      M_AXIMM_62_ARLOCK,
    output wire [3:0]                      M_AXIMM_62_ARCACHE,
    output wire [2:0]                      M_AXIMM_62_ARPROT,
    output wire [3:0]                      M_AXIMM_62_ARREGION,
    output wire [3:0]                      M_AXIMM_62_ARQOS,
    output wire                            M_AXIMM_62_ARVALID,
    input  wire                            M_AXIMM_62_ARREADY,
    input  wire [M_AXIMM_62_DATA_WIDTH-1:0]   M_AXIMM_62_RDATA,
    input  wire [1:0]                      M_AXIMM_62_RRESP,
    input  wire                            M_AXIMM_62_RLAST,
    input  wire                            M_AXIMM_62_RVALID,
    output wire                            M_AXIMM_62_RREADY,
    //AXI-MM pass-through interface 63
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_63_AWADDR,
    input wire [7:0]                      AP_AXIMM_63_AWLEN,
    input wire [2:0]                      AP_AXIMM_63_AWSIZE,
    input wire [1:0]                      AP_AXIMM_63_AWBURST,
    input wire [1:0]                      AP_AXIMM_63_AWLOCK,
    input wire [3:0]                      AP_AXIMM_63_AWCACHE,
    input wire [2:0]                      AP_AXIMM_63_AWPROT,
    input wire [3:0]                      AP_AXIMM_63_AWREGION,
    input wire [3:0]                      AP_AXIMM_63_AWQOS,
    input wire                            AP_AXIMM_63_AWVALID,
    output  wire                            AP_AXIMM_63_AWREADY,
    input wire [M_AXIMM_63_DATA_WIDTH-1:0]   AP_AXIMM_63_WDATA,
    input wire [M_AXIMM_63_DATA_WIDTH/8-1:0] AP_AXIMM_63_WSTRB,
    input wire                            AP_AXIMM_63_WLAST,
    input wire                            AP_AXIMM_63_WVALID,
    output  wire                            AP_AXIMM_63_WREADY,
    output  wire [1:0]                      AP_AXIMM_63_BRESP,
    output  wire                            AP_AXIMM_63_BVALID,
    input wire                            AP_AXIMM_63_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_63_ARADDR,
    input wire [7:0]                      AP_AXIMM_63_ARLEN,
    input wire [2:0]                      AP_AXIMM_63_ARSIZE,
    input wire [1:0]                      AP_AXIMM_63_ARBURST,
    input wire [1:0]                      AP_AXIMM_63_ARLOCK,
    input wire [3:0]                      AP_AXIMM_63_ARCACHE,
    input wire [2:0]                      AP_AXIMM_63_ARPROT,
    input wire [3:0]                      AP_AXIMM_63_ARREGION,
    input wire [3:0]                      AP_AXIMM_63_ARQOS,
    input wire                            AP_AXIMM_63_ARVALID,
    output  wire                            AP_AXIMM_63_ARREADY,
    output  wire [M_AXIMM_63_DATA_WIDTH-1:0]   AP_AXIMM_63_RDATA,
    output  wire [1:0]                      AP_AXIMM_63_RRESP,
    output  wire                            AP_AXIMM_63_RLAST,
    output  wire                            AP_AXIMM_63_RVALID,
    input  wire                            AP_AXIMM_63_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_63_AWADDR,
    output wire [7:0]                      M_AXIMM_63_AWLEN,
    output wire [2:0]                      M_AXIMM_63_AWSIZE,
    output wire [1:0]                      M_AXIMM_63_AWBURST,
    output wire [1:0]                      M_AXIMM_63_AWLOCK,
    output wire [3:0]                      M_AXIMM_63_AWCACHE,
    output wire [2:0]                      M_AXIMM_63_AWPROT,
    output wire [3:0]                      M_AXIMM_63_AWREGION,
    output wire [3:0]                      M_AXIMM_63_AWQOS,
    output wire                            M_AXIMM_63_AWVALID,
    input  wire                            M_AXIMM_63_AWREADY,
    output wire [M_AXIMM_63_DATA_WIDTH-1:0]   M_AXIMM_63_WDATA,
    output wire [M_AXIMM_63_DATA_WIDTH/8-1:0] M_AXIMM_63_WSTRB,
    output wire                            M_AXIMM_63_WLAST,
    output wire                            M_AXIMM_63_WVALID,
    input  wire                            M_AXIMM_63_WREADY,
    input  wire [1:0]                      M_AXIMM_63_BRESP,
    input  wire                            M_AXIMM_63_BVALID,
    output wire                            M_AXIMM_63_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_63_ARADDR,
    output wire [7:0]                      M_AXIMM_63_ARLEN,
    output wire [2:0]                      M_AXIMM_63_ARSIZE,
    output wire [1:0]                      M_AXIMM_63_ARBURST,
    output wire [1:0]                      M_AXIMM_63_ARLOCK,
    output wire [3:0]                      M_AXIMM_63_ARCACHE,
    output wire [2:0]                      M_AXIMM_63_ARPROT,
    output wire [3:0]                      M_AXIMM_63_ARREGION,
    output wire [3:0]                      M_AXIMM_63_ARQOS,
    output wire                            M_AXIMM_63_ARVALID,
    input  wire                            M_AXIMM_63_ARREADY,
    input  wire [M_AXIMM_63_DATA_WIDTH-1:0]   M_AXIMM_63_RDATA,
    input  wire [1:0]                      M_AXIMM_63_RRESP,
    input  wire                            M_AXIMM_63_RLAST,
    input  wire                            M_AXIMM_63_RVALID,
    output wire                            M_AXIMM_63_RREADY,
    //AXI-MM pass-through interface 64
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_64_AWADDR,
    input wire [7:0]                      AP_AXIMM_64_AWLEN,
    input wire [2:0]                      AP_AXIMM_64_AWSIZE,
    input wire [1:0]                      AP_AXIMM_64_AWBURST,
    input wire [1:0]                      AP_AXIMM_64_AWLOCK,
    input wire [3:0]                      AP_AXIMM_64_AWCACHE,
    input wire [2:0]                      AP_AXIMM_64_AWPROT,
    input wire [3:0]                      AP_AXIMM_64_AWREGION,
    input wire [3:0]                      AP_AXIMM_64_AWQOS,
    input wire                            AP_AXIMM_64_AWVALID,
    output  wire                            AP_AXIMM_64_AWREADY,
    input wire [M_AXIMM_64_DATA_WIDTH-1:0]   AP_AXIMM_64_WDATA,
    input wire [M_AXIMM_64_DATA_WIDTH/8-1:0] AP_AXIMM_64_WSTRB,
    input wire                            AP_AXIMM_64_WLAST,
    input wire                            AP_AXIMM_64_WVALID,
    output  wire                            AP_AXIMM_64_WREADY,
    output  wire [1:0]                      AP_AXIMM_64_BRESP,
    output  wire                            AP_AXIMM_64_BVALID,
    input wire                            AP_AXIMM_64_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_64_ARADDR,
    input wire [7:0]                      AP_AXIMM_64_ARLEN,
    input wire [2:0]                      AP_AXIMM_64_ARSIZE,
    input wire [1:0]                      AP_AXIMM_64_ARBURST,
    input wire [1:0]                      AP_AXIMM_64_ARLOCK,
    input wire [3:0]                      AP_AXIMM_64_ARCACHE,
    input wire [2:0]                      AP_AXIMM_64_ARPROT,
    input wire [3:0]                      AP_AXIMM_64_ARREGION,
    input wire [3:0]                      AP_AXIMM_64_ARQOS,
    input wire                            AP_AXIMM_64_ARVALID,
    output  wire                            AP_AXIMM_64_ARREADY,
    output  wire [M_AXIMM_64_DATA_WIDTH-1:0]   AP_AXIMM_64_RDATA,
    output  wire [1:0]                      AP_AXIMM_64_RRESP,
    output  wire                            AP_AXIMM_64_RLAST,
    output  wire                            AP_AXIMM_64_RVALID,
    input  wire                            AP_AXIMM_64_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_64_AWADDR,
    output wire [7:0]                      M_AXIMM_64_AWLEN,
    output wire [2:0]                      M_AXIMM_64_AWSIZE,
    output wire [1:0]                      M_AXIMM_64_AWBURST,
    output wire [1:0]                      M_AXIMM_64_AWLOCK,
    output wire [3:0]                      M_AXIMM_64_AWCACHE,
    output wire [2:0]                      M_AXIMM_64_AWPROT,
    output wire [3:0]                      M_AXIMM_64_AWREGION,
    output wire [3:0]                      M_AXIMM_64_AWQOS,
    output wire                            M_AXIMM_64_AWVALID,
    input  wire                            M_AXIMM_64_AWREADY,
    output wire [M_AXIMM_64_DATA_WIDTH-1:0]   M_AXIMM_64_WDATA,
    output wire [M_AXIMM_64_DATA_WIDTH/8-1:0] M_AXIMM_64_WSTRB,
    output wire                            M_AXIMM_64_WLAST,
    output wire                            M_AXIMM_64_WVALID,
    input  wire                            M_AXIMM_64_WREADY,
    input  wire [1:0]                      M_AXIMM_64_BRESP,
    input  wire                            M_AXIMM_64_BVALID,
    output wire                            M_AXIMM_64_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_64_ARADDR,
    output wire [7:0]                      M_AXIMM_64_ARLEN,
    output wire [2:0]                      M_AXIMM_64_ARSIZE,
    output wire [1:0]                      M_AXIMM_64_ARBURST,
    output wire [1:0]                      M_AXIMM_64_ARLOCK,
    output wire [3:0]                      M_AXIMM_64_ARCACHE,
    output wire [2:0]                      M_AXIMM_64_ARPROT,
    output wire [3:0]                      M_AXIMM_64_ARREGION,
    output wire [3:0]                      M_AXIMM_64_ARQOS,
    output wire                            M_AXIMM_64_ARVALID,
    input  wire                            M_AXIMM_64_ARREADY,
    input  wire [M_AXIMM_64_DATA_WIDTH-1:0]   M_AXIMM_64_RDATA,
    input  wire [1:0]                      M_AXIMM_64_RRESP,
    input  wire                            M_AXIMM_64_RLAST,
    input  wire                            M_AXIMM_64_RVALID,
    output wire                            M_AXIMM_64_RREADY,
    //AXI-MM pass-through interface 65
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_65_AWADDR,
    input wire [7:0]                      AP_AXIMM_65_AWLEN,
    input wire [2:0]                      AP_AXIMM_65_AWSIZE,
    input wire [1:0]                      AP_AXIMM_65_AWBURST,
    input wire [1:0]                      AP_AXIMM_65_AWLOCK,
    input wire [3:0]                      AP_AXIMM_65_AWCACHE,
    input wire [2:0]                      AP_AXIMM_65_AWPROT,
    input wire [3:0]                      AP_AXIMM_65_AWREGION,
    input wire [3:0]                      AP_AXIMM_65_AWQOS,
    input wire                            AP_AXIMM_65_AWVALID,
    output  wire                            AP_AXIMM_65_AWREADY,
    input wire [M_AXIMM_65_DATA_WIDTH-1:0]   AP_AXIMM_65_WDATA,
    input wire [M_AXIMM_65_DATA_WIDTH/8-1:0] AP_AXIMM_65_WSTRB,
    input wire                            AP_AXIMM_65_WLAST,
    input wire                            AP_AXIMM_65_WVALID,
    output  wire                            AP_AXIMM_65_WREADY,
    output  wire [1:0]                      AP_AXIMM_65_BRESP,
    output  wire                            AP_AXIMM_65_BVALID,
    input wire                            AP_AXIMM_65_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_65_ARADDR,
    input wire [7:0]                      AP_AXIMM_65_ARLEN,
    input wire [2:0]                      AP_AXIMM_65_ARSIZE,
    input wire [1:0]                      AP_AXIMM_65_ARBURST,
    input wire [1:0]                      AP_AXIMM_65_ARLOCK,
    input wire [3:0]                      AP_AXIMM_65_ARCACHE,
    input wire [2:0]                      AP_AXIMM_65_ARPROT,
    input wire [3:0]                      AP_AXIMM_65_ARREGION,
    input wire [3:0]                      AP_AXIMM_65_ARQOS,
    input wire                            AP_AXIMM_65_ARVALID,
    output  wire                            AP_AXIMM_65_ARREADY,
    output  wire [M_AXIMM_65_DATA_WIDTH-1:0]   AP_AXIMM_65_RDATA,
    output  wire [1:0]                      AP_AXIMM_65_RRESP,
    output  wire                            AP_AXIMM_65_RLAST,
    output  wire                            AP_AXIMM_65_RVALID,
    input  wire                            AP_AXIMM_65_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_65_AWADDR,
    output wire [7:0]                      M_AXIMM_65_AWLEN,
    output wire [2:0]                      M_AXIMM_65_AWSIZE,
    output wire [1:0]                      M_AXIMM_65_AWBURST,
    output wire [1:0]                      M_AXIMM_65_AWLOCK,
    output wire [3:0]                      M_AXIMM_65_AWCACHE,
    output wire [2:0]                      M_AXIMM_65_AWPROT,
    output wire [3:0]                      M_AXIMM_65_AWREGION,
    output wire [3:0]                      M_AXIMM_65_AWQOS,
    output wire                            M_AXIMM_65_AWVALID,
    input  wire                            M_AXIMM_65_AWREADY,
    output wire [M_AXIMM_65_DATA_WIDTH-1:0]   M_AXIMM_65_WDATA,
    output wire [M_AXIMM_65_DATA_WIDTH/8-1:0] M_AXIMM_65_WSTRB,
    output wire                            M_AXIMM_65_WLAST,
    output wire                            M_AXIMM_65_WVALID,
    input  wire                            M_AXIMM_65_WREADY,
    input  wire [1:0]                      M_AXIMM_65_BRESP,
    input  wire                            M_AXIMM_65_BVALID,
    output wire                            M_AXIMM_65_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_65_ARADDR,
    output wire [7:0]                      M_AXIMM_65_ARLEN,
    output wire [2:0]                      M_AXIMM_65_ARSIZE,
    output wire [1:0]                      M_AXIMM_65_ARBURST,
    output wire [1:0]                      M_AXIMM_65_ARLOCK,
    output wire [3:0]                      M_AXIMM_65_ARCACHE,
    output wire [2:0]                      M_AXIMM_65_ARPROT,
    output wire [3:0]                      M_AXIMM_65_ARREGION,
    output wire [3:0]                      M_AXIMM_65_ARQOS,
    output wire                            M_AXIMM_65_ARVALID,
    input  wire                            M_AXIMM_65_ARREADY,
    input  wire [M_AXIMM_65_DATA_WIDTH-1:0]   M_AXIMM_65_RDATA,
    input  wire [1:0]                      M_AXIMM_65_RRESP,
    input  wire                            M_AXIMM_65_RLAST,
    input  wire                            M_AXIMM_65_RVALID,
    output wire                            M_AXIMM_65_RREADY,
    //AXI-MM pass-through interface 66
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_66_AWADDR,
    input wire [7:0]                      AP_AXIMM_66_AWLEN,
    input wire [2:0]                      AP_AXIMM_66_AWSIZE,
    input wire [1:0]                      AP_AXIMM_66_AWBURST,
    input wire [1:0]                      AP_AXIMM_66_AWLOCK,
    input wire [3:0]                      AP_AXIMM_66_AWCACHE,
    input wire [2:0]                      AP_AXIMM_66_AWPROT,
    input wire [3:0]                      AP_AXIMM_66_AWREGION,
    input wire [3:0]                      AP_AXIMM_66_AWQOS,
    input wire                            AP_AXIMM_66_AWVALID,
    output  wire                            AP_AXIMM_66_AWREADY,
    input wire [M_AXIMM_66_DATA_WIDTH-1:0]   AP_AXIMM_66_WDATA,
    input wire [M_AXIMM_66_DATA_WIDTH/8-1:0] AP_AXIMM_66_WSTRB,
    input wire                            AP_AXIMM_66_WLAST,
    input wire                            AP_AXIMM_66_WVALID,
    output  wire                            AP_AXIMM_66_WREADY,
    output  wire [1:0]                      AP_AXIMM_66_BRESP,
    output  wire                            AP_AXIMM_66_BVALID,
    input wire                            AP_AXIMM_66_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_66_ARADDR,
    input wire [7:0]                      AP_AXIMM_66_ARLEN,
    input wire [2:0]                      AP_AXIMM_66_ARSIZE,
    input wire [1:0]                      AP_AXIMM_66_ARBURST,
    input wire [1:0]                      AP_AXIMM_66_ARLOCK,
    input wire [3:0]                      AP_AXIMM_66_ARCACHE,
    input wire [2:0]                      AP_AXIMM_66_ARPROT,
    input wire [3:0]                      AP_AXIMM_66_ARREGION,
    input wire [3:0]                      AP_AXIMM_66_ARQOS,
    input wire                            AP_AXIMM_66_ARVALID,
    output  wire                            AP_AXIMM_66_ARREADY,
    output  wire [M_AXIMM_66_DATA_WIDTH-1:0]   AP_AXIMM_66_RDATA,
    output  wire [1:0]                      AP_AXIMM_66_RRESP,
    output  wire                            AP_AXIMM_66_RLAST,
    output  wire                            AP_AXIMM_66_RVALID,
    input  wire                            AP_AXIMM_66_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_66_AWADDR,
    output wire [7:0]                      M_AXIMM_66_AWLEN,
    output wire [2:0]                      M_AXIMM_66_AWSIZE,
    output wire [1:0]                      M_AXIMM_66_AWBURST,
    output wire [1:0]                      M_AXIMM_66_AWLOCK,
    output wire [3:0]                      M_AXIMM_66_AWCACHE,
    output wire [2:0]                      M_AXIMM_66_AWPROT,
    output wire [3:0]                      M_AXIMM_66_AWREGION,
    output wire [3:0]                      M_AXIMM_66_AWQOS,
    output wire                            M_AXIMM_66_AWVALID,
    input  wire                            M_AXIMM_66_AWREADY,
    output wire [M_AXIMM_66_DATA_WIDTH-1:0]   M_AXIMM_66_WDATA,
    output wire [M_AXIMM_66_DATA_WIDTH/8-1:0] M_AXIMM_66_WSTRB,
    output wire                            M_AXIMM_66_WLAST,
    output wire                            M_AXIMM_66_WVALID,
    input  wire                            M_AXIMM_66_WREADY,
    input  wire [1:0]                      M_AXIMM_66_BRESP,
    input  wire                            M_AXIMM_66_BVALID,
    output wire                            M_AXIMM_66_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_66_ARADDR,
    output wire [7:0]                      M_AXIMM_66_ARLEN,
    output wire [2:0]                      M_AXIMM_66_ARSIZE,
    output wire [1:0]                      M_AXIMM_66_ARBURST,
    output wire [1:0]                      M_AXIMM_66_ARLOCK,
    output wire [3:0]                      M_AXIMM_66_ARCACHE,
    output wire [2:0]                      M_AXIMM_66_ARPROT,
    output wire [3:0]                      M_AXIMM_66_ARREGION,
    output wire [3:0]                      M_AXIMM_66_ARQOS,
    output wire                            M_AXIMM_66_ARVALID,
    input  wire                            M_AXIMM_66_ARREADY,
    input  wire [M_AXIMM_66_DATA_WIDTH-1:0]   M_AXIMM_66_RDATA,
    input  wire [1:0]                      M_AXIMM_66_RRESP,
    input  wire                            M_AXIMM_66_RLAST,
    input  wire                            M_AXIMM_66_RVALID,
    output wire                            M_AXIMM_66_RREADY,
    //AXI-MM pass-through interface 67
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_67_AWADDR,
    input wire [7:0]                      AP_AXIMM_67_AWLEN,
    input wire [2:0]                      AP_AXIMM_67_AWSIZE,
    input wire [1:0]                      AP_AXIMM_67_AWBURST,
    input wire [1:0]                      AP_AXIMM_67_AWLOCK,
    input wire [3:0]                      AP_AXIMM_67_AWCACHE,
    input wire [2:0]                      AP_AXIMM_67_AWPROT,
    input wire [3:0]                      AP_AXIMM_67_AWREGION,
    input wire [3:0]                      AP_AXIMM_67_AWQOS,
    input wire                            AP_AXIMM_67_AWVALID,
    output  wire                            AP_AXIMM_67_AWREADY,
    input wire [M_AXIMM_67_DATA_WIDTH-1:0]   AP_AXIMM_67_WDATA,
    input wire [M_AXIMM_67_DATA_WIDTH/8-1:0] AP_AXIMM_67_WSTRB,
    input wire                            AP_AXIMM_67_WLAST,
    input wire                            AP_AXIMM_67_WVALID,
    output  wire                            AP_AXIMM_67_WREADY,
    output  wire [1:0]                      AP_AXIMM_67_BRESP,
    output  wire                            AP_AXIMM_67_BVALID,
    input wire                            AP_AXIMM_67_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_67_ARADDR,
    input wire [7:0]                      AP_AXIMM_67_ARLEN,
    input wire [2:0]                      AP_AXIMM_67_ARSIZE,
    input wire [1:0]                      AP_AXIMM_67_ARBURST,
    input wire [1:0]                      AP_AXIMM_67_ARLOCK,
    input wire [3:0]                      AP_AXIMM_67_ARCACHE,
    input wire [2:0]                      AP_AXIMM_67_ARPROT,
    input wire [3:0]                      AP_AXIMM_67_ARREGION,
    input wire [3:0]                      AP_AXIMM_67_ARQOS,
    input wire                            AP_AXIMM_67_ARVALID,
    output  wire                            AP_AXIMM_67_ARREADY,
    output  wire [M_AXIMM_67_DATA_WIDTH-1:0]   AP_AXIMM_67_RDATA,
    output  wire [1:0]                      AP_AXIMM_67_RRESP,
    output  wire                            AP_AXIMM_67_RLAST,
    output  wire                            AP_AXIMM_67_RVALID,
    input  wire                            AP_AXIMM_67_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_67_AWADDR,
    output wire [7:0]                      M_AXIMM_67_AWLEN,
    output wire [2:0]                      M_AXIMM_67_AWSIZE,
    output wire [1:0]                      M_AXIMM_67_AWBURST,
    output wire [1:0]                      M_AXIMM_67_AWLOCK,
    output wire [3:0]                      M_AXIMM_67_AWCACHE,
    output wire [2:0]                      M_AXIMM_67_AWPROT,
    output wire [3:0]                      M_AXIMM_67_AWREGION,
    output wire [3:0]                      M_AXIMM_67_AWQOS,
    output wire                            M_AXIMM_67_AWVALID,
    input  wire                            M_AXIMM_67_AWREADY,
    output wire [M_AXIMM_67_DATA_WIDTH-1:0]   M_AXIMM_67_WDATA,
    output wire [M_AXIMM_67_DATA_WIDTH/8-1:0] M_AXIMM_67_WSTRB,
    output wire                            M_AXIMM_67_WLAST,
    output wire                            M_AXIMM_67_WVALID,
    input  wire                            M_AXIMM_67_WREADY,
    input  wire [1:0]                      M_AXIMM_67_BRESP,
    input  wire                            M_AXIMM_67_BVALID,
    output wire                            M_AXIMM_67_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_67_ARADDR,
    output wire [7:0]                      M_AXIMM_67_ARLEN,
    output wire [2:0]                      M_AXIMM_67_ARSIZE,
    output wire [1:0]                      M_AXIMM_67_ARBURST,
    output wire [1:0]                      M_AXIMM_67_ARLOCK,
    output wire [3:0]                      M_AXIMM_67_ARCACHE,
    output wire [2:0]                      M_AXIMM_67_ARPROT,
    output wire [3:0]                      M_AXIMM_67_ARREGION,
    output wire [3:0]                      M_AXIMM_67_ARQOS,
    output wire                            M_AXIMM_67_ARVALID,
    input  wire                            M_AXIMM_67_ARREADY,
    input  wire [M_AXIMM_67_DATA_WIDTH-1:0]   M_AXIMM_67_RDATA,
    input  wire [1:0]                      M_AXIMM_67_RRESP,
    input  wire                            M_AXIMM_67_RLAST,
    input  wire                            M_AXIMM_67_RVALID,
    output wire                            M_AXIMM_67_RREADY,
    //AXI-MM pass-through interface 68
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_68_AWADDR,
    input wire [7:0]                      AP_AXIMM_68_AWLEN,
    input wire [2:0]                      AP_AXIMM_68_AWSIZE,
    input wire [1:0]                      AP_AXIMM_68_AWBURST,
    input wire [1:0]                      AP_AXIMM_68_AWLOCK,
    input wire [3:0]                      AP_AXIMM_68_AWCACHE,
    input wire [2:0]                      AP_AXIMM_68_AWPROT,
    input wire [3:0]                      AP_AXIMM_68_AWREGION,
    input wire [3:0]                      AP_AXIMM_68_AWQOS,
    input wire                            AP_AXIMM_68_AWVALID,
    output  wire                            AP_AXIMM_68_AWREADY,
    input wire [M_AXIMM_68_DATA_WIDTH-1:0]   AP_AXIMM_68_WDATA,
    input wire [M_AXIMM_68_DATA_WIDTH/8-1:0] AP_AXIMM_68_WSTRB,
    input wire                            AP_AXIMM_68_WLAST,
    input wire                            AP_AXIMM_68_WVALID,
    output  wire                            AP_AXIMM_68_WREADY,
    output  wire [1:0]                      AP_AXIMM_68_BRESP,
    output  wire                            AP_AXIMM_68_BVALID,
    input wire                            AP_AXIMM_68_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_68_ARADDR,
    input wire [7:0]                      AP_AXIMM_68_ARLEN,
    input wire [2:0]                      AP_AXIMM_68_ARSIZE,
    input wire [1:0]                      AP_AXIMM_68_ARBURST,
    input wire [1:0]                      AP_AXIMM_68_ARLOCK,
    input wire [3:0]                      AP_AXIMM_68_ARCACHE,
    input wire [2:0]                      AP_AXIMM_68_ARPROT,
    input wire [3:0]                      AP_AXIMM_68_ARREGION,
    input wire [3:0]                      AP_AXIMM_68_ARQOS,
    input wire                            AP_AXIMM_68_ARVALID,
    output  wire                            AP_AXIMM_68_ARREADY,
    output  wire [M_AXIMM_68_DATA_WIDTH-1:0]   AP_AXIMM_68_RDATA,
    output  wire [1:0]                      AP_AXIMM_68_RRESP,
    output  wire                            AP_AXIMM_68_RLAST,
    output  wire                            AP_AXIMM_68_RVALID,
    input  wire                            AP_AXIMM_68_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_68_AWADDR,
    output wire [7:0]                      M_AXIMM_68_AWLEN,
    output wire [2:0]                      M_AXIMM_68_AWSIZE,
    output wire [1:0]                      M_AXIMM_68_AWBURST,
    output wire [1:0]                      M_AXIMM_68_AWLOCK,
    output wire [3:0]                      M_AXIMM_68_AWCACHE,
    output wire [2:0]                      M_AXIMM_68_AWPROT,
    output wire [3:0]                      M_AXIMM_68_AWREGION,
    output wire [3:0]                      M_AXIMM_68_AWQOS,
    output wire                            M_AXIMM_68_AWVALID,
    input  wire                            M_AXIMM_68_AWREADY,
    output wire [M_AXIMM_68_DATA_WIDTH-1:0]   M_AXIMM_68_WDATA,
    output wire [M_AXIMM_68_DATA_WIDTH/8-1:0] M_AXIMM_68_WSTRB,
    output wire                            M_AXIMM_68_WLAST,
    output wire                            M_AXIMM_68_WVALID,
    input  wire                            M_AXIMM_68_WREADY,
    input  wire [1:0]                      M_AXIMM_68_BRESP,
    input  wire                            M_AXIMM_68_BVALID,
    output wire                            M_AXIMM_68_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_68_ARADDR,
    output wire [7:0]                      M_AXIMM_68_ARLEN,
    output wire [2:0]                      M_AXIMM_68_ARSIZE,
    output wire [1:0]                      M_AXIMM_68_ARBURST,
    output wire [1:0]                      M_AXIMM_68_ARLOCK,
    output wire [3:0]                      M_AXIMM_68_ARCACHE,
    output wire [2:0]                      M_AXIMM_68_ARPROT,
    output wire [3:0]                      M_AXIMM_68_ARREGION,
    output wire [3:0]                      M_AXIMM_68_ARQOS,
    output wire                            M_AXIMM_68_ARVALID,
    input  wire                            M_AXIMM_68_ARREADY,
    input  wire [M_AXIMM_68_DATA_WIDTH-1:0]   M_AXIMM_68_RDATA,
    input  wire [1:0]                      M_AXIMM_68_RRESP,
    input  wire                            M_AXIMM_68_RLAST,
    input  wire                            M_AXIMM_68_RVALID,
    output wire                            M_AXIMM_68_RREADY,
    //AXI-MM pass-through interface 69
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_69_AWADDR,
    input wire [7:0]                      AP_AXIMM_69_AWLEN,
    input wire [2:0]                      AP_AXIMM_69_AWSIZE,
    input wire [1:0]                      AP_AXIMM_69_AWBURST,
    input wire [1:0]                      AP_AXIMM_69_AWLOCK,
    input wire [3:0]                      AP_AXIMM_69_AWCACHE,
    input wire [2:0]                      AP_AXIMM_69_AWPROT,
    input wire [3:0]                      AP_AXIMM_69_AWREGION,
    input wire [3:0]                      AP_AXIMM_69_AWQOS,
    input wire                            AP_AXIMM_69_AWVALID,
    output  wire                            AP_AXIMM_69_AWREADY,
    input wire [M_AXIMM_69_DATA_WIDTH-1:0]   AP_AXIMM_69_WDATA,
    input wire [M_AXIMM_69_DATA_WIDTH/8-1:0] AP_AXIMM_69_WSTRB,
    input wire                            AP_AXIMM_69_WLAST,
    input wire                            AP_AXIMM_69_WVALID,
    output  wire                            AP_AXIMM_69_WREADY,
    output  wire [1:0]                      AP_AXIMM_69_BRESP,
    output  wire                            AP_AXIMM_69_BVALID,
    input wire                            AP_AXIMM_69_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_69_ARADDR,
    input wire [7:0]                      AP_AXIMM_69_ARLEN,
    input wire [2:0]                      AP_AXIMM_69_ARSIZE,
    input wire [1:0]                      AP_AXIMM_69_ARBURST,
    input wire [1:0]                      AP_AXIMM_69_ARLOCK,
    input wire [3:0]                      AP_AXIMM_69_ARCACHE,
    input wire [2:0]                      AP_AXIMM_69_ARPROT,
    input wire [3:0]                      AP_AXIMM_69_ARREGION,
    input wire [3:0]                      AP_AXIMM_69_ARQOS,
    input wire                            AP_AXIMM_69_ARVALID,
    output  wire                            AP_AXIMM_69_ARREADY,
    output  wire [M_AXIMM_69_DATA_WIDTH-1:0]   AP_AXIMM_69_RDATA,
    output  wire [1:0]                      AP_AXIMM_69_RRESP,
    output  wire                            AP_AXIMM_69_RLAST,
    output  wire                            AP_AXIMM_69_RVALID,
    input  wire                            AP_AXIMM_69_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_69_AWADDR,
    output wire [7:0]                      M_AXIMM_69_AWLEN,
    output wire [2:0]                      M_AXIMM_69_AWSIZE,
    output wire [1:0]                      M_AXIMM_69_AWBURST,
    output wire [1:0]                      M_AXIMM_69_AWLOCK,
    output wire [3:0]                      M_AXIMM_69_AWCACHE,
    output wire [2:0]                      M_AXIMM_69_AWPROT,
    output wire [3:0]                      M_AXIMM_69_AWREGION,
    output wire [3:0]                      M_AXIMM_69_AWQOS,
    output wire                            M_AXIMM_69_AWVALID,
    input  wire                            M_AXIMM_69_AWREADY,
    output wire [M_AXIMM_69_DATA_WIDTH-1:0]   M_AXIMM_69_WDATA,
    output wire [M_AXIMM_69_DATA_WIDTH/8-1:0] M_AXIMM_69_WSTRB,
    output wire                            M_AXIMM_69_WLAST,
    output wire                            M_AXIMM_69_WVALID,
    input  wire                            M_AXIMM_69_WREADY,
    input  wire [1:0]                      M_AXIMM_69_BRESP,
    input  wire                            M_AXIMM_69_BVALID,
    output wire                            M_AXIMM_69_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_69_ARADDR,
    output wire [7:0]                      M_AXIMM_69_ARLEN,
    output wire [2:0]                      M_AXIMM_69_ARSIZE,
    output wire [1:0]                      M_AXIMM_69_ARBURST,
    output wire [1:0]                      M_AXIMM_69_ARLOCK,
    output wire [3:0]                      M_AXIMM_69_ARCACHE,
    output wire [2:0]                      M_AXIMM_69_ARPROT,
    output wire [3:0]                      M_AXIMM_69_ARREGION,
    output wire [3:0]                      M_AXIMM_69_ARQOS,
    output wire                            M_AXIMM_69_ARVALID,
    input  wire                            M_AXIMM_69_ARREADY,
    input  wire [M_AXIMM_69_DATA_WIDTH-1:0]   M_AXIMM_69_RDATA,
    input  wire [1:0]                      M_AXIMM_69_RRESP,
    input  wire                            M_AXIMM_69_RLAST,
    input  wire                            M_AXIMM_69_RVALID,
    output wire                            M_AXIMM_69_RREADY,
    //AXI-MM pass-through interface 70
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_70_AWADDR,
    input wire [7:0]                      AP_AXIMM_70_AWLEN,
    input wire [2:0]                      AP_AXIMM_70_AWSIZE,
    input wire [1:0]                      AP_AXIMM_70_AWBURST,
    input wire [1:0]                      AP_AXIMM_70_AWLOCK,
    input wire [3:0]                      AP_AXIMM_70_AWCACHE,
    input wire [2:0]                      AP_AXIMM_70_AWPROT,
    input wire [3:0]                      AP_AXIMM_70_AWREGION,
    input wire [3:0]                      AP_AXIMM_70_AWQOS,
    input wire                            AP_AXIMM_70_AWVALID,
    output  wire                            AP_AXIMM_70_AWREADY,
    input wire [M_AXIMM_70_DATA_WIDTH-1:0]   AP_AXIMM_70_WDATA,
    input wire [M_AXIMM_70_DATA_WIDTH/8-1:0] AP_AXIMM_70_WSTRB,
    input wire                            AP_AXIMM_70_WLAST,
    input wire                            AP_AXIMM_70_WVALID,
    output  wire                            AP_AXIMM_70_WREADY,
    output  wire [1:0]                      AP_AXIMM_70_BRESP,
    output  wire                            AP_AXIMM_70_BVALID,
    input wire                            AP_AXIMM_70_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_70_ARADDR,
    input wire [7:0]                      AP_AXIMM_70_ARLEN,
    input wire [2:0]                      AP_AXIMM_70_ARSIZE,
    input wire [1:0]                      AP_AXIMM_70_ARBURST,
    input wire [1:0]                      AP_AXIMM_70_ARLOCK,
    input wire [3:0]                      AP_AXIMM_70_ARCACHE,
    input wire [2:0]                      AP_AXIMM_70_ARPROT,
    input wire [3:0]                      AP_AXIMM_70_ARREGION,
    input wire [3:0]                      AP_AXIMM_70_ARQOS,
    input wire                            AP_AXIMM_70_ARVALID,
    output  wire                            AP_AXIMM_70_ARREADY,
    output  wire [M_AXIMM_70_DATA_WIDTH-1:0]   AP_AXIMM_70_RDATA,
    output  wire [1:0]                      AP_AXIMM_70_RRESP,
    output  wire                            AP_AXIMM_70_RLAST,
    output  wire                            AP_AXIMM_70_RVALID,
    input  wire                            AP_AXIMM_70_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_70_AWADDR,
    output wire [7:0]                      M_AXIMM_70_AWLEN,
    output wire [2:0]                      M_AXIMM_70_AWSIZE,
    output wire [1:0]                      M_AXIMM_70_AWBURST,
    output wire [1:0]                      M_AXIMM_70_AWLOCK,
    output wire [3:0]                      M_AXIMM_70_AWCACHE,
    output wire [2:0]                      M_AXIMM_70_AWPROT,
    output wire [3:0]                      M_AXIMM_70_AWREGION,
    output wire [3:0]                      M_AXIMM_70_AWQOS,
    output wire                            M_AXIMM_70_AWVALID,
    input  wire                            M_AXIMM_70_AWREADY,
    output wire [M_AXIMM_70_DATA_WIDTH-1:0]   M_AXIMM_70_WDATA,
    output wire [M_AXIMM_70_DATA_WIDTH/8-1:0] M_AXIMM_70_WSTRB,
    output wire                            M_AXIMM_70_WLAST,
    output wire                            M_AXIMM_70_WVALID,
    input  wire                            M_AXIMM_70_WREADY,
    input  wire [1:0]                      M_AXIMM_70_BRESP,
    input  wire                            M_AXIMM_70_BVALID,
    output wire                            M_AXIMM_70_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_70_ARADDR,
    output wire [7:0]                      M_AXIMM_70_ARLEN,
    output wire [2:0]                      M_AXIMM_70_ARSIZE,
    output wire [1:0]                      M_AXIMM_70_ARBURST,
    output wire [1:0]                      M_AXIMM_70_ARLOCK,
    output wire [3:0]                      M_AXIMM_70_ARCACHE,
    output wire [2:0]                      M_AXIMM_70_ARPROT,
    output wire [3:0]                      M_AXIMM_70_ARREGION,
    output wire [3:0]                      M_AXIMM_70_ARQOS,
    output wire                            M_AXIMM_70_ARVALID,
    input  wire                            M_AXIMM_70_ARREADY,
    input  wire [M_AXIMM_70_DATA_WIDTH-1:0]   M_AXIMM_70_RDATA,
    input  wire [1:0]                      M_AXIMM_70_RRESP,
    input  wire                            M_AXIMM_70_RLAST,
    input  wire                            M_AXIMM_70_RVALID,
    output wire                            M_AXIMM_70_RREADY,
    //AXI-MM pass-through interface 71
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_71_AWADDR,
    input wire [7:0]                      AP_AXIMM_71_AWLEN,
    input wire [2:0]                      AP_AXIMM_71_AWSIZE,
    input wire [1:0]                      AP_AXIMM_71_AWBURST,
    input wire [1:0]                      AP_AXIMM_71_AWLOCK,
    input wire [3:0]                      AP_AXIMM_71_AWCACHE,
    input wire [2:0]                      AP_AXIMM_71_AWPROT,
    input wire [3:0]                      AP_AXIMM_71_AWREGION,
    input wire [3:0]                      AP_AXIMM_71_AWQOS,
    input wire                            AP_AXIMM_71_AWVALID,
    output  wire                            AP_AXIMM_71_AWREADY,
    input wire [M_AXIMM_71_DATA_WIDTH-1:0]   AP_AXIMM_71_WDATA,
    input wire [M_AXIMM_71_DATA_WIDTH/8-1:0] AP_AXIMM_71_WSTRB,
    input wire                            AP_AXIMM_71_WLAST,
    input wire                            AP_AXIMM_71_WVALID,
    output  wire                            AP_AXIMM_71_WREADY,
    output  wire [1:0]                      AP_AXIMM_71_BRESP,
    output  wire                            AP_AXIMM_71_BVALID,
    input wire                            AP_AXIMM_71_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_71_ARADDR,
    input wire [7:0]                      AP_AXIMM_71_ARLEN,
    input wire [2:0]                      AP_AXIMM_71_ARSIZE,
    input wire [1:0]                      AP_AXIMM_71_ARBURST,
    input wire [1:0]                      AP_AXIMM_71_ARLOCK,
    input wire [3:0]                      AP_AXIMM_71_ARCACHE,
    input wire [2:0]                      AP_AXIMM_71_ARPROT,
    input wire [3:0]                      AP_AXIMM_71_ARREGION,
    input wire [3:0]                      AP_AXIMM_71_ARQOS,
    input wire                            AP_AXIMM_71_ARVALID,
    output  wire                            AP_AXIMM_71_ARREADY,
    output  wire [M_AXIMM_71_DATA_WIDTH-1:0]   AP_AXIMM_71_RDATA,
    output  wire [1:0]                      AP_AXIMM_71_RRESP,
    output  wire                            AP_AXIMM_71_RLAST,
    output  wire                            AP_AXIMM_71_RVALID,
    input  wire                            AP_AXIMM_71_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_71_AWADDR,
    output wire [7:0]                      M_AXIMM_71_AWLEN,
    output wire [2:0]                      M_AXIMM_71_AWSIZE,
    output wire [1:0]                      M_AXIMM_71_AWBURST,
    output wire [1:0]                      M_AXIMM_71_AWLOCK,
    output wire [3:0]                      M_AXIMM_71_AWCACHE,
    output wire [2:0]                      M_AXIMM_71_AWPROT,
    output wire [3:0]                      M_AXIMM_71_AWREGION,
    output wire [3:0]                      M_AXIMM_71_AWQOS,
    output wire                            M_AXIMM_71_AWVALID,
    input  wire                            M_AXIMM_71_AWREADY,
    output wire [M_AXIMM_71_DATA_WIDTH-1:0]   M_AXIMM_71_WDATA,
    output wire [M_AXIMM_71_DATA_WIDTH/8-1:0] M_AXIMM_71_WSTRB,
    output wire                            M_AXIMM_71_WLAST,
    output wire                            M_AXIMM_71_WVALID,
    input  wire                            M_AXIMM_71_WREADY,
    input  wire [1:0]                      M_AXIMM_71_BRESP,
    input  wire                            M_AXIMM_71_BVALID,
    output wire                            M_AXIMM_71_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_71_ARADDR,
    output wire [7:0]                      M_AXIMM_71_ARLEN,
    output wire [2:0]                      M_AXIMM_71_ARSIZE,
    output wire [1:0]                      M_AXIMM_71_ARBURST,
    output wire [1:0]                      M_AXIMM_71_ARLOCK,
    output wire [3:0]                      M_AXIMM_71_ARCACHE,
    output wire [2:0]                      M_AXIMM_71_ARPROT,
    output wire [3:0]                      M_AXIMM_71_ARREGION,
    output wire [3:0]                      M_AXIMM_71_ARQOS,
    output wire                            M_AXIMM_71_ARVALID,
    input  wire                            M_AXIMM_71_ARREADY,
    input  wire [M_AXIMM_71_DATA_WIDTH-1:0]   M_AXIMM_71_RDATA,
    input  wire [1:0]                      M_AXIMM_71_RRESP,
    input  wire                            M_AXIMM_71_RLAST,
    input  wire                            M_AXIMM_71_RVALID,
    output wire                            M_AXIMM_71_RREADY,
    //AXI-MM pass-through interface 72
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_72_AWADDR,
    input wire [7:0]                      AP_AXIMM_72_AWLEN,
    input wire [2:0]                      AP_AXIMM_72_AWSIZE,
    input wire [1:0]                      AP_AXIMM_72_AWBURST,
    input wire [1:0]                      AP_AXIMM_72_AWLOCK,
    input wire [3:0]                      AP_AXIMM_72_AWCACHE,
    input wire [2:0]                      AP_AXIMM_72_AWPROT,
    input wire [3:0]                      AP_AXIMM_72_AWREGION,
    input wire [3:0]                      AP_AXIMM_72_AWQOS,
    input wire                            AP_AXIMM_72_AWVALID,
    output  wire                            AP_AXIMM_72_AWREADY,
    input wire [M_AXIMM_72_DATA_WIDTH-1:0]   AP_AXIMM_72_WDATA,
    input wire [M_AXIMM_72_DATA_WIDTH/8-1:0] AP_AXIMM_72_WSTRB,
    input wire                            AP_AXIMM_72_WLAST,
    input wire                            AP_AXIMM_72_WVALID,
    output  wire                            AP_AXIMM_72_WREADY,
    output  wire [1:0]                      AP_AXIMM_72_BRESP,
    output  wire                            AP_AXIMM_72_BVALID,
    input wire                            AP_AXIMM_72_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_72_ARADDR,
    input wire [7:0]                      AP_AXIMM_72_ARLEN,
    input wire [2:0]                      AP_AXIMM_72_ARSIZE,
    input wire [1:0]                      AP_AXIMM_72_ARBURST,
    input wire [1:0]                      AP_AXIMM_72_ARLOCK,
    input wire [3:0]                      AP_AXIMM_72_ARCACHE,
    input wire [2:0]                      AP_AXIMM_72_ARPROT,
    input wire [3:0]                      AP_AXIMM_72_ARREGION,
    input wire [3:0]                      AP_AXIMM_72_ARQOS,
    input wire                            AP_AXIMM_72_ARVALID,
    output  wire                            AP_AXIMM_72_ARREADY,
    output  wire [M_AXIMM_72_DATA_WIDTH-1:0]   AP_AXIMM_72_RDATA,
    output  wire [1:0]                      AP_AXIMM_72_RRESP,
    output  wire                            AP_AXIMM_72_RLAST,
    output  wire                            AP_AXIMM_72_RVALID,
    input  wire                            AP_AXIMM_72_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_72_AWADDR,
    output wire [7:0]                      M_AXIMM_72_AWLEN,
    output wire [2:0]                      M_AXIMM_72_AWSIZE,
    output wire [1:0]                      M_AXIMM_72_AWBURST,
    output wire [1:0]                      M_AXIMM_72_AWLOCK,
    output wire [3:0]                      M_AXIMM_72_AWCACHE,
    output wire [2:0]                      M_AXIMM_72_AWPROT,
    output wire [3:0]                      M_AXIMM_72_AWREGION,
    output wire [3:0]                      M_AXIMM_72_AWQOS,
    output wire                            M_AXIMM_72_AWVALID,
    input  wire                            M_AXIMM_72_AWREADY,
    output wire [M_AXIMM_72_DATA_WIDTH-1:0]   M_AXIMM_72_WDATA,
    output wire [M_AXIMM_72_DATA_WIDTH/8-1:0] M_AXIMM_72_WSTRB,
    output wire                            M_AXIMM_72_WLAST,
    output wire                            M_AXIMM_72_WVALID,
    input  wire                            M_AXIMM_72_WREADY,
    input  wire [1:0]                      M_AXIMM_72_BRESP,
    input  wire                            M_AXIMM_72_BVALID,
    output wire                            M_AXIMM_72_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_72_ARADDR,
    output wire [7:0]                      M_AXIMM_72_ARLEN,
    output wire [2:0]                      M_AXIMM_72_ARSIZE,
    output wire [1:0]                      M_AXIMM_72_ARBURST,
    output wire [1:0]                      M_AXIMM_72_ARLOCK,
    output wire [3:0]                      M_AXIMM_72_ARCACHE,
    output wire [2:0]                      M_AXIMM_72_ARPROT,
    output wire [3:0]                      M_AXIMM_72_ARREGION,
    output wire [3:0]                      M_AXIMM_72_ARQOS,
    output wire                            M_AXIMM_72_ARVALID,
    input  wire                            M_AXIMM_72_ARREADY,
    input  wire [M_AXIMM_72_DATA_WIDTH-1:0]   M_AXIMM_72_RDATA,
    input  wire [1:0]                      M_AXIMM_72_RRESP,
    input  wire                            M_AXIMM_72_RLAST,
    input  wire                            M_AXIMM_72_RVALID,
    output wire                            M_AXIMM_72_RREADY,
    //AXI-MM pass-through interface 73
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_73_AWADDR,
    input wire [7:0]                      AP_AXIMM_73_AWLEN,
    input wire [2:0]                      AP_AXIMM_73_AWSIZE,
    input wire [1:0]                      AP_AXIMM_73_AWBURST,
    input wire [1:0]                      AP_AXIMM_73_AWLOCK,
    input wire [3:0]                      AP_AXIMM_73_AWCACHE,
    input wire [2:0]                      AP_AXIMM_73_AWPROT,
    input wire [3:0]                      AP_AXIMM_73_AWREGION,
    input wire [3:0]                      AP_AXIMM_73_AWQOS,
    input wire                            AP_AXIMM_73_AWVALID,
    output  wire                            AP_AXIMM_73_AWREADY,
    input wire [M_AXIMM_73_DATA_WIDTH-1:0]   AP_AXIMM_73_WDATA,
    input wire [M_AXIMM_73_DATA_WIDTH/8-1:0] AP_AXIMM_73_WSTRB,
    input wire                            AP_AXIMM_73_WLAST,
    input wire                            AP_AXIMM_73_WVALID,
    output  wire                            AP_AXIMM_73_WREADY,
    output  wire [1:0]                      AP_AXIMM_73_BRESP,
    output  wire                            AP_AXIMM_73_BVALID,
    input wire                            AP_AXIMM_73_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_73_ARADDR,
    input wire [7:0]                      AP_AXIMM_73_ARLEN,
    input wire [2:0]                      AP_AXIMM_73_ARSIZE,
    input wire [1:0]                      AP_AXIMM_73_ARBURST,
    input wire [1:0]                      AP_AXIMM_73_ARLOCK,
    input wire [3:0]                      AP_AXIMM_73_ARCACHE,
    input wire [2:0]                      AP_AXIMM_73_ARPROT,
    input wire [3:0]                      AP_AXIMM_73_ARREGION,
    input wire [3:0]                      AP_AXIMM_73_ARQOS,
    input wire                            AP_AXIMM_73_ARVALID,
    output  wire                            AP_AXIMM_73_ARREADY,
    output  wire [M_AXIMM_73_DATA_WIDTH-1:0]   AP_AXIMM_73_RDATA,
    output  wire [1:0]                      AP_AXIMM_73_RRESP,
    output  wire                            AP_AXIMM_73_RLAST,
    output  wire                            AP_AXIMM_73_RVALID,
    input  wire                            AP_AXIMM_73_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_73_AWADDR,
    output wire [7:0]                      M_AXIMM_73_AWLEN,
    output wire [2:0]                      M_AXIMM_73_AWSIZE,
    output wire [1:0]                      M_AXIMM_73_AWBURST,
    output wire [1:0]                      M_AXIMM_73_AWLOCK,
    output wire [3:0]                      M_AXIMM_73_AWCACHE,
    output wire [2:0]                      M_AXIMM_73_AWPROT,
    output wire [3:0]                      M_AXIMM_73_AWREGION,
    output wire [3:0]                      M_AXIMM_73_AWQOS,
    output wire                            M_AXIMM_73_AWVALID,
    input  wire                            M_AXIMM_73_AWREADY,
    output wire [M_AXIMM_73_DATA_WIDTH-1:0]   M_AXIMM_73_WDATA,
    output wire [M_AXIMM_73_DATA_WIDTH/8-1:0] M_AXIMM_73_WSTRB,
    output wire                            M_AXIMM_73_WLAST,
    output wire                            M_AXIMM_73_WVALID,
    input  wire                            M_AXIMM_73_WREADY,
    input  wire [1:0]                      M_AXIMM_73_BRESP,
    input  wire                            M_AXIMM_73_BVALID,
    output wire                            M_AXIMM_73_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_73_ARADDR,
    output wire [7:0]                      M_AXIMM_73_ARLEN,
    output wire [2:0]                      M_AXIMM_73_ARSIZE,
    output wire [1:0]                      M_AXIMM_73_ARBURST,
    output wire [1:0]                      M_AXIMM_73_ARLOCK,
    output wire [3:0]                      M_AXIMM_73_ARCACHE,
    output wire [2:0]                      M_AXIMM_73_ARPROT,
    output wire [3:0]                      M_AXIMM_73_ARREGION,
    output wire [3:0]                      M_AXIMM_73_ARQOS,
    output wire                            M_AXIMM_73_ARVALID,
    input  wire                            M_AXIMM_73_ARREADY,
    input  wire [M_AXIMM_73_DATA_WIDTH-1:0]   M_AXIMM_73_RDATA,
    input  wire [1:0]                      M_AXIMM_73_RRESP,
    input  wire                            M_AXIMM_73_RLAST,
    input  wire                            M_AXIMM_73_RVALID,
    output wire                            M_AXIMM_73_RREADY,
    //AXI-MM pass-through interface 74
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_74_AWADDR,
    input wire [7:0]                      AP_AXIMM_74_AWLEN,
    input wire [2:0]                      AP_AXIMM_74_AWSIZE,
    input wire [1:0]                      AP_AXIMM_74_AWBURST,
    input wire [1:0]                      AP_AXIMM_74_AWLOCK,
    input wire [3:0]                      AP_AXIMM_74_AWCACHE,
    input wire [2:0]                      AP_AXIMM_74_AWPROT,
    input wire [3:0]                      AP_AXIMM_74_AWREGION,
    input wire [3:0]                      AP_AXIMM_74_AWQOS,
    input wire                            AP_AXIMM_74_AWVALID,
    output  wire                            AP_AXIMM_74_AWREADY,
    input wire [M_AXIMM_74_DATA_WIDTH-1:0]   AP_AXIMM_74_WDATA,
    input wire [M_AXIMM_74_DATA_WIDTH/8-1:0] AP_AXIMM_74_WSTRB,
    input wire                            AP_AXIMM_74_WLAST,
    input wire                            AP_AXIMM_74_WVALID,
    output  wire                            AP_AXIMM_74_WREADY,
    output  wire [1:0]                      AP_AXIMM_74_BRESP,
    output  wire                            AP_AXIMM_74_BVALID,
    input wire                            AP_AXIMM_74_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_74_ARADDR,
    input wire [7:0]                      AP_AXIMM_74_ARLEN,
    input wire [2:0]                      AP_AXIMM_74_ARSIZE,
    input wire [1:0]                      AP_AXIMM_74_ARBURST,
    input wire [1:0]                      AP_AXIMM_74_ARLOCK,
    input wire [3:0]                      AP_AXIMM_74_ARCACHE,
    input wire [2:0]                      AP_AXIMM_74_ARPROT,
    input wire [3:0]                      AP_AXIMM_74_ARREGION,
    input wire [3:0]                      AP_AXIMM_74_ARQOS,
    input wire                            AP_AXIMM_74_ARVALID,
    output  wire                            AP_AXIMM_74_ARREADY,
    output  wire [M_AXIMM_74_DATA_WIDTH-1:0]   AP_AXIMM_74_RDATA,
    output  wire [1:0]                      AP_AXIMM_74_RRESP,
    output  wire                            AP_AXIMM_74_RLAST,
    output  wire                            AP_AXIMM_74_RVALID,
    input  wire                            AP_AXIMM_74_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_74_AWADDR,
    output wire [7:0]                      M_AXIMM_74_AWLEN,
    output wire [2:0]                      M_AXIMM_74_AWSIZE,
    output wire [1:0]                      M_AXIMM_74_AWBURST,
    output wire [1:0]                      M_AXIMM_74_AWLOCK,
    output wire [3:0]                      M_AXIMM_74_AWCACHE,
    output wire [2:0]                      M_AXIMM_74_AWPROT,
    output wire [3:0]                      M_AXIMM_74_AWREGION,
    output wire [3:0]                      M_AXIMM_74_AWQOS,
    output wire                            M_AXIMM_74_AWVALID,
    input  wire                            M_AXIMM_74_AWREADY,
    output wire [M_AXIMM_74_DATA_WIDTH-1:0]   M_AXIMM_74_WDATA,
    output wire [M_AXIMM_74_DATA_WIDTH/8-1:0] M_AXIMM_74_WSTRB,
    output wire                            M_AXIMM_74_WLAST,
    output wire                            M_AXIMM_74_WVALID,
    input  wire                            M_AXIMM_74_WREADY,
    input  wire [1:0]                      M_AXIMM_74_BRESP,
    input  wire                            M_AXIMM_74_BVALID,
    output wire                            M_AXIMM_74_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_74_ARADDR,
    output wire [7:0]                      M_AXIMM_74_ARLEN,
    output wire [2:0]                      M_AXIMM_74_ARSIZE,
    output wire [1:0]                      M_AXIMM_74_ARBURST,
    output wire [1:0]                      M_AXIMM_74_ARLOCK,
    output wire [3:0]                      M_AXIMM_74_ARCACHE,
    output wire [2:0]                      M_AXIMM_74_ARPROT,
    output wire [3:0]                      M_AXIMM_74_ARREGION,
    output wire [3:0]                      M_AXIMM_74_ARQOS,
    output wire                            M_AXIMM_74_ARVALID,
    input  wire                            M_AXIMM_74_ARREADY,
    input  wire [M_AXIMM_74_DATA_WIDTH-1:0]   M_AXIMM_74_RDATA,
    input  wire [1:0]                      M_AXIMM_74_RRESP,
    input  wire                            M_AXIMM_74_RLAST,
    input  wire                            M_AXIMM_74_RVALID,
    output wire                            M_AXIMM_74_RREADY,
    //AXI-MM pass-through interface 75
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_75_AWADDR,
    input wire [7:0]                      AP_AXIMM_75_AWLEN,
    input wire [2:0]                      AP_AXIMM_75_AWSIZE,
    input wire [1:0]                      AP_AXIMM_75_AWBURST,
    input wire [1:0]                      AP_AXIMM_75_AWLOCK,
    input wire [3:0]                      AP_AXIMM_75_AWCACHE,
    input wire [2:0]                      AP_AXIMM_75_AWPROT,
    input wire [3:0]                      AP_AXIMM_75_AWREGION,
    input wire [3:0]                      AP_AXIMM_75_AWQOS,
    input wire                            AP_AXIMM_75_AWVALID,
    output  wire                            AP_AXIMM_75_AWREADY,
    input wire [M_AXIMM_75_DATA_WIDTH-1:0]   AP_AXIMM_75_WDATA,
    input wire [M_AXIMM_75_DATA_WIDTH/8-1:0] AP_AXIMM_75_WSTRB,
    input wire                            AP_AXIMM_75_WLAST,
    input wire                            AP_AXIMM_75_WVALID,
    output  wire                            AP_AXIMM_75_WREADY,
    output  wire [1:0]                      AP_AXIMM_75_BRESP,
    output  wire                            AP_AXIMM_75_BVALID,
    input wire                            AP_AXIMM_75_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_75_ARADDR,
    input wire [7:0]                      AP_AXIMM_75_ARLEN,
    input wire [2:0]                      AP_AXIMM_75_ARSIZE,
    input wire [1:0]                      AP_AXIMM_75_ARBURST,
    input wire [1:0]                      AP_AXIMM_75_ARLOCK,
    input wire [3:0]                      AP_AXIMM_75_ARCACHE,
    input wire [2:0]                      AP_AXIMM_75_ARPROT,
    input wire [3:0]                      AP_AXIMM_75_ARREGION,
    input wire [3:0]                      AP_AXIMM_75_ARQOS,
    input wire                            AP_AXIMM_75_ARVALID,
    output  wire                            AP_AXIMM_75_ARREADY,
    output  wire [M_AXIMM_75_DATA_WIDTH-1:0]   AP_AXIMM_75_RDATA,
    output  wire [1:0]                      AP_AXIMM_75_RRESP,
    output  wire                            AP_AXIMM_75_RLAST,
    output  wire                            AP_AXIMM_75_RVALID,
    input  wire                            AP_AXIMM_75_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_75_AWADDR,
    output wire [7:0]                      M_AXIMM_75_AWLEN,
    output wire [2:0]                      M_AXIMM_75_AWSIZE,
    output wire [1:0]                      M_AXIMM_75_AWBURST,
    output wire [1:0]                      M_AXIMM_75_AWLOCK,
    output wire [3:0]                      M_AXIMM_75_AWCACHE,
    output wire [2:0]                      M_AXIMM_75_AWPROT,
    output wire [3:0]                      M_AXIMM_75_AWREGION,
    output wire [3:0]                      M_AXIMM_75_AWQOS,
    output wire                            M_AXIMM_75_AWVALID,
    input  wire                            M_AXIMM_75_AWREADY,
    output wire [M_AXIMM_75_DATA_WIDTH-1:0]   M_AXIMM_75_WDATA,
    output wire [M_AXIMM_75_DATA_WIDTH/8-1:0] M_AXIMM_75_WSTRB,
    output wire                            M_AXIMM_75_WLAST,
    output wire                            M_AXIMM_75_WVALID,
    input  wire                            M_AXIMM_75_WREADY,
    input  wire [1:0]                      M_AXIMM_75_BRESP,
    input  wire                            M_AXIMM_75_BVALID,
    output wire                            M_AXIMM_75_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_75_ARADDR,
    output wire [7:0]                      M_AXIMM_75_ARLEN,
    output wire [2:0]                      M_AXIMM_75_ARSIZE,
    output wire [1:0]                      M_AXIMM_75_ARBURST,
    output wire [1:0]                      M_AXIMM_75_ARLOCK,
    output wire [3:0]                      M_AXIMM_75_ARCACHE,
    output wire [2:0]                      M_AXIMM_75_ARPROT,
    output wire [3:0]                      M_AXIMM_75_ARREGION,
    output wire [3:0]                      M_AXIMM_75_ARQOS,
    output wire                            M_AXIMM_75_ARVALID,
    input  wire                            M_AXIMM_75_ARREADY,
    input  wire [M_AXIMM_75_DATA_WIDTH-1:0]   M_AXIMM_75_RDATA,
    input  wire [1:0]                      M_AXIMM_75_RRESP,
    input  wire                            M_AXIMM_75_RLAST,
    input  wire                            M_AXIMM_75_RVALID,
    output wire                            M_AXIMM_75_RREADY,
    //AXI-MM pass-through interface 76
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_76_AWADDR,
    input wire [7:0]                      AP_AXIMM_76_AWLEN,
    input wire [2:0]                      AP_AXIMM_76_AWSIZE,
    input wire [1:0]                      AP_AXIMM_76_AWBURST,
    input wire [1:0]                      AP_AXIMM_76_AWLOCK,
    input wire [3:0]                      AP_AXIMM_76_AWCACHE,
    input wire [2:0]                      AP_AXIMM_76_AWPROT,
    input wire [3:0]                      AP_AXIMM_76_AWREGION,
    input wire [3:0]                      AP_AXIMM_76_AWQOS,
    input wire                            AP_AXIMM_76_AWVALID,
    output  wire                            AP_AXIMM_76_AWREADY,
    input wire [M_AXIMM_76_DATA_WIDTH-1:0]   AP_AXIMM_76_WDATA,
    input wire [M_AXIMM_76_DATA_WIDTH/8-1:0] AP_AXIMM_76_WSTRB,
    input wire                            AP_AXIMM_76_WLAST,
    input wire                            AP_AXIMM_76_WVALID,
    output  wire                            AP_AXIMM_76_WREADY,
    output  wire [1:0]                      AP_AXIMM_76_BRESP,
    output  wire                            AP_AXIMM_76_BVALID,
    input wire                            AP_AXIMM_76_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_76_ARADDR,
    input wire [7:0]                      AP_AXIMM_76_ARLEN,
    input wire [2:0]                      AP_AXIMM_76_ARSIZE,
    input wire [1:0]                      AP_AXIMM_76_ARBURST,
    input wire [1:0]                      AP_AXIMM_76_ARLOCK,
    input wire [3:0]                      AP_AXIMM_76_ARCACHE,
    input wire [2:0]                      AP_AXIMM_76_ARPROT,
    input wire [3:0]                      AP_AXIMM_76_ARREGION,
    input wire [3:0]                      AP_AXIMM_76_ARQOS,
    input wire                            AP_AXIMM_76_ARVALID,
    output  wire                            AP_AXIMM_76_ARREADY,
    output  wire [M_AXIMM_76_DATA_WIDTH-1:0]   AP_AXIMM_76_RDATA,
    output  wire [1:0]                      AP_AXIMM_76_RRESP,
    output  wire                            AP_AXIMM_76_RLAST,
    output  wire                            AP_AXIMM_76_RVALID,
    input  wire                            AP_AXIMM_76_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_76_AWADDR,
    output wire [7:0]                      M_AXIMM_76_AWLEN,
    output wire [2:0]                      M_AXIMM_76_AWSIZE,
    output wire [1:0]                      M_AXIMM_76_AWBURST,
    output wire [1:0]                      M_AXIMM_76_AWLOCK,
    output wire [3:0]                      M_AXIMM_76_AWCACHE,
    output wire [2:0]                      M_AXIMM_76_AWPROT,
    output wire [3:0]                      M_AXIMM_76_AWREGION,
    output wire [3:0]                      M_AXIMM_76_AWQOS,
    output wire                            M_AXIMM_76_AWVALID,
    input  wire                            M_AXIMM_76_AWREADY,
    output wire [M_AXIMM_76_DATA_WIDTH-1:0]   M_AXIMM_76_WDATA,
    output wire [M_AXIMM_76_DATA_WIDTH/8-1:0] M_AXIMM_76_WSTRB,
    output wire                            M_AXIMM_76_WLAST,
    output wire                            M_AXIMM_76_WVALID,
    input  wire                            M_AXIMM_76_WREADY,
    input  wire [1:0]                      M_AXIMM_76_BRESP,
    input  wire                            M_AXIMM_76_BVALID,
    output wire                            M_AXIMM_76_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_76_ARADDR,
    output wire [7:0]                      M_AXIMM_76_ARLEN,
    output wire [2:0]                      M_AXIMM_76_ARSIZE,
    output wire [1:0]                      M_AXIMM_76_ARBURST,
    output wire [1:0]                      M_AXIMM_76_ARLOCK,
    output wire [3:0]                      M_AXIMM_76_ARCACHE,
    output wire [2:0]                      M_AXIMM_76_ARPROT,
    output wire [3:0]                      M_AXIMM_76_ARREGION,
    output wire [3:0]                      M_AXIMM_76_ARQOS,
    output wire                            M_AXIMM_76_ARVALID,
    input  wire                            M_AXIMM_76_ARREADY,
    input  wire [M_AXIMM_76_DATA_WIDTH-1:0]   M_AXIMM_76_RDATA,
    input  wire [1:0]                      M_AXIMM_76_RRESP,
    input  wire                            M_AXIMM_76_RLAST,
    input  wire                            M_AXIMM_76_RVALID,
    output wire                            M_AXIMM_76_RREADY,
    //AXI-MM pass-through interface 77
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_77_AWADDR,
    input wire [7:0]                      AP_AXIMM_77_AWLEN,
    input wire [2:0]                      AP_AXIMM_77_AWSIZE,
    input wire [1:0]                      AP_AXIMM_77_AWBURST,
    input wire [1:0]                      AP_AXIMM_77_AWLOCK,
    input wire [3:0]                      AP_AXIMM_77_AWCACHE,
    input wire [2:0]                      AP_AXIMM_77_AWPROT,
    input wire [3:0]                      AP_AXIMM_77_AWREGION,
    input wire [3:0]                      AP_AXIMM_77_AWQOS,
    input wire                            AP_AXIMM_77_AWVALID,
    output  wire                            AP_AXIMM_77_AWREADY,
    input wire [M_AXIMM_77_DATA_WIDTH-1:0]   AP_AXIMM_77_WDATA,
    input wire [M_AXIMM_77_DATA_WIDTH/8-1:0] AP_AXIMM_77_WSTRB,
    input wire                            AP_AXIMM_77_WLAST,
    input wire                            AP_AXIMM_77_WVALID,
    output  wire                            AP_AXIMM_77_WREADY,
    output  wire [1:0]                      AP_AXIMM_77_BRESP,
    output  wire                            AP_AXIMM_77_BVALID,
    input wire                            AP_AXIMM_77_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_77_ARADDR,
    input wire [7:0]                      AP_AXIMM_77_ARLEN,
    input wire [2:0]                      AP_AXIMM_77_ARSIZE,
    input wire [1:0]                      AP_AXIMM_77_ARBURST,
    input wire [1:0]                      AP_AXIMM_77_ARLOCK,
    input wire [3:0]                      AP_AXIMM_77_ARCACHE,
    input wire [2:0]                      AP_AXIMM_77_ARPROT,
    input wire [3:0]                      AP_AXIMM_77_ARREGION,
    input wire [3:0]                      AP_AXIMM_77_ARQOS,
    input wire                            AP_AXIMM_77_ARVALID,
    output  wire                            AP_AXIMM_77_ARREADY,
    output  wire [M_AXIMM_77_DATA_WIDTH-1:0]   AP_AXIMM_77_RDATA,
    output  wire [1:0]                      AP_AXIMM_77_RRESP,
    output  wire                            AP_AXIMM_77_RLAST,
    output  wire                            AP_AXIMM_77_RVALID,
    input  wire                            AP_AXIMM_77_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_77_AWADDR,
    output wire [7:0]                      M_AXIMM_77_AWLEN,
    output wire [2:0]                      M_AXIMM_77_AWSIZE,
    output wire [1:0]                      M_AXIMM_77_AWBURST,
    output wire [1:0]                      M_AXIMM_77_AWLOCK,
    output wire [3:0]                      M_AXIMM_77_AWCACHE,
    output wire [2:0]                      M_AXIMM_77_AWPROT,
    output wire [3:0]                      M_AXIMM_77_AWREGION,
    output wire [3:0]                      M_AXIMM_77_AWQOS,
    output wire                            M_AXIMM_77_AWVALID,
    input  wire                            M_AXIMM_77_AWREADY,
    output wire [M_AXIMM_77_DATA_WIDTH-1:0]   M_AXIMM_77_WDATA,
    output wire [M_AXIMM_77_DATA_WIDTH/8-1:0] M_AXIMM_77_WSTRB,
    output wire                            M_AXIMM_77_WLAST,
    output wire                            M_AXIMM_77_WVALID,
    input  wire                            M_AXIMM_77_WREADY,
    input  wire [1:0]                      M_AXIMM_77_BRESP,
    input  wire                            M_AXIMM_77_BVALID,
    output wire                            M_AXIMM_77_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_77_ARADDR,
    output wire [7:0]                      M_AXIMM_77_ARLEN,
    output wire [2:0]                      M_AXIMM_77_ARSIZE,
    output wire [1:0]                      M_AXIMM_77_ARBURST,
    output wire [1:0]                      M_AXIMM_77_ARLOCK,
    output wire [3:0]                      M_AXIMM_77_ARCACHE,
    output wire [2:0]                      M_AXIMM_77_ARPROT,
    output wire [3:0]                      M_AXIMM_77_ARREGION,
    output wire [3:0]                      M_AXIMM_77_ARQOS,
    output wire                            M_AXIMM_77_ARVALID,
    input  wire                            M_AXIMM_77_ARREADY,
    input  wire [M_AXIMM_77_DATA_WIDTH-1:0]   M_AXIMM_77_RDATA,
    input  wire [1:0]                      M_AXIMM_77_RRESP,
    input  wire                            M_AXIMM_77_RLAST,
    input  wire                            M_AXIMM_77_RVALID,
    output wire                            M_AXIMM_77_RREADY,
    //AXI-MM pass-through interface 78
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_78_AWADDR,
    input wire [7:0]                      AP_AXIMM_78_AWLEN,
    input wire [2:0]                      AP_AXIMM_78_AWSIZE,
    input wire [1:0]                      AP_AXIMM_78_AWBURST,
    input wire [1:0]                      AP_AXIMM_78_AWLOCK,
    input wire [3:0]                      AP_AXIMM_78_AWCACHE,
    input wire [2:0]                      AP_AXIMM_78_AWPROT,
    input wire [3:0]                      AP_AXIMM_78_AWREGION,
    input wire [3:0]                      AP_AXIMM_78_AWQOS,
    input wire                            AP_AXIMM_78_AWVALID,
    output  wire                            AP_AXIMM_78_AWREADY,
    input wire [M_AXIMM_78_DATA_WIDTH-1:0]   AP_AXIMM_78_WDATA,
    input wire [M_AXIMM_78_DATA_WIDTH/8-1:0] AP_AXIMM_78_WSTRB,
    input wire                            AP_AXIMM_78_WLAST,
    input wire                            AP_AXIMM_78_WVALID,
    output  wire                            AP_AXIMM_78_WREADY,
    output  wire [1:0]                      AP_AXIMM_78_BRESP,
    output  wire                            AP_AXIMM_78_BVALID,
    input wire                            AP_AXIMM_78_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_78_ARADDR,
    input wire [7:0]                      AP_AXIMM_78_ARLEN,
    input wire [2:0]                      AP_AXIMM_78_ARSIZE,
    input wire [1:0]                      AP_AXIMM_78_ARBURST,
    input wire [1:0]                      AP_AXIMM_78_ARLOCK,
    input wire [3:0]                      AP_AXIMM_78_ARCACHE,
    input wire [2:0]                      AP_AXIMM_78_ARPROT,
    input wire [3:0]                      AP_AXIMM_78_ARREGION,
    input wire [3:0]                      AP_AXIMM_78_ARQOS,
    input wire                            AP_AXIMM_78_ARVALID,
    output  wire                            AP_AXIMM_78_ARREADY,
    output  wire [M_AXIMM_78_DATA_WIDTH-1:0]   AP_AXIMM_78_RDATA,
    output  wire [1:0]                      AP_AXIMM_78_RRESP,
    output  wire                            AP_AXIMM_78_RLAST,
    output  wire                            AP_AXIMM_78_RVALID,
    input  wire                            AP_AXIMM_78_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_78_AWADDR,
    output wire [7:0]                      M_AXIMM_78_AWLEN,
    output wire [2:0]                      M_AXIMM_78_AWSIZE,
    output wire [1:0]                      M_AXIMM_78_AWBURST,
    output wire [1:0]                      M_AXIMM_78_AWLOCK,
    output wire [3:0]                      M_AXIMM_78_AWCACHE,
    output wire [2:0]                      M_AXIMM_78_AWPROT,
    output wire [3:0]                      M_AXIMM_78_AWREGION,
    output wire [3:0]                      M_AXIMM_78_AWQOS,
    output wire                            M_AXIMM_78_AWVALID,
    input  wire                            M_AXIMM_78_AWREADY,
    output wire [M_AXIMM_78_DATA_WIDTH-1:0]   M_AXIMM_78_WDATA,
    output wire [M_AXIMM_78_DATA_WIDTH/8-1:0] M_AXIMM_78_WSTRB,
    output wire                            M_AXIMM_78_WLAST,
    output wire                            M_AXIMM_78_WVALID,
    input  wire                            M_AXIMM_78_WREADY,
    input  wire [1:0]                      M_AXIMM_78_BRESP,
    input  wire                            M_AXIMM_78_BVALID,
    output wire                            M_AXIMM_78_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_78_ARADDR,
    output wire [7:0]                      M_AXIMM_78_ARLEN,
    output wire [2:0]                      M_AXIMM_78_ARSIZE,
    output wire [1:0]                      M_AXIMM_78_ARBURST,
    output wire [1:0]                      M_AXIMM_78_ARLOCK,
    output wire [3:0]                      M_AXIMM_78_ARCACHE,
    output wire [2:0]                      M_AXIMM_78_ARPROT,
    output wire [3:0]                      M_AXIMM_78_ARREGION,
    output wire [3:0]                      M_AXIMM_78_ARQOS,
    output wire                            M_AXIMM_78_ARVALID,
    input  wire                            M_AXIMM_78_ARREADY,
    input  wire [M_AXIMM_78_DATA_WIDTH-1:0]   M_AXIMM_78_RDATA,
    input  wire [1:0]                      M_AXIMM_78_RRESP,
    input  wire                            M_AXIMM_78_RLAST,
    input  wire                            M_AXIMM_78_RVALID,
    output wire                            M_AXIMM_78_RREADY,
    //AXI-MM pass-through interface 79
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_79_AWADDR,
    input wire [7:0]                      AP_AXIMM_79_AWLEN,
    input wire [2:0]                      AP_AXIMM_79_AWSIZE,
    input wire [1:0]                      AP_AXIMM_79_AWBURST,
    input wire [1:0]                      AP_AXIMM_79_AWLOCK,
    input wire [3:0]                      AP_AXIMM_79_AWCACHE,
    input wire [2:0]                      AP_AXIMM_79_AWPROT,
    input wire [3:0]                      AP_AXIMM_79_AWREGION,
    input wire [3:0]                      AP_AXIMM_79_AWQOS,
    input wire                            AP_AXIMM_79_AWVALID,
    output  wire                            AP_AXIMM_79_AWREADY,
    input wire [M_AXIMM_79_DATA_WIDTH-1:0]   AP_AXIMM_79_WDATA,
    input wire [M_AXIMM_79_DATA_WIDTH/8-1:0] AP_AXIMM_79_WSTRB,
    input wire                            AP_AXIMM_79_WLAST,
    input wire                            AP_AXIMM_79_WVALID,
    output  wire                            AP_AXIMM_79_WREADY,
    output  wire [1:0]                      AP_AXIMM_79_BRESP,
    output  wire                            AP_AXIMM_79_BVALID,
    input wire                            AP_AXIMM_79_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_79_ARADDR,
    input wire [7:0]                      AP_AXIMM_79_ARLEN,
    input wire [2:0]                      AP_AXIMM_79_ARSIZE,
    input wire [1:0]                      AP_AXIMM_79_ARBURST,
    input wire [1:0]                      AP_AXIMM_79_ARLOCK,
    input wire [3:0]                      AP_AXIMM_79_ARCACHE,
    input wire [2:0]                      AP_AXIMM_79_ARPROT,
    input wire [3:0]                      AP_AXIMM_79_ARREGION,
    input wire [3:0]                      AP_AXIMM_79_ARQOS,
    input wire                            AP_AXIMM_79_ARVALID,
    output  wire                            AP_AXIMM_79_ARREADY,
    output  wire [M_AXIMM_79_DATA_WIDTH-1:0]   AP_AXIMM_79_RDATA,
    output  wire [1:0]                      AP_AXIMM_79_RRESP,
    output  wire                            AP_AXIMM_79_RLAST,
    output  wire                            AP_AXIMM_79_RVALID,
    input  wire                            AP_AXIMM_79_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_79_AWADDR,
    output wire [7:0]                      M_AXIMM_79_AWLEN,
    output wire [2:0]                      M_AXIMM_79_AWSIZE,
    output wire [1:0]                      M_AXIMM_79_AWBURST,
    output wire [1:0]                      M_AXIMM_79_AWLOCK,
    output wire [3:0]                      M_AXIMM_79_AWCACHE,
    output wire [2:0]                      M_AXIMM_79_AWPROT,
    output wire [3:0]                      M_AXIMM_79_AWREGION,
    output wire [3:0]                      M_AXIMM_79_AWQOS,
    output wire                            M_AXIMM_79_AWVALID,
    input  wire                            M_AXIMM_79_AWREADY,
    output wire [M_AXIMM_79_DATA_WIDTH-1:0]   M_AXIMM_79_WDATA,
    output wire [M_AXIMM_79_DATA_WIDTH/8-1:0] M_AXIMM_79_WSTRB,
    output wire                            M_AXIMM_79_WLAST,
    output wire                            M_AXIMM_79_WVALID,
    input  wire                            M_AXIMM_79_WREADY,
    input  wire [1:0]                      M_AXIMM_79_BRESP,
    input  wire                            M_AXIMM_79_BVALID,
    output wire                            M_AXIMM_79_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_79_ARADDR,
    output wire [7:0]                      M_AXIMM_79_ARLEN,
    output wire [2:0]                      M_AXIMM_79_ARSIZE,
    output wire [1:0]                      M_AXIMM_79_ARBURST,
    output wire [1:0]                      M_AXIMM_79_ARLOCK,
    output wire [3:0]                      M_AXIMM_79_ARCACHE,
    output wire [2:0]                      M_AXIMM_79_ARPROT,
    output wire [3:0]                      M_AXIMM_79_ARREGION,
    output wire [3:0]                      M_AXIMM_79_ARQOS,
    output wire                            M_AXIMM_79_ARVALID,
    input  wire                            M_AXIMM_79_ARREADY,
    input  wire [M_AXIMM_79_DATA_WIDTH-1:0]   M_AXIMM_79_RDATA,
    input  wire [1:0]                      M_AXIMM_79_RRESP,
    input  wire                            M_AXIMM_79_RLAST,
    input  wire                            M_AXIMM_79_RVALID,
    output wire                            M_AXIMM_79_RREADY,
    //AXI-MM pass-through interface 80
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_80_AWADDR,
    input wire [7:0]                      AP_AXIMM_80_AWLEN,
    input wire [2:0]                      AP_AXIMM_80_AWSIZE,
    input wire [1:0]                      AP_AXIMM_80_AWBURST,
    input wire [1:0]                      AP_AXIMM_80_AWLOCK,
    input wire [3:0]                      AP_AXIMM_80_AWCACHE,
    input wire [2:0]                      AP_AXIMM_80_AWPROT,
    input wire [3:0]                      AP_AXIMM_80_AWREGION,
    input wire [3:0]                      AP_AXIMM_80_AWQOS,
    input wire                            AP_AXIMM_80_AWVALID,
    output  wire                            AP_AXIMM_80_AWREADY,
    input wire [M_AXIMM_80_DATA_WIDTH-1:0]   AP_AXIMM_80_WDATA,
    input wire [M_AXIMM_80_DATA_WIDTH/8-1:0] AP_AXIMM_80_WSTRB,
    input wire                            AP_AXIMM_80_WLAST,
    input wire                            AP_AXIMM_80_WVALID,
    output  wire                            AP_AXIMM_80_WREADY,
    output  wire [1:0]                      AP_AXIMM_80_BRESP,
    output  wire                            AP_AXIMM_80_BVALID,
    input wire                            AP_AXIMM_80_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_80_ARADDR,
    input wire [7:0]                      AP_AXIMM_80_ARLEN,
    input wire [2:0]                      AP_AXIMM_80_ARSIZE,
    input wire [1:0]                      AP_AXIMM_80_ARBURST,
    input wire [1:0]                      AP_AXIMM_80_ARLOCK,
    input wire [3:0]                      AP_AXIMM_80_ARCACHE,
    input wire [2:0]                      AP_AXIMM_80_ARPROT,
    input wire [3:0]                      AP_AXIMM_80_ARREGION,
    input wire [3:0]                      AP_AXIMM_80_ARQOS,
    input wire                            AP_AXIMM_80_ARVALID,
    output  wire                            AP_AXIMM_80_ARREADY,
    output  wire [M_AXIMM_80_DATA_WIDTH-1:0]   AP_AXIMM_80_RDATA,
    output  wire [1:0]                      AP_AXIMM_80_RRESP,
    output  wire                            AP_AXIMM_80_RLAST,
    output  wire                            AP_AXIMM_80_RVALID,
    input  wire                            AP_AXIMM_80_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_80_AWADDR,
    output wire [7:0]                      M_AXIMM_80_AWLEN,
    output wire [2:0]                      M_AXIMM_80_AWSIZE,
    output wire [1:0]                      M_AXIMM_80_AWBURST,
    output wire [1:0]                      M_AXIMM_80_AWLOCK,
    output wire [3:0]                      M_AXIMM_80_AWCACHE,
    output wire [2:0]                      M_AXIMM_80_AWPROT,
    output wire [3:0]                      M_AXIMM_80_AWREGION,
    output wire [3:0]                      M_AXIMM_80_AWQOS,
    output wire                            M_AXIMM_80_AWVALID,
    input  wire                            M_AXIMM_80_AWREADY,
    output wire [M_AXIMM_80_DATA_WIDTH-1:0]   M_AXIMM_80_WDATA,
    output wire [M_AXIMM_80_DATA_WIDTH/8-1:0] M_AXIMM_80_WSTRB,
    output wire                            M_AXIMM_80_WLAST,
    output wire                            M_AXIMM_80_WVALID,
    input  wire                            M_AXIMM_80_WREADY,
    input  wire [1:0]                      M_AXIMM_80_BRESP,
    input  wire                            M_AXIMM_80_BVALID,
    output wire                            M_AXIMM_80_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_80_ARADDR,
    output wire [7:0]                      M_AXIMM_80_ARLEN,
    output wire [2:0]                      M_AXIMM_80_ARSIZE,
    output wire [1:0]                      M_AXIMM_80_ARBURST,
    output wire [1:0]                      M_AXIMM_80_ARLOCK,
    output wire [3:0]                      M_AXIMM_80_ARCACHE,
    output wire [2:0]                      M_AXIMM_80_ARPROT,
    output wire [3:0]                      M_AXIMM_80_ARREGION,
    output wire [3:0]                      M_AXIMM_80_ARQOS,
    output wire                            M_AXIMM_80_ARVALID,
    input  wire                            M_AXIMM_80_ARREADY,
    input  wire [M_AXIMM_80_DATA_WIDTH-1:0]   M_AXIMM_80_RDATA,
    input  wire [1:0]                      M_AXIMM_80_RRESP,
    input  wire                            M_AXIMM_80_RLAST,
    input  wire                            M_AXIMM_80_RVALID,
    output wire                            M_AXIMM_80_RREADY,
    //AXI-MM pass-through interface 81
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_81_AWADDR,
    input wire [7:0]                      AP_AXIMM_81_AWLEN,
    input wire [2:0]                      AP_AXIMM_81_AWSIZE,
    input wire [1:0]                      AP_AXIMM_81_AWBURST,
    input wire [1:0]                      AP_AXIMM_81_AWLOCK,
    input wire [3:0]                      AP_AXIMM_81_AWCACHE,
    input wire [2:0]                      AP_AXIMM_81_AWPROT,
    input wire [3:0]                      AP_AXIMM_81_AWREGION,
    input wire [3:0]                      AP_AXIMM_81_AWQOS,
    input wire                            AP_AXIMM_81_AWVALID,
    output  wire                            AP_AXIMM_81_AWREADY,
    input wire [M_AXIMM_81_DATA_WIDTH-1:0]   AP_AXIMM_81_WDATA,
    input wire [M_AXIMM_81_DATA_WIDTH/8-1:0] AP_AXIMM_81_WSTRB,
    input wire                            AP_AXIMM_81_WLAST,
    input wire                            AP_AXIMM_81_WVALID,
    output  wire                            AP_AXIMM_81_WREADY,
    output  wire [1:0]                      AP_AXIMM_81_BRESP,
    output  wire                            AP_AXIMM_81_BVALID,
    input wire                            AP_AXIMM_81_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_81_ARADDR,
    input wire [7:0]                      AP_AXIMM_81_ARLEN,
    input wire [2:0]                      AP_AXIMM_81_ARSIZE,
    input wire [1:0]                      AP_AXIMM_81_ARBURST,
    input wire [1:0]                      AP_AXIMM_81_ARLOCK,
    input wire [3:0]                      AP_AXIMM_81_ARCACHE,
    input wire [2:0]                      AP_AXIMM_81_ARPROT,
    input wire [3:0]                      AP_AXIMM_81_ARREGION,
    input wire [3:0]                      AP_AXIMM_81_ARQOS,
    input wire                            AP_AXIMM_81_ARVALID,
    output  wire                            AP_AXIMM_81_ARREADY,
    output  wire [M_AXIMM_81_DATA_WIDTH-1:0]   AP_AXIMM_81_RDATA,
    output  wire [1:0]                      AP_AXIMM_81_RRESP,
    output  wire                            AP_AXIMM_81_RLAST,
    output  wire                            AP_AXIMM_81_RVALID,
    input  wire                            AP_AXIMM_81_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_81_AWADDR,
    output wire [7:0]                      M_AXIMM_81_AWLEN,
    output wire [2:0]                      M_AXIMM_81_AWSIZE,
    output wire [1:0]                      M_AXIMM_81_AWBURST,
    output wire [1:0]                      M_AXIMM_81_AWLOCK,
    output wire [3:0]                      M_AXIMM_81_AWCACHE,
    output wire [2:0]                      M_AXIMM_81_AWPROT,
    output wire [3:0]                      M_AXIMM_81_AWREGION,
    output wire [3:0]                      M_AXIMM_81_AWQOS,
    output wire                            M_AXIMM_81_AWVALID,
    input  wire                            M_AXIMM_81_AWREADY,
    output wire [M_AXIMM_81_DATA_WIDTH-1:0]   M_AXIMM_81_WDATA,
    output wire [M_AXIMM_81_DATA_WIDTH/8-1:0] M_AXIMM_81_WSTRB,
    output wire                            M_AXIMM_81_WLAST,
    output wire                            M_AXIMM_81_WVALID,
    input  wire                            M_AXIMM_81_WREADY,
    input  wire [1:0]                      M_AXIMM_81_BRESP,
    input  wire                            M_AXIMM_81_BVALID,
    output wire                            M_AXIMM_81_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_81_ARADDR,
    output wire [7:0]                      M_AXIMM_81_ARLEN,
    output wire [2:0]                      M_AXIMM_81_ARSIZE,
    output wire [1:0]                      M_AXIMM_81_ARBURST,
    output wire [1:0]                      M_AXIMM_81_ARLOCK,
    output wire [3:0]                      M_AXIMM_81_ARCACHE,
    output wire [2:0]                      M_AXIMM_81_ARPROT,
    output wire [3:0]                      M_AXIMM_81_ARREGION,
    output wire [3:0]                      M_AXIMM_81_ARQOS,
    output wire                            M_AXIMM_81_ARVALID,
    input  wire                            M_AXIMM_81_ARREADY,
    input  wire [M_AXIMM_81_DATA_WIDTH-1:0]   M_AXIMM_81_RDATA,
    input  wire [1:0]                      M_AXIMM_81_RRESP,
    input  wire                            M_AXIMM_81_RLAST,
    input  wire                            M_AXIMM_81_RVALID,
    output wire                            M_AXIMM_81_RREADY,
    //AXI-MM pass-through interface 82
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_82_AWADDR,
    input wire [7:0]                      AP_AXIMM_82_AWLEN,
    input wire [2:0]                      AP_AXIMM_82_AWSIZE,
    input wire [1:0]                      AP_AXIMM_82_AWBURST,
    input wire [1:0]                      AP_AXIMM_82_AWLOCK,
    input wire [3:0]                      AP_AXIMM_82_AWCACHE,
    input wire [2:0]                      AP_AXIMM_82_AWPROT,
    input wire [3:0]                      AP_AXIMM_82_AWREGION,
    input wire [3:0]                      AP_AXIMM_82_AWQOS,
    input wire                            AP_AXIMM_82_AWVALID,
    output  wire                            AP_AXIMM_82_AWREADY,
    input wire [M_AXIMM_82_DATA_WIDTH-1:0]   AP_AXIMM_82_WDATA,
    input wire [M_AXIMM_82_DATA_WIDTH/8-1:0] AP_AXIMM_82_WSTRB,
    input wire                            AP_AXIMM_82_WLAST,
    input wire                            AP_AXIMM_82_WVALID,
    output  wire                            AP_AXIMM_82_WREADY,
    output  wire [1:0]                      AP_AXIMM_82_BRESP,
    output  wire                            AP_AXIMM_82_BVALID,
    input wire                            AP_AXIMM_82_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_82_ARADDR,
    input wire [7:0]                      AP_AXIMM_82_ARLEN,
    input wire [2:0]                      AP_AXIMM_82_ARSIZE,
    input wire [1:0]                      AP_AXIMM_82_ARBURST,
    input wire [1:0]                      AP_AXIMM_82_ARLOCK,
    input wire [3:0]                      AP_AXIMM_82_ARCACHE,
    input wire [2:0]                      AP_AXIMM_82_ARPROT,
    input wire [3:0]                      AP_AXIMM_82_ARREGION,
    input wire [3:0]                      AP_AXIMM_82_ARQOS,
    input wire                            AP_AXIMM_82_ARVALID,
    output  wire                            AP_AXIMM_82_ARREADY,
    output  wire [M_AXIMM_82_DATA_WIDTH-1:0]   AP_AXIMM_82_RDATA,
    output  wire [1:0]                      AP_AXIMM_82_RRESP,
    output  wire                            AP_AXIMM_82_RLAST,
    output  wire                            AP_AXIMM_82_RVALID,
    input  wire                            AP_AXIMM_82_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_82_AWADDR,
    output wire [7:0]                      M_AXIMM_82_AWLEN,
    output wire [2:0]                      M_AXIMM_82_AWSIZE,
    output wire [1:0]                      M_AXIMM_82_AWBURST,
    output wire [1:0]                      M_AXIMM_82_AWLOCK,
    output wire [3:0]                      M_AXIMM_82_AWCACHE,
    output wire [2:0]                      M_AXIMM_82_AWPROT,
    output wire [3:0]                      M_AXIMM_82_AWREGION,
    output wire [3:0]                      M_AXIMM_82_AWQOS,
    output wire                            M_AXIMM_82_AWVALID,
    input  wire                            M_AXIMM_82_AWREADY,
    output wire [M_AXIMM_82_DATA_WIDTH-1:0]   M_AXIMM_82_WDATA,
    output wire [M_AXIMM_82_DATA_WIDTH/8-1:0] M_AXIMM_82_WSTRB,
    output wire                            M_AXIMM_82_WLAST,
    output wire                            M_AXIMM_82_WVALID,
    input  wire                            M_AXIMM_82_WREADY,
    input  wire [1:0]                      M_AXIMM_82_BRESP,
    input  wire                            M_AXIMM_82_BVALID,
    output wire                            M_AXIMM_82_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_82_ARADDR,
    output wire [7:0]                      M_AXIMM_82_ARLEN,
    output wire [2:0]                      M_AXIMM_82_ARSIZE,
    output wire [1:0]                      M_AXIMM_82_ARBURST,
    output wire [1:0]                      M_AXIMM_82_ARLOCK,
    output wire [3:0]                      M_AXIMM_82_ARCACHE,
    output wire [2:0]                      M_AXIMM_82_ARPROT,
    output wire [3:0]                      M_AXIMM_82_ARREGION,
    output wire [3:0]                      M_AXIMM_82_ARQOS,
    output wire                            M_AXIMM_82_ARVALID,
    input  wire                            M_AXIMM_82_ARREADY,
    input  wire [M_AXIMM_82_DATA_WIDTH-1:0]   M_AXIMM_82_RDATA,
    input  wire [1:0]                      M_AXIMM_82_RRESP,
    input  wire                            M_AXIMM_82_RLAST,
    input  wire                            M_AXIMM_82_RVALID,
    output wire                            M_AXIMM_82_RREADY,
    //AXI-MM pass-through interface 83
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_83_AWADDR,
    input wire [7:0]                      AP_AXIMM_83_AWLEN,
    input wire [2:0]                      AP_AXIMM_83_AWSIZE,
    input wire [1:0]                      AP_AXIMM_83_AWBURST,
    input wire [1:0]                      AP_AXIMM_83_AWLOCK,
    input wire [3:0]                      AP_AXIMM_83_AWCACHE,
    input wire [2:0]                      AP_AXIMM_83_AWPROT,
    input wire [3:0]                      AP_AXIMM_83_AWREGION,
    input wire [3:0]                      AP_AXIMM_83_AWQOS,
    input wire                            AP_AXIMM_83_AWVALID,
    output  wire                            AP_AXIMM_83_AWREADY,
    input wire [M_AXIMM_83_DATA_WIDTH-1:0]   AP_AXIMM_83_WDATA,
    input wire [M_AXIMM_83_DATA_WIDTH/8-1:0] AP_AXIMM_83_WSTRB,
    input wire                            AP_AXIMM_83_WLAST,
    input wire                            AP_AXIMM_83_WVALID,
    output  wire                            AP_AXIMM_83_WREADY,
    output  wire [1:0]                      AP_AXIMM_83_BRESP,
    output  wire                            AP_AXIMM_83_BVALID,
    input wire                            AP_AXIMM_83_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_83_ARADDR,
    input wire [7:0]                      AP_AXIMM_83_ARLEN,
    input wire [2:0]                      AP_AXIMM_83_ARSIZE,
    input wire [1:0]                      AP_AXIMM_83_ARBURST,
    input wire [1:0]                      AP_AXIMM_83_ARLOCK,
    input wire [3:0]                      AP_AXIMM_83_ARCACHE,
    input wire [2:0]                      AP_AXIMM_83_ARPROT,
    input wire [3:0]                      AP_AXIMM_83_ARREGION,
    input wire [3:0]                      AP_AXIMM_83_ARQOS,
    input wire                            AP_AXIMM_83_ARVALID,
    output  wire                            AP_AXIMM_83_ARREADY,
    output  wire [M_AXIMM_83_DATA_WIDTH-1:0]   AP_AXIMM_83_RDATA,
    output  wire [1:0]                      AP_AXIMM_83_RRESP,
    output  wire                            AP_AXIMM_83_RLAST,
    output  wire                            AP_AXIMM_83_RVALID,
    input  wire                            AP_AXIMM_83_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_83_AWADDR,
    output wire [7:0]                      M_AXIMM_83_AWLEN,
    output wire [2:0]                      M_AXIMM_83_AWSIZE,
    output wire [1:0]                      M_AXIMM_83_AWBURST,
    output wire [1:0]                      M_AXIMM_83_AWLOCK,
    output wire [3:0]                      M_AXIMM_83_AWCACHE,
    output wire [2:0]                      M_AXIMM_83_AWPROT,
    output wire [3:0]                      M_AXIMM_83_AWREGION,
    output wire [3:0]                      M_AXIMM_83_AWQOS,
    output wire                            M_AXIMM_83_AWVALID,
    input  wire                            M_AXIMM_83_AWREADY,
    output wire [M_AXIMM_83_DATA_WIDTH-1:0]   M_AXIMM_83_WDATA,
    output wire [M_AXIMM_83_DATA_WIDTH/8-1:0] M_AXIMM_83_WSTRB,
    output wire                            M_AXIMM_83_WLAST,
    output wire                            M_AXIMM_83_WVALID,
    input  wire                            M_AXIMM_83_WREADY,
    input  wire [1:0]                      M_AXIMM_83_BRESP,
    input  wire                            M_AXIMM_83_BVALID,
    output wire                            M_AXIMM_83_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_83_ARADDR,
    output wire [7:0]                      M_AXIMM_83_ARLEN,
    output wire [2:0]                      M_AXIMM_83_ARSIZE,
    output wire [1:0]                      M_AXIMM_83_ARBURST,
    output wire [1:0]                      M_AXIMM_83_ARLOCK,
    output wire [3:0]                      M_AXIMM_83_ARCACHE,
    output wire [2:0]                      M_AXIMM_83_ARPROT,
    output wire [3:0]                      M_AXIMM_83_ARREGION,
    output wire [3:0]                      M_AXIMM_83_ARQOS,
    output wire                            M_AXIMM_83_ARVALID,
    input  wire                            M_AXIMM_83_ARREADY,
    input  wire [M_AXIMM_83_DATA_WIDTH-1:0]   M_AXIMM_83_RDATA,
    input  wire [1:0]                      M_AXIMM_83_RRESP,
    input  wire                            M_AXIMM_83_RLAST,
    input  wire                            M_AXIMM_83_RVALID,
    output wire                            M_AXIMM_83_RREADY,
    //AXI-MM pass-through interface 84
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_84_AWADDR,
    input wire [7:0]                      AP_AXIMM_84_AWLEN,
    input wire [2:0]                      AP_AXIMM_84_AWSIZE,
    input wire [1:0]                      AP_AXIMM_84_AWBURST,
    input wire [1:0]                      AP_AXIMM_84_AWLOCK,
    input wire [3:0]                      AP_AXIMM_84_AWCACHE,
    input wire [2:0]                      AP_AXIMM_84_AWPROT,
    input wire [3:0]                      AP_AXIMM_84_AWREGION,
    input wire [3:0]                      AP_AXIMM_84_AWQOS,
    input wire                            AP_AXIMM_84_AWVALID,
    output  wire                            AP_AXIMM_84_AWREADY,
    input wire [M_AXIMM_84_DATA_WIDTH-1:0]   AP_AXIMM_84_WDATA,
    input wire [M_AXIMM_84_DATA_WIDTH/8-1:0] AP_AXIMM_84_WSTRB,
    input wire                            AP_AXIMM_84_WLAST,
    input wire                            AP_AXIMM_84_WVALID,
    output  wire                            AP_AXIMM_84_WREADY,
    output  wire [1:0]                      AP_AXIMM_84_BRESP,
    output  wire                            AP_AXIMM_84_BVALID,
    input wire                            AP_AXIMM_84_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_84_ARADDR,
    input wire [7:0]                      AP_AXIMM_84_ARLEN,
    input wire [2:0]                      AP_AXIMM_84_ARSIZE,
    input wire [1:0]                      AP_AXIMM_84_ARBURST,
    input wire [1:0]                      AP_AXIMM_84_ARLOCK,
    input wire [3:0]                      AP_AXIMM_84_ARCACHE,
    input wire [2:0]                      AP_AXIMM_84_ARPROT,
    input wire [3:0]                      AP_AXIMM_84_ARREGION,
    input wire [3:0]                      AP_AXIMM_84_ARQOS,
    input wire                            AP_AXIMM_84_ARVALID,
    output  wire                            AP_AXIMM_84_ARREADY,
    output  wire [M_AXIMM_84_DATA_WIDTH-1:0]   AP_AXIMM_84_RDATA,
    output  wire [1:0]                      AP_AXIMM_84_RRESP,
    output  wire                            AP_AXIMM_84_RLAST,
    output  wire                            AP_AXIMM_84_RVALID,
    input  wire                            AP_AXIMM_84_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_84_AWADDR,
    output wire [7:0]                      M_AXIMM_84_AWLEN,
    output wire [2:0]                      M_AXIMM_84_AWSIZE,
    output wire [1:0]                      M_AXIMM_84_AWBURST,
    output wire [1:0]                      M_AXIMM_84_AWLOCK,
    output wire [3:0]                      M_AXIMM_84_AWCACHE,
    output wire [2:0]                      M_AXIMM_84_AWPROT,
    output wire [3:0]                      M_AXIMM_84_AWREGION,
    output wire [3:0]                      M_AXIMM_84_AWQOS,
    output wire                            M_AXIMM_84_AWVALID,
    input  wire                            M_AXIMM_84_AWREADY,
    output wire [M_AXIMM_84_DATA_WIDTH-1:0]   M_AXIMM_84_WDATA,
    output wire [M_AXIMM_84_DATA_WIDTH/8-1:0] M_AXIMM_84_WSTRB,
    output wire                            M_AXIMM_84_WLAST,
    output wire                            M_AXIMM_84_WVALID,
    input  wire                            M_AXIMM_84_WREADY,
    input  wire [1:0]                      M_AXIMM_84_BRESP,
    input  wire                            M_AXIMM_84_BVALID,
    output wire                            M_AXIMM_84_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_84_ARADDR,
    output wire [7:0]                      M_AXIMM_84_ARLEN,
    output wire [2:0]                      M_AXIMM_84_ARSIZE,
    output wire [1:0]                      M_AXIMM_84_ARBURST,
    output wire [1:0]                      M_AXIMM_84_ARLOCK,
    output wire [3:0]                      M_AXIMM_84_ARCACHE,
    output wire [2:0]                      M_AXIMM_84_ARPROT,
    output wire [3:0]                      M_AXIMM_84_ARREGION,
    output wire [3:0]                      M_AXIMM_84_ARQOS,
    output wire                            M_AXIMM_84_ARVALID,
    input  wire                            M_AXIMM_84_ARREADY,
    input  wire [M_AXIMM_84_DATA_WIDTH-1:0]   M_AXIMM_84_RDATA,
    input  wire [1:0]                      M_AXIMM_84_RRESP,
    input  wire                            M_AXIMM_84_RLAST,
    input  wire                            M_AXIMM_84_RVALID,
    output wire                            M_AXIMM_84_RREADY,
    //AXI-MM pass-through interface 85
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_85_AWADDR,
    input wire [7:0]                      AP_AXIMM_85_AWLEN,
    input wire [2:0]                      AP_AXIMM_85_AWSIZE,
    input wire [1:0]                      AP_AXIMM_85_AWBURST,
    input wire [1:0]                      AP_AXIMM_85_AWLOCK,
    input wire [3:0]                      AP_AXIMM_85_AWCACHE,
    input wire [2:0]                      AP_AXIMM_85_AWPROT,
    input wire [3:0]                      AP_AXIMM_85_AWREGION,
    input wire [3:0]                      AP_AXIMM_85_AWQOS,
    input wire                            AP_AXIMM_85_AWVALID,
    output  wire                            AP_AXIMM_85_AWREADY,
    input wire [M_AXIMM_85_DATA_WIDTH-1:0]   AP_AXIMM_85_WDATA,
    input wire [M_AXIMM_85_DATA_WIDTH/8-1:0] AP_AXIMM_85_WSTRB,
    input wire                            AP_AXIMM_85_WLAST,
    input wire                            AP_AXIMM_85_WVALID,
    output  wire                            AP_AXIMM_85_WREADY,
    output  wire [1:0]                      AP_AXIMM_85_BRESP,
    output  wire                            AP_AXIMM_85_BVALID,
    input wire                            AP_AXIMM_85_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_85_ARADDR,
    input wire [7:0]                      AP_AXIMM_85_ARLEN,
    input wire [2:0]                      AP_AXIMM_85_ARSIZE,
    input wire [1:0]                      AP_AXIMM_85_ARBURST,
    input wire [1:0]                      AP_AXIMM_85_ARLOCK,
    input wire [3:0]                      AP_AXIMM_85_ARCACHE,
    input wire [2:0]                      AP_AXIMM_85_ARPROT,
    input wire [3:0]                      AP_AXIMM_85_ARREGION,
    input wire [3:0]                      AP_AXIMM_85_ARQOS,
    input wire                            AP_AXIMM_85_ARVALID,
    output  wire                            AP_AXIMM_85_ARREADY,
    output  wire [M_AXIMM_85_DATA_WIDTH-1:0]   AP_AXIMM_85_RDATA,
    output  wire [1:0]                      AP_AXIMM_85_RRESP,
    output  wire                            AP_AXIMM_85_RLAST,
    output  wire                            AP_AXIMM_85_RVALID,
    input  wire                            AP_AXIMM_85_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_85_AWADDR,
    output wire [7:0]                      M_AXIMM_85_AWLEN,
    output wire [2:0]                      M_AXIMM_85_AWSIZE,
    output wire [1:0]                      M_AXIMM_85_AWBURST,
    output wire [1:0]                      M_AXIMM_85_AWLOCK,
    output wire [3:0]                      M_AXIMM_85_AWCACHE,
    output wire [2:0]                      M_AXIMM_85_AWPROT,
    output wire [3:0]                      M_AXIMM_85_AWREGION,
    output wire [3:0]                      M_AXIMM_85_AWQOS,
    output wire                            M_AXIMM_85_AWVALID,
    input  wire                            M_AXIMM_85_AWREADY,
    output wire [M_AXIMM_85_DATA_WIDTH-1:0]   M_AXIMM_85_WDATA,
    output wire [M_AXIMM_85_DATA_WIDTH/8-1:0] M_AXIMM_85_WSTRB,
    output wire                            M_AXIMM_85_WLAST,
    output wire                            M_AXIMM_85_WVALID,
    input  wire                            M_AXIMM_85_WREADY,
    input  wire [1:0]                      M_AXIMM_85_BRESP,
    input  wire                            M_AXIMM_85_BVALID,
    output wire                            M_AXIMM_85_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_85_ARADDR,
    output wire [7:0]                      M_AXIMM_85_ARLEN,
    output wire [2:0]                      M_AXIMM_85_ARSIZE,
    output wire [1:0]                      M_AXIMM_85_ARBURST,
    output wire [1:0]                      M_AXIMM_85_ARLOCK,
    output wire [3:0]                      M_AXIMM_85_ARCACHE,
    output wire [2:0]                      M_AXIMM_85_ARPROT,
    output wire [3:0]                      M_AXIMM_85_ARREGION,
    output wire [3:0]                      M_AXIMM_85_ARQOS,
    output wire                            M_AXIMM_85_ARVALID,
    input  wire                            M_AXIMM_85_ARREADY,
    input  wire [M_AXIMM_85_DATA_WIDTH-1:0]   M_AXIMM_85_RDATA,
    input  wire [1:0]                      M_AXIMM_85_RRESP,
    input  wire                            M_AXIMM_85_RLAST,
    input  wire                            M_AXIMM_85_RVALID,
    output wire                            M_AXIMM_85_RREADY,
    //AXI-MM pass-through interface 86
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_86_AWADDR,
    input wire [7:0]                      AP_AXIMM_86_AWLEN,
    input wire [2:0]                      AP_AXIMM_86_AWSIZE,
    input wire [1:0]                      AP_AXIMM_86_AWBURST,
    input wire [1:0]                      AP_AXIMM_86_AWLOCK,
    input wire [3:0]                      AP_AXIMM_86_AWCACHE,
    input wire [2:0]                      AP_AXIMM_86_AWPROT,
    input wire [3:0]                      AP_AXIMM_86_AWREGION,
    input wire [3:0]                      AP_AXIMM_86_AWQOS,
    input wire                            AP_AXIMM_86_AWVALID,
    output  wire                            AP_AXIMM_86_AWREADY,
    input wire [M_AXIMM_86_DATA_WIDTH-1:0]   AP_AXIMM_86_WDATA,
    input wire [M_AXIMM_86_DATA_WIDTH/8-1:0] AP_AXIMM_86_WSTRB,
    input wire                            AP_AXIMM_86_WLAST,
    input wire                            AP_AXIMM_86_WVALID,
    output  wire                            AP_AXIMM_86_WREADY,
    output  wire [1:0]                      AP_AXIMM_86_BRESP,
    output  wire                            AP_AXIMM_86_BVALID,
    input wire                            AP_AXIMM_86_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_86_ARADDR,
    input wire [7:0]                      AP_AXIMM_86_ARLEN,
    input wire [2:0]                      AP_AXIMM_86_ARSIZE,
    input wire [1:0]                      AP_AXIMM_86_ARBURST,
    input wire [1:0]                      AP_AXIMM_86_ARLOCK,
    input wire [3:0]                      AP_AXIMM_86_ARCACHE,
    input wire [2:0]                      AP_AXIMM_86_ARPROT,
    input wire [3:0]                      AP_AXIMM_86_ARREGION,
    input wire [3:0]                      AP_AXIMM_86_ARQOS,
    input wire                            AP_AXIMM_86_ARVALID,
    output  wire                            AP_AXIMM_86_ARREADY,
    output  wire [M_AXIMM_86_DATA_WIDTH-1:0]   AP_AXIMM_86_RDATA,
    output  wire [1:0]                      AP_AXIMM_86_RRESP,
    output  wire                            AP_AXIMM_86_RLAST,
    output  wire                            AP_AXIMM_86_RVALID,
    input  wire                            AP_AXIMM_86_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_86_AWADDR,
    output wire [7:0]                      M_AXIMM_86_AWLEN,
    output wire [2:0]                      M_AXIMM_86_AWSIZE,
    output wire [1:0]                      M_AXIMM_86_AWBURST,
    output wire [1:0]                      M_AXIMM_86_AWLOCK,
    output wire [3:0]                      M_AXIMM_86_AWCACHE,
    output wire [2:0]                      M_AXIMM_86_AWPROT,
    output wire [3:0]                      M_AXIMM_86_AWREGION,
    output wire [3:0]                      M_AXIMM_86_AWQOS,
    output wire                            M_AXIMM_86_AWVALID,
    input  wire                            M_AXIMM_86_AWREADY,
    output wire [M_AXIMM_86_DATA_WIDTH-1:0]   M_AXIMM_86_WDATA,
    output wire [M_AXIMM_86_DATA_WIDTH/8-1:0] M_AXIMM_86_WSTRB,
    output wire                            M_AXIMM_86_WLAST,
    output wire                            M_AXIMM_86_WVALID,
    input  wire                            M_AXIMM_86_WREADY,
    input  wire [1:0]                      M_AXIMM_86_BRESP,
    input  wire                            M_AXIMM_86_BVALID,
    output wire                            M_AXIMM_86_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_86_ARADDR,
    output wire [7:0]                      M_AXIMM_86_ARLEN,
    output wire [2:0]                      M_AXIMM_86_ARSIZE,
    output wire [1:0]                      M_AXIMM_86_ARBURST,
    output wire [1:0]                      M_AXIMM_86_ARLOCK,
    output wire [3:0]                      M_AXIMM_86_ARCACHE,
    output wire [2:0]                      M_AXIMM_86_ARPROT,
    output wire [3:0]                      M_AXIMM_86_ARREGION,
    output wire [3:0]                      M_AXIMM_86_ARQOS,
    output wire                            M_AXIMM_86_ARVALID,
    input  wire                            M_AXIMM_86_ARREADY,
    input  wire [M_AXIMM_86_DATA_WIDTH-1:0]   M_AXIMM_86_RDATA,
    input  wire [1:0]                      M_AXIMM_86_RRESP,
    input  wire                            M_AXIMM_86_RLAST,
    input  wire                            M_AXIMM_86_RVALID,
    output wire                            M_AXIMM_86_RREADY,
    //AXI-MM pass-through interface 87
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_87_AWADDR,
    input wire [7:0]                      AP_AXIMM_87_AWLEN,
    input wire [2:0]                      AP_AXIMM_87_AWSIZE,
    input wire [1:0]                      AP_AXIMM_87_AWBURST,
    input wire [1:0]                      AP_AXIMM_87_AWLOCK,
    input wire [3:0]                      AP_AXIMM_87_AWCACHE,
    input wire [2:0]                      AP_AXIMM_87_AWPROT,
    input wire [3:0]                      AP_AXIMM_87_AWREGION,
    input wire [3:0]                      AP_AXIMM_87_AWQOS,
    input wire                            AP_AXIMM_87_AWVALID,
    output  wire                            AP_AXIMM_87_AWREADY,
    input wire [M_AXIMM_87_DATA_WIDTH-1:0]   AP_AXIMM_87_WDATA,
    input wire [M_AXIMM_87_DATA_WIDTH/8-1:0] AP_AXIMM_87_WSTRB,
    input wire                            AP_AXIMM_87_WLAST,
    input wire                            AP_AXIMM_87_WVALID,
    output  wire                            AP_AXIMM_87_WREADY,
    output  wire [1:0]                      AP_AXIMM_87_BRESP,
    output  wire                            AP_AXIMM_87_BVALID,
    input wire                            AP_AXIMM_87_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_87_ARADDR,
    input wire [7:0]                      AP_AXIMM_87_ARLEN,
    input wire [2:0]                      AP_AXIMM_87_ARSIZE,
    input wire [1:0]                      AP_AXIMM_87_ARBURST,
    input wire [1:0]                      AP_AXIMM_87_ARLOCK,
    input wire [3:0]                      AP_AXIMM_87_ARCACHE,
    input wire [2:0]                      AP_AXIMM_87_ARPROT,
    input wire [3:0]                      AP_AXIMM_87_ARREGION,
    input wire [3:0]                      AP_AXIMM_87_ARQOS,
    input wire                            AP_AXIMM_87_ARVALID,
    output  wire                            AP_AXIMM_87_ARREADY,
    output  wire [M_AXIMM_87_DATA_WIDTH-1:0]   AP_AXIMM_87_RDATA,
    output  wire [1:0]                      AP_AXIMM_87_RRESP,
    output  wire                            AP_AXIMM_87_RLAST,
    output  wire                            AP_AXIMM_87_RVALID,
    input  wire                            AP_AXIMM_87_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_87_AWADDR,
    output wire [7:0]                      M_AXIMM_87_AWLEN,
    output wire [2:0]                      M_AXIMM_87_AWSIZE,
    output wire [1:0]                      M_AXIMM_87_AWBURST,
    output wire [1:0]                      M_AXIMM_87_AWLOCK,
    output wire [3:0]                      M_AXIMM_87_AWCACHE,
    output wire [2:0]                      M_AXIMM_87_AWPROT,
    output wire [3:0]                      M_AXIMM_87_AWREGION,
    output wire [3:0]                      M_AXIMM_87_AWQOS,
    output wire                            M_AXIMM_87_AWVALID,
    input  wire                            M_AXIMM_87_AWREADY,
    output wire [M_AXIMM_87_DATA_WIDTH-1:0]   M_AXIMM_87_WDATA,
    output wire [M_AXIMM_87_DATA_WIDTH/8-1:0] M_AXIMM_87_WSTRB,
    output wire                            M_AXIMM_87_WLAST,
    output wire                            M_AXIMM_87_WVALID,
    input  wire                            M_AXIMM_87_WREADY,
    input  wire [1:0]                      M_AXIMM_87_BRESP,
    input  wire                            M_AXIMM_87_BVALID,
    output wire                            M_AXIMM_87_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_87_ARADDR,
    output wire [7:0]                      M_AXIMM_87_ARLEN,
    output wire [2:0]                      M_AXIMM_87_ARSIZE,
    output wire [1:0]                      M_AXIMM_87_ARBURST,
    output wire [1:0]                      M_AXIMM_87_ARLOCK,
    output wire [3:0]                      M_AXIMM_87_ARCACHE,
    output wire [2:0]                      M_AXIMM_87_ARPROT,
    output wire [3:0]                      M_AXIMM_87_ARREGION,
    output wire [3:0]                      M_AXIMM_87_ARQOS,
    output wire                            M_AXIMM_87_ARVALID,
    input  wire                            M_AXIMM_87_ARREADY,
    input  wire [M_AXIMM_87_DATA_WIDTH-1:0]   M_AXIMM_87_RDATA,
    input  wire [1:0]                      M_AXIMM_87_RRESP,
    input  wire                            M_AXIMM_87_RLAST,
    input  wire                            M_AXIMM_87_RVALID,
    output wire                            M_AXIMM_87_RREADY,
    //AXI-MM pass-through interface 88
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_88_AWADDR,
    input wire [7:0]                      AP_AXIMM_88_AWLEN,
    input wire [2:0]                      AP_AXIMM_88_AWSIZE,
    input wire [1:0]                      AP_AXIMM_88_AWBURST,
    input wire [1:0]                      AP_AXIMM_88_AWLOCK,
    input wire [3:0]                      AP_AXIMM_88_AWCACHE,
    input wire [2:0]                      AP_AXIMM_88_AWPROT,
    input wire [3:0]                      AP_AXIMM_88_AWREGION,
    input wire [3:0]                      AP_AXIMM_88_AWQOS,
    input wire                            AP_AXIMM_88_AWVALID,
    output  wire                            AP_AXIMM_88_AWREADY,
    input wire [M_AXIMM_88_DATA_WIDTH-1:0]   AP_AXIMM_88_WDATA,
    input wire [M_AXIMM_88_DATA_WIDTH/8-1:0] AP_AXIMM_88_WSTRB,
    input wire                            AP_AXIMM_88_WLAST,
    input wire                            AP_AXIMM_88_WVALID,
    output  wire                            AP_AXIMM_88_WREADY,
    output  wire [1:0]                      AP_AXIMM_88_BRESP,
    output  wire                            AP_AXIMM_88_BVALID,
    input wire                            AP_AXIMM_88_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_88_ARADDR,
    input wire [7:0]                      AP_AXIMM_88_ARLEN,
    input wire [2:0]                      AP_AXIMM_88_ARSIZE,
    input wire [1:0]                      AP_AXIMM_88_ARBURST,
    input wire [1:0]                      AP_AXIMM_88_ARLOCK,
    input wire [3:0]                      AP_AXIMM_88_ARCACHE,
    input wire [2:0]                      AP_AXIMM_88_ARPROT,
    input wire [3:0]                      AP_AXIMM_88_ARREGION,
    input wire [3:0]                      AP_AXIMM_88_ARQOS,
    input wire                            AP_AXIMM_88_ARVALID,
    output  wire                            AP_AXIMM_88_ARREADY,
    output  wire [M_AXIMM_88_DATA_WIDTH-1:0]   AP_AXIMM_88_RDATA,
    output  wire [1:0]                      AP_AXIMM_88_RRESP,
    output  wire                            AP_AXIMM_88_RLAST,
    output  wire                            AP_AXIMM_88_RVALID,
    input  wire                            AP_AXIMM_88_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_88_AWADDR,
    output wire [7:0]                      M_AXIMM_88_AWLEN,
    output wire [2:0]                      M_AXIMM_88_AWSIZE,
    output wire [1:0]                      M_AXIMM_88_AWBURST,
    output wire [1:0]                      M_AXIMM_88_AWLOCK,
    output wire [3:0]                      M_AXIMM_88_AWCACHE,
    output wire [2:0]                      M_AXIMM_88_AWPROT,
    output wire [3:0]                      M_AXIMM_88_AWREGION,
    output wire [3:0]                      M_AXIMM_88_AWQOS,
    output wire                            M_AXIMM_88_AWVALID,
    input  wire                            M_AXIMM_88_AWREADY,
    output wire [M_AXIMM_88_DATA_WIDTH-1:0]   M_AXIMM_88_WDATA,
    output wire [M_AXIMM_88_DATA_WIDTH/8-1:0] M_AXIMM_88_WSTRB,
    output wire                            M_AXIMM_88_WLAST,
    output wire                            M_AXIMM_88_WVALID,
    input  wire                            M_AXIMM_88_WREADY,
    input  wire [1:0]                      M_AXIMM_88_BRESP,
    input  wire                            M_AXIMM_88_BVALID,
    output wire                            M_AXIMM_88_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_88_ARADDR,
    output wire [7:0]                      M_AXIMM_88_ARLEN,
    output wire [2:0]                      M_AXIMM_88_ARSIZE,
    output wire [1:0]                      M_AXIMM_88_ARBURST,
    output wire [1:0]                      M_AXIMM_88_ARLOCK,
    output wire [3:0]                      M_AXIMM_88_ARCACHE,
    output wire [2:0]                      M_AXIMM_88_ARPROT,
    output wire [3:0]                      M_AXIMM_88_ARREGION,
    output wire [3:0]                      M_AXIMM_88_ARQOS,
    output wire                            M_AXIMM_88_ARVALID,
    input  wire                            M_AXIMM_88_ARREADY,
    input  wire [M_AXIMM_88_DATA_WIDTH-1:0]   M_AXIMM_88_RDATA,
    input  wire [1:0]                      M_AXIMM_88_RRESP,
    input  wire                            M_AXIMM_88_RLAST,
    input  wire                            M_AXIMM_88_RVALID,
    output wire                            M_AXIMM_88_RREADY,
    //AXI-MM pass-through interface 89
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_89_AWADDR,
    input wire [7:0]                      AP_AXIMM_89_AWLEN,
    input wire [2:0]                      AP_AXIMM_89_AWSIZE,
    input wire [1:0]                      AP_AXIMM_89_AWBURST,
    input wire [1:0]                      AP_AXIMM_89_AWLOCK,
    input wire [3:0]                      AP_AXIMM_89_AWCACHE,
    input wire [2:0]                      AP_AXIMM_89_AWPROT,
    input wire [3:0]                      AP_AXIMM_89_AWREGION,
    input wire [3:0]                      AP_AXIMM_89_AWQOS,
    input wire                            AP_AXIMM_89_AWVALID,
    output  wire                            AP_AXIMM_89_AWREADY,
    input wire [M_AXIMM_89_DATA_WIDTH-1:0]   AP_AXIMM_89_WDATA,
    input wire [M_AXIMM_89_DATA_WIDTH/8-1:0] AP_AXIMM_89_WSTRB,
    input wire                            AP_AXIMM_89_WLAST,
    input wire                            AP_AXIMM_89_WVALID,
    output  wire                            AP_AXIMM_89_WREADY,
    output  wire [1:0]                      AP_AXIMM_89_BRESP,
    output  wire                            AP_AXIMM_89_BVALID,
    input wire                            AP_AXIMM_89_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_89_ARADDR,
    input wire [7:0]                      AP_AXIMM_89_ARLEN,
    input wire [2:0]                      AP_AXIMM_89_ARSIZE,
    input wire [1:0]                      AP_AXIMM_89_ARBURST,
    input wire [1:0]                      AP_AXIMM_89_ARLOCK,
    input wire [3:0]                      AP_AXIMM_89_ARCACHE,
    input wire [2:0]                      AP_AXIMM_89_ARPROT,
    input wire [3:0]                      AP_AXIMM_89_ARREGION,
    input wire [3:0]                      AP_AXIMM_89_ARQOS,
    input wire                            AP_AXIMM_89_ARVALID,
    output  wire                            AP_AXIMM_89_ARREADY,
    output  wire [M_AXIMM_89_DATA_WIDTH-1:0]   AP_AXIMM_89_RDATA,
    output  wire [1:0]                      AP_AXIMM_89_RRESP,
    output  wire                            AP_AXIMM_89_RLAST,
    output  wire                            AP_AXIMM_89_RVALID,
    input  wire                            AP_AXIMM_89_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_89_AWADDR,
    output wire [7:0]                      M_AXIMM_89_AWLEN,
    output wire [2:0]                      M_AXIMM_89_AWSIZE,
    output wire [1:0]                      M_AXIMM_89_AWBURST,
    output wire [1:0]                      M_AXIMM_89_AWLOCK,
    output wire [3:0]                      M_AXIMM_89_AWCACHE,
    output wire [2:0]                      M_AXIMM_89_AWPROT,
    output wire [3:0]                      M_AXIMM_89_AWREGION,
    output wire [3:0]                      M_AXIMM_89_AWQOS,
    output wire                            M_AXIMM_89_AWVALID,
    input  wire                            M_AXIMM_89_AWREADY,
    output wire [M_AXIMM_89_DATA_WIDTH-1:0]   M_AXIMM_89_WDATA,
    output wire [M_AXIMM_89_DATA_WIDTH/8-1:0] M_AXIMM_89_WSTRB,
    output wire                            M_AXIMM_89_WLAST,
    output wire                            M_AXIMM_89_WVALID,
    input  wire                            M_AXIMM_89_WREADY,
    input  wire [1:0]                      M_AXIMM_89_BRESP,
    input  wire                            M_AXIMM_89_BVALID,
    output wire                            M_AXIMM_89_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_89_ARADDR,
    output wire [7:0]                      M_AXIMM_89_ARLEN,
    output wire [2:0]                      M_AXIMM_89_ARSIZE,
    output wire [1:0]                      M_AXIMM_89_ARBURST,
    output wire [1:0]                      M_AXIMM_89_ARLOCK,
    output wire [3:0]                      M_AXIMM_89_ARCACHE,
    output wire [2:0]                      M_AXIMM_89_ARPROT,
    output wire [3:0]                      M_AXIMM_89_ARREGION,
    output wire [3:0]                      M_AXIMM_89_ARQOS,
    output wire                            M_AXIMM_89_ARVALID,
    input  wire                            M_AXIMM_89_ARREADY,
    input  wire [M_AXIMM_89_DATA_WIDTH-1:0]   M_AXIMM_89_RDATA,
    input  wire [1:0]                      M_AXIMM_89_RRESP,
    input  wire                            M_AXIMM_89_RLAST,
    input  wire                            M_AXIMM_89_RVALID,
    output wire                            M_AXIMM_89_RREADY,
    //AXI-MM pass-through interface 90
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_90_AWADDR,
    input wire [7:0]                      AP_AXIMM_90_AWLEN,
    input wire [2:0]                      AP_AXIMM_90_AWSIZE,
    input wire [1:0]                      AP_AXIMM_90_AWBURST,
    input wire [1:0]                      AP_AXIMM_90_AWLOCK,
    input wire [3:0]                      AP_AXIMM_90_AWCACHE,
    input wire [2:0]                      AP_AXIMM_90_AWPROT,
    input wire [3:0]                      AP_AXIMM_90_AWREGION,
    input wire [3:0]                      AP_AXIMM_90_AWQOS,
    input wire                            AP_AXIMM_90_AWVALID,
    output  wire                            AP_AXIMM_90_AWREADY,
    input wire [M_AXIMM_90_DATA_WIDTH-1:0]   AP_AXIMM_90_WDATA,
    input wire [M_AXIMM_90_DATA_WIDTH/8-1:0] AP_AXIMM_90_WSTRB,
    input wire                            AP_AXIMM_90_WLAST,
    input wire                            AP_AXIMM_90_WVALID,
    output  wire                            AP_AXIMM_90_WREADY,
    output  wire [1:0]                      AP_AXIMM_90_BRESP,
    output  wire                            AP_AXIMM_90_BVALID,
    input wire                            AP_AXIMM_90_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_90_ARADDR,
    input wire [7:0]                      AP_AXIMM_90_ARLEN,
    input wire [2:0]                      AP_AXIMM_90_ARSIZE,
    input wire [1:0]                      AP_AXIMM_90_ARBURST,
    input wire [1:0]                      AP_AXIMM_90_ARLOCK,
    input wire [3:0]                      AP_AXIMM_90_ARCACHE,
    input wire [2:0]                      AP_AXIMM_90_ARPROT,
    input wire [3:0]                      AP_AXIMM_90_ARREGION,
    input wire [3:0]                      AP_AXIMM_90_ARQOS,
    input wire                            AP_AXIMM_90_ARVALID,
    output  wire                            AP_AXIMM_90_ARREADY,
    output  wire [M_AXIMM_90_DATA_WIDTH-1:0]   AP_AXIMM_90_RDATA,
    output  wire [1:0]                      AP_AXIMM_90_RRESP,
    output  wire                            AP_AXIMM_90_RLAST,
    output  wire                            AP_AXIMM_90_RVALID,
    input  wire                            AP_AXIMM_90_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_90_AWADDR,
    output wire [7:0]                      M_AXIMM_90_AWLEN,
    output wire [2:0]                      M_AXIMM_90_AWSIZE,
    output wire [1:0]                      M_AXIMM_90_AWBURST,
    output wire [1:0]                      M_AXIMM_90_AWLOCK,
    output wire [3:0]                      M_AXIMM_90_AWCACHE,
    output wire [2:0]                      M_AXIMM_90_AWPROT,
    output wire [3:0]                      M_AXIMM_90_AWREGION,
    output wire [3:0]                      M_AXIMM_90_AWQOS,
    output wire                            M_AXIMM_90_AWVALID,
    input  wire                            M_AXIMM_90_AWREADY,
    output wire [M_AXIMM_90_DATA_WIDTH-1:0]   M_AXIMM_90_WDATA,
    output wire [M_AXIMM_90_DATA_WIDTH/8-1:0] M_AXIMM_90_WSTRB,
    output wire                            M_AXIMM_90_WLAST,
    output wire                            M_AXIMM_90_WVALID,
    input  wire                            M_AXIMM_90_WREADY,
    input  wire [1:0]                      M_AXIMM_90_BRESP,
    input  wire                            M_AXIMM_90_BVALID,
    output wire                            M_AXIMM_90_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_90_ARADDR,
    output wire [7:0]                      M_AXIMM_90_ARLEN,
    output wire [2:0]                      M_AXIMM_90_ARSIZE,
    output wire [1:0]                      M_AXIMM_90_ARBURST,
    output wire [1:0]                      M_AXIMM_90_ARLOCK,
    output wire [3:0]                      M_AXIMM_90_ARCACHE,
    output wire [2:0]                      M_AXIMM_90_ARPROT,
    output wire [3:0]                      M_AXIMM_90_ARREGION,
    output wire [3:0]                      M_AXIMM_90_ARQOS,
    output wire                            M_AXIMM_90_ARVALID,
    input  wire                            M_AXIMM_90_ARREADY,
    input  wire [M_AXIMM_90_DATA_WIDTH-1:0]   M_AXIMM_90_RDATA,
    input  wire [1:0]                      M_AXIMM_90_RRESP,
    input  wire                            M_AXIMM_90_RLAST,
    input  wire                            M_AXIMM_90_RVALID,
    output wire                            M_AXIMM_90_RREADY,
    //AXI-MM pass-through interface 91
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_91_AWADDR,
    input wire [7:0]                      AP_AXIMM_91_AWLEN,
    input wire [2:0]                      AP_AXIMM_91_AWSIZE,
    input wire [1:0]                      AP_AXIMM_91_AWBURST,
    input wire [1:0]                      AP_AXIMM_91_AWLOCK,
    input wire [3:0]                      AP_AXIMM_91_AWCACHE,
    input wire [2:0]                      AP_AXIMM_91_AWPROT,
    input wire [3:0]                      AP_AXIMM_91_AWREGION,
    input wire [3:0]                      AP_AXIMM_91_AWQOS,
    input wire                            AP_AXIMM_91_AWVALID,
    output  wire                            AP_AXIMM_91_AWREADY,
    input wire [M_AXIMM_91_DATA_WIDTH-1:0]   AP_AXIMM_91_WDATA,
    input wire [M_AXIMM_91_DATA_WIDTH/8-1:0] AP_AXIMM_91_WSTRB,
    input wire                            AP_AXIMM_91_WLAST,
    input wire                            AP_AXIMM_91_WVALID,
    output  wire                            AP_AXIMM_91_WREADY,
    output  wire [1:0]                      AP_AXIMM_91_BRESP,
    output  wire                            AP_AXIMM_91_BVALID,
    input wire                            AP_AXIMM_91_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_91_ARADDR,
    input wire [7:0]                      AP_AXIMM_91_ARLEN,
    input wire [2:0]                      AP_AXIMM_91_ARSIZE,
    input wire [1:0]                      AP_AXIMM_91_ARBURST,
    input wire [1:0]                      AP_AXIMM_91_ARLOCK,
    input wire [3:0]                      AP_AXIMM_91_ARCACHE,
    input wire [2:0]                      AP_AXIMM_91_ARPROT,
    input wire [3:0]                      AP_AXIMM_91_ARREGION,
    input wire [3:0]                      AP_AXIMM_91_ARQOS,
    input wire                            AP_AXIMM_91_ARVALID,
    output  wire                            AP_AXIMM_91_ARREADY,
    output  wire [M_AXIMM_91_DATA_WIDTH-1:0]   AP_AXIMM_91_RDATA,
    output  wire [1:0]                      AP_AXIMM_91_RRESP,
    output  wire                            AP_AXIMM_91_RLAST,
    output  wire                            AP_AXIMM_91_RVALID,
    input  wire                            AP_AXIMM_91_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_91_AWADDR,
    output wire [7:0]                      M_AXIMM_91_AWLEN,
    output wire [2:0]                      M_AXIMM_91_AWSIZE,
    output wire [1:0]                      M_AXIMM_91_AWBURST,
    output wire [1:0]                      M_AXIMM_91_AWLOCK,
    output wire [3:0]                      M_AXIMM_91_AWCACHE,
    output wire [2:0]                      M_AXIMM_91_AWPROT,
    output wire [3:0]                      M_AXIMM_91_AWREGION,
    output wire [3:0]                      M_AXIMM_91_AWQOS,
    output wire                            M_AXIMM_91_AWVALID,
    input  wire                            M_AXIMM_91_AWREADY,
    output wire [M_AXIMM_91_DATA_WIDTH-1:0]   M_AXIMM_91_WDATA,
    output wire [M_AXIMM_91_DATA_WIDTH/8-1:0] M_AXIMM_91_WSTRB,
    output wire                            M_AXIMM_91_WLAST,
    output wire                            M_AXIMM_91_WVALID,
    input  wire                            M_AXIMM_91_WREADY,
    input  wire [1:0]                      M_AXIMM_91_BRESP,
    input  wire                            M_AXIMM_91_BVALID,
    output wire                            M_AXIMM_91_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_91_ARADDR,
    output wire [7:0]                      M_AXIMM_91_ARLEN,
    output wire [2:0]                      M_AXIMM_91_ARSIZE,
    output wire [1:0]                      M_AXIMM_91_ARBURST,
    output wire [1:0]                      M_AXIMM_91_ARLOCK,
    output wire [3:0]                      M_AXIMM_91_ARCACHE,
    output wire [2:0]                      M_AXIMM_91_ARPROT,
    output wire [3:0]                      M_AXIMM_91_ARREGION,
    output wire [3:0]                      M_AXIMM_91_ARQOS,
    output wire                            M_AXIMM_91_ARVALID,
    input  wire                            M_AXIMM_91_ARREADY,
    input  wire [M_AXIMM_91_DATA_WIDTH-1:0]   M_AXIMM_91_RDATA,
    input  wire [1:0]                      M_AXIMM_91_RRESP,
    input  wire                            M_AXIMM_91_RLAST,
    input  wire                            M_AXIMM_91_RVALID,
    output wire                            M_AXIMM_91_RREADY,
    //AXI-MM pass-through interface 92
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_92_AWADDR,
    input wire [7:0]                      AP_AXIMM_92_AWLEN,
    input wire [2:0]                      AP_AXIMM_92_AWSIZE,
    input wire [1:0]                      AP_AXIMM_92_AWBURST,
    input wire [1:0]                      AP_AXIMM_92_AWLOCK,
    input wire [3:0]                      AP_AXIMM_92_AWCACHE,
    input wire [2:0]                      AP_AXIMM_92_AWPROT,
    input wire [3:0]                      AP_AXIMM_92_AWREGION,
    input wire [3:0]                      AP_AXIMM_92_AWQOS,
    input wire                            AP_AXIMM_92_AWVALID,
    output  wire                            AP_AXIMM_92_AWREADY,
    input wire [M_AXIMM_92_DATA_WIDTH-1:0]   AP_AXIMM_92_WDATA,
    input wire [M_AXIMM_92_DATA_WIDTH/8-1:0] AP_AXIMM_92_WSTRB,
    input wire                            AP_AXIMM_92_WLAST,
    input wire                            AP_AXIMM_92_WVALID,
    output  wire                            AP_AXIMM_92_WREADY,
    output  wire [1:0]                      AP_AXIMM_92_BRESP,
    output  wire                            AP_AXIMM_92_BVALID,
    input wire                            AP_AXIMM_92_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_92_ARADDR,
    input wire [7:0]                      AP_AXIMM_92_ARLEN,
    input wire [2:0]                      AP_AXIMM_92_ARSIZE,
    input wire [1:0]                      AP_AXIMM_92_ARBURST,
    input wire [1:0]                      AP_AXIMM_92_ARLOCK,
    input wire [3:0]                      AP_AXIMM_92_ARCACHE,
    input wire [2:0]                      AP_AXIMM_92_ARPROT,
    input wire [3:0]                      AP_AXIMM_92_ARREGION,
    input wire [3:0]                      AP_AXIMM_92_ARQOS,
    input wire                            AP_AXIMM_92_ARVALID,
    output  wire                            AP_AXIMM_92_ARREADY,
    output  wire [M_AXIMM_92_DATA_WIDTH-1:0]   AP_AXIMM_92_RDATA,
    output  wire [1:0]                      AP_AXIMM_92_RRESP,
    output  wire                            AP_AXIMM_92_RLAST,
    output  wire                            AP_AXIMM_92_RVALID,
    input  wire                            AP_AXIMM_92_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_92_AWADDR,
    output wire [7:0]                      M_AXIMM_92_AWLEN,
    output wire [2:0]                      M_AXIMM_92_AWSIZE,
    output wire [1:0]                      M_AXIMM_92_AWBURST,
    output wire [1:0]                      M_AXIMM_92_AWLOCK,
    output wire [3:0]                      M_AXIMM_92_AWCACHE,
    output wire [2:0]                      M_AXIMM_92_AWPROT,
    output wire [3:0]                      M_AXIMM_92_AWREGION,
    output wire [3:0]                      M_AXIMM_92_AWQOS,
    output wire                            M_AXIMM_92_AWVALID,
    input  wire                            M_AXIMM_92_AWREADY,
    output wire [M_AXIMM_92_DATA_WIDTH-1:0]   M_AXIMM_92_WDATA,
    output wire [M_AXIMM_92_DATA_WIDTH/8-1:0] M_AXIMM_92_WSTRB,
    output wire                            M_AXIMM_92_WLAST,
    output wire                            M_AXIMM_92_WVALID,
    input  wire                            M_AXIMM_92_WREADY,
    input  wire [1:0]                      M_AXIMM_92_BRESP,
    input  wire                            M_AXIMM_92_BVALID,
    output wire                            M_AXIMM_92_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_92_ARADDR,
    output wire [7:0]                      M_AXIMM_92_ARLEN,
    output wire [2:0]                      M_AXIMM_92_ARSIZE,
    output wire [1:0]                      M_AXIMM_92_ARBURST,
    output wire [1:0]                      M_AXIMM_92_ARLOCK,
    output wire [3:0]                      M_AXIMM_92_ARCACHE,
    output wire [2:0]                      M_AXIMM_92_ARPROT,
    output wire [3:0]                      M_AXIMM_92_ARREGION,
    output wire [3:0]                      M_AXIMM_92_ARQOS,
    output wire                            M_AXIMM_92_ARVALID,
    input  wire                            M_AXIMM_92_ARREADY,
    input  wire [M_AXIMM_92_DATA_WIDTH-1:0]   M_AXIMM_92_RDATA,
    input  wire [1:0]                      M_AXIMM_92_RRESP,
    input  wire                            M_AXIMM_92_RLAST,
    input  wire                            M_AXIMM_92_RVALID,
    output wire                            M_AXIMM_92_RREADY,
    //AXI-MM pass-through interface 93
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_93_AWADDR,
    input wire [7:0]                      AP_AXIMM_93_AWLEN,
    input wire [2:0]                      AP_AXIMM_93_AWSIZE,
    input wire [1:0]                      AP_AXIMM_93_AWBURST,
    input wire [1:0]                      AP_AXIMM_93_AWLOCK,
    input wire [3:0]                      AP_AXIMM_93_AWCACHE,
    input wire [2:0]                      AP_AXIMM_93_AWPROT,
    input wire [3:0]                      AP_AXIMM_93_AWREGION,
    input wire [3:0]                      AP_AXIMM_93_AWQOS,
    input wire                            AP_AXIMM_93_AWVALID,
    output  wire                            AP_AXIMM_93_AWREADY,
    input wire [M_AXIMM_93_DATA_WIDTH-1:0]   AP_AXIMM_93_WDATA,
    input wire [M_AXIMM_93_DATA_WIDTH/8-1:0] AP_AXIMM_93_WSTRB,
    input wire                            AP_AXIMM_93_WLAST,
    input wire                            AP_AXIMM_93_WVALID,
    output  wire                            AP_AXIMM_93_WREADY,
    output  wire [1:0]                      AP_AXIMM_93_BRESP,
    output  wire                            AP_AXIMM_93_BVALID,
    input wire                            AP_AXIMM_93_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_93_ARADDR,
    input wire [7:0]                      AP_AXIMM_93_ARLEN,
    input wire [2:0]                      AP_AXIMM_93_ARSIZE,
    input wire [1:0]                      AP_AXIMM_93_ARBURST,
    input wire [1:0]                      AP_AXIMM_93_ARLOCK,
    input wire [3:0]                      AP_AXIMM_93_ARCACHE,
    input wire [2:0]                      AP_AXIMM_93_ARPROT,
    input wire [3:0]                      AP_AXIMM_93_ARREGION,
    input wire [3:0]                      AP_AXIMM_93_ARQOS,
    input wire                            AP_AXIMM_93_ARVALID,
    output  wire                            AP_AXIMM_93_ARREADY,
    output  wire [M_AXIMM_93_DATA_WIDTH-1:0]   AP_AXIMM_93_RDATA,
    output  wire [1:0]                      AP_AXIMM_93_RRESP,
    output  wire                            AP_AXIMM_93_RLAST,
    output  wire                            AP_AXIMM_93_RVALID,
    input  wire                            AP_AXIMM_93_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_93_AWADDR,
    output wire [7:0]                      M_AXIMM_93_AWLEN,
    output wire [2:0]                      M_AXIMM_93_AWSIZE,
    output wire [1:0]                      M_AXIMM_93_AWBURST,
    output wire [1:0]                      M_AXIMM_93_AWLOCK,
    output wire [3:0]                      M_AXIMM_93_AWCACHE,
    output wire [2:0]                      M_AXIMM_93_AWPROT,
    output wire [3:0]                      M_AXIMM_93_AWREGION,
    output wire [3:0]                      M_AXIMM_93_AWQOS,
    output wire                            M_AXIMM_93_AWVALID,
    input  wire                            M_AXIMM_93_AWREADY,
    output wire [M_AXIMM_93_DATA_WIDTH-1:0]   M_AXIMM_93_WDATA,
    output wire [M_AXIMM_93_DATA_WIDTH/8-1:0] M_AXIMM_93_WSTRB,
    output wire                            M_AXIMM_93_WLAST,
    output wire                            M_AXIMM_93_WVALID,
    input  wire                            M_AXIMM_93_WREADY,
    input  wire [1:0]                      M_AXIMM_93_BRESP,
    input  wire                            M_AXIMM_93_BVALID,
    output wire                            M_AXIMM_93_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_93_ARADDR,
    output wire [7:0]                      M_AXIMM_93_ARLEN,
    output wire [2:0]                      M_AXIMM_93_ARSIZE,
    output wire [1:0]                      M_AXIMM_93_ARBURST,
    output wire [1:0]                      M_AXIMM_93_ARLOCK,
    output wire [3:0]                      M_AXIMM_93_ARCACHE,
    output wire [2:0]                      M_AXIMM_93_ARPROT,
    output wire [3:0]                      M_AXIMM_93_ARREGION,
    output wire [3:0]                      M_AXIMM_93_ARQOS,
    output wire                            M_AXIMM_93_ARVALID,
    input  wire                            M_AXIMM_93_ARREADY,
    input  wire [M_AXIMM_93_DATA_WIDTH-1:0]   M_AXIMM_93_RDATA,
    input  wire [1:0]                      M_AXIMM_93_RRESP,
    input  wire                            M_AXIMM_93_RLAST,
    input  wire                            M_AXIMM_93_RVALID,
    output wire                            M_AXIMM_93_RREADY,
    //AXI-MM pass-through interface 94
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_94_AWADDR,
    input wire [7:0]                      AP_AXIMM_94_AWLEN,
    input wire [2:0]                      AP_AXIMM_94_AWSIZE,
    input wire [1:0]                      AP_AXIMM_94_AWBURST,
    input wire [1:0]                      AP_AXIMM_94_AWLOCK,
    input wire [3:0]                      AP_AXIMM_94_AWCACHE,
    input wire [2:0]                      AP_AXIMM_94_AWPROT,
    input wire [3:0]                      AP_AXIMM_94_AWREGION,
    input wire [3:0]                      AP_AXIMM_94_AWQOS,
    input wire                            AP_AXIMM_94_AWVALID,
    output  wire                            AP_AXIMM_94_AWREADY,
    input wire [M_AXIMM_94_DATA_WIDTH-1:0]   AP_AXIMM_94_WDATA,
    input wire [M_AXIMM_94_DATA_WIDTH/8-1:0] AP_AXIMM_94_WSTRB,
    input wire                            AP_AXIMM_94_WLAST,
    input wire                            AP_AXIMM_94_WVALID,
    output  wire                            AP_AXIMM_94_WREADY,
    output  wire [1:0]                      AP_AXIMM_94_BRESP,
    output  wire                            AP_AXIMM_94_BVALID,
    input wire                            AP_AXIMM_94_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_94_ARADDR,
    input wire [7:0]                      AP_AXIMM_94_ARLEN,
    input wire [2:0]                      AP_AXIMM_94_ARSIZE,
    input wire [1:0]                      AP_AXIMM_94_ARBURST,
    input wire [1:0]                      AP_AXIMM_94_ARLOCK,
    input wire [3:0]                      AP_AXIMM_94_ARCACHE,
    input wire [2:0]                      AP_AXIMM_94_ARPROT,
    input wire [3:0]                      AP_AXIMM_94_ARREGION,
    input wire [3:0]                      AP_AXIMM_94_ARQOS,
    input wire                            AP_AXIMM_94_ARVALID,
    output  wire                            AP_AXIMM_94_ARREADY,
    output  wire [M_AXIMM_94_DATA_WIDTH-1:0]   AP_AXIMM_94_RDATA,
    output  wire [1:0]                      AP_AXIMM_94_RRESP,
    output  wire                            AP_AXIMM_94_RLAST,
    output  wire                            AP_AXIMM_94_RVALID,
    input  wire                            AP_AXIMM_94_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_94_AWADDR,
    output wire [7:0]                      M_AXIMM_94_AWLEN,
    output wire [2:0]                      M_AXIMM_94_AWSIZE,
    output wire [1:0]                      M_AXIMM_94_AWBURST,
    output wire [1:0]                      M_AXIMM_94_AWLOCK,
    output wire [3:0]                      M_AXIMM_94_AWCACHE,
    output wire [2:0]                      M_AXIMM_94_AWPROT,
    output wire [3:0]                      M_AXIMM_94_AWREGION,
    output wire [3:0]                      M_AXIMM_94_AWQOS,
    output wire                            M_AXIMM_94_AWVALID,
    input  wire                            M_AXIMM_94_AWREADY,
    output wire [M_AXIMM_94_DATA_WIDTH-1:0]   M_AXIMM_94_WDATA,
    output wire [M_AXIMM_94_DATA_WIDTH/8-1:0] M_AXIMM_94_WSTRB,
    output wire                            M_AXIMM_94_WLAST,
    output wire                            M_AXIMM_94_WVALID,
    input  wire                            M_AXIMM_94_WREADY,
    input  wire [1:0]                      M_AXIMM_94_BRESP,
    input  wire                            M_AXIMM_94_BVALID,
    output wire                            M_AXIMM_94_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_94_ARADDR,
    output wire [7:0]                      M_AXIMM_94_ARLEN,
    output wire [2:0]                      M_AXIMM_94_ARSIZE,
    output wire [1:0]                      M_AXIMM_94_ARBURST,
    output wire [1:0]                      M_AXIMM_94_ARLOCK,
    output wire [3:0]                      M_AXIMM_94_ARCACHE,
    output wire [2:0]                      M_AXIMM_94_ARPROT,
    output wire [3:0]                      M_AXIMM_94_ARREGION,
    output wire [3:0]                      M_AXIMM_94_ARQOS,
    output wire                            M_AXIMM_94_ARVALID,
    input  wire                            M_AXIMM_94_ARREADY,
    input  wire [M_AXIMM_94_DATA_WIDTH-1:0]   M_AXIMM_94_RDATA,
    input  wire [1:0]                      M_AXIMM_94_RRESP,
    input  wire                            M_AXIMM_94_RLAST,
    input  wire                            M_AXIMM_94_RVALID,
    output wire                            M_AXIMM_94_RREADY,
    //AXI-MM pass-through interface 95
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_95_AWADDR,
    input wire [7:0]                      AP_AXIMM_95_AWLEN,
    input wire [2:0]                      AP_AXIMM_95_AWSIZE,
    input wire [1:0]                      AP_AXIMM_95_AWBURST,
    input wire [1:0]                      AP_AXIMM_95_AWLOCK,
    input wire [3:0]                      AP_AXIMM_95_AWCACHE,
    input wire [2:0]                      AP_AXIMM_95_AWPROT,
    input wire [3:0]                      AP_AXIMM_95_AWREGION,
    input wire [3:0]                      AP_AXIMM_95_AWQOS,
    input wire                            AP_AXIMM_95_AWVALID,
    output  wire                            AP_AXIMM_95_AWREADY,
    input wire [M_AXIMM_95_DATA_WIDTH-1:0]   AP_AXIMM_95_WDATA,
    input wire [M_AXIMM_95_DATA_WIDTH/8-1:0] AP_AXIMM_95_WSTRB,
    input wire                            AP_AXIMM_95_WLAST,
    input wire                            AP_AXIMM_95_WVALID,
    output  wire                            AP_AXIMM_95_WREADY,
    output  wire [1:0]                      AP_AXIMM_95_BRESP,
    output  wire                            AP_AXIMM_95_BVALID,
    input wire                            AP_AXIMM_95_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_95_ARADDR,
    input wire [7:0]                      AP_AXIMM_95_ARLEN,
    input wire [2:0]                      AP_AXIMM_95_ARSIZE,
    input wire [1:0]                      AP_AXIMM_95_ARBURST,
    input wire [1:0]                      AP_AXIMM_95_ARLOCK,
    input wire [3:0]                      AP_AXIMM_95_ARCACHE,
    input wire [2:0]                      AP_AXIMM_95_ARPROT,
    input wire [3:0]                      AP_AXIMM_95_ARREGION,
    input wire [3:0]                      AP_AXIMM_95_ARQOS,
    input wire                            AP_AXIMM_95_ARVALID,
    output  wire                            AP_AXIMM_95_ARREADY,
    output  wire [M_AXIMM_95_DATA_WIDTH-1:0]   AP_AXIMM_95_RDATA,
    output  wire [1:0]                      AP_AXIMM_95_RRESP,
    output  wire                            AP_AXIMM_95_RLAST,
    output  wire                            AP_AXIMM_95_RVALID,
    input  wire                            AP_AXIMM_95_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_95_AWADDR,
    output wire [7:0]                      M_AXIMM_95_AWLEN,
    output wire [2:0]                      M_AXIMM_95_AWSIZE,
    output wire [1:0]                      M_AXIMM_95_AWBURST,
    output wire [1:0]                      M_AXIMM_95_AWLOCK,
    output wire [3:0]                      M_AXIMM_95_AWCACHE,
    output wire [2:0]                      M_AXIMM_95_AWPROT,
    output wire [3:0]                      M_AXIMM_95_AWREGION,
    output wire [3:0]                      M_AXIMM_95_AWQOS,
    output wire                            M_AXIMM_95_AWVALID,
    input  wire                            M_AXIMM_95_AWREADY,
    output wire [M_AXIMM_95_DATA_WIDTH-1:0]   M_AXIMM_95_WDATA,
    output wire [M_AXIMM_95_DATA_WIDTH/8-1:0] M_AXIMM_95_WSTRB,
    output wire                            M_AXIMM_95_WLAST,
    output wire                            M_AXIMM_95_WVALID,
    input  wire                            M_AXIMM_95_WREADY,
    input  wire [1:0]                      M_AXIMM_95_BRESP,
    input  wire                            M_AXIMM_95_BVALID,
    output wire                            M_AXIMM_95_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_95_ARADDR,
    output wire [7:0]                      M_AXIMM_95_ARLEN,
    output wire [2:0]                      M_AXIMM_95_ARSIZE,
    output wire [1:0]                      M_AXIMM_95_ARBURST,
    output wire [1:0]                      M_AXIMM_95_ARLOCK,
    output wire [3:0]                      M_AXIMM_95_ARCACHE,
    output wire [2:0]                      M_AXIMM_95_ARPROT,
    output wire [3:0]                      M_AXIMM_95_ARREGION,
    output wire [3:0]                      M_AXIMM_95_ARQOS,
    output wire                            M_AXIMM_95_ARVALID,
    input  wire                            M_AXIMM_95_ARREADY,
    input  wire [M_AXIMM_95_DATA_WIDTH-1:0]   M_AXIMM_95_RDATA,
    input  wire [1:0]                      M_AXIMM_95_RRESP,
    input  wire                            M_AXIMM_95_RLAST,
    input  wire                            M_AXIMM_95_RVALID,
    output wire                            M_AXIMM_95_RREADY,
    //AXI-MM pass-through interface 96
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_96_AWADDR,
    input wire [7:0]                      AP_AXIMM_96_AWLEN,
    input wire [2:0]                      AP_AXIMM_96_AWSIZE,
    input wire [1:0]                      AP_AXIMM_96_AWBURST,
    input wire [1:0]                      AP_AXIMM_96_AWLOCK,
    input wire [3:0]                      AP_AXIMM_96_AWCACHE,
    input wire [2:0]                      AP_AXIMM_96_AWPROT,
    input wire [3:0]                      AP_AXIMM_96_AWREGION,
    input wire [3:0]                      AP_AXIMM_96_AWQOS,
    input wire                            AP_AXIMM_96_AWVALID,
    output  wire                            AP_AXIMM_96_AWREADY,
    input wire [M_AXIMM_96_DATA_WIDTH-1:0]   AP_AXIMM_96_WDATA,
    input wire [M_AXIMM_96_DATA_WIDTH/8-1:0] AP_AXIMM_96_WSTRB,
    input wire                            AP_AXIMM_96_WLAST,
    input wire                            AP_AXIMM_96_WVALID,
    output  wire                            AP_AXIMM_96_WREADY,
    output  wire [1:0]                      AP_AXIMM_96_BRESP,
    output  wire                            AP_AXIMM_96_BVALID,
    input wire                            AP_AXIMM_96_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_96_ARADDR,
    input wire [7:0]                      AP_AXIMM_96_ARLEN,
    input wire [2:0]                      AP_AXIMM_96_ARSIZE,
    input wire [1:0]                      AP_AXIMM_96_ARBURST,
    input wire [1:0]                      AP_AXIMM_96_ARLOCK,
    input wire [3:0]                      AP_AXIMM_96_ARCACHE,
    input wire [2:0]                      AP_AXIMM_96_ARPROT,
    input wire [3:0]                      AP_AXIMM_96_ARREGION,
    input wire [3:0]                      AP_AXIMM_96_ARQOS,
    input wire                            AP_AXIMM_96_ARVALID,
    output  wire                            AP_AXIMM_96_ARREADY,
    output  wire [M_AXIMM_96_DATA_WIDTH-1:0]   AP_AXIMM_96_RDATA,
    output  wire [1:0]                      AP_AXIMM_96_RRESP,
    output  wire                            AP_AXIMM_96_RLAST,
    output  wire                            AP_AXIMM_96_RVALID,
    input  wire                            AP_AXIMM_96_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_96_AWADDR,
    output wire [7:0]                      M_AXIMM_96_AWLEN,
    output wire [2:0]                      M_AXIMM_96_AWSIZE,
    output wire [1:0]                      M_AXIMM_96_AWBURST,
    output wire [1:0]                      M_AXIMM_96_AWLOCK,
    output wire [3:0]                      M_AXIMM_96_AWCACHE,
    output wire [2:0]                      M_AXIMM_96_AWPROT,
    output wire [3:0]                      M_AXIMM_96_AWREGION,
    output wire [3:0]                      M_AXIMM_96_AWQOS,
    output wire                            M_AXIMM_96_AWVALID,
    input  wire                            M_AXIMM_96_AWREADY,
    output wire [M_AXIMM_96_DATA_WIDTH-1:0]   M_AXIMM_96_WDATA,
    output wire [M_AXIMM_96_DATA_WIDTH/8-1:0] M_AXIMM_96_WSTRB,
    output wire                            M_AXIMM_96_WLAST,
    output wire                            M_AXIMM_96_WVALID,
    input  wire                            M_AXIMM_96_WREADY,
    input  wire [1:0]                      M_AXIMM_96_BRESP,
    input  wire                            M_AXIMM_96_BVALID,
    output wire                            M_AXIMM_96_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_96_ARADDR,
    output wire [7:0]                      M_AXIMM_96_ARLEN,
    output wire [2:0]                      M_AXIMM_96_ARSIZE,
    output wire [1:0]                      M_AXIMM_96_ARBURST,
    output wire [1:0]                      M_AXIMM_96_ARLOCK,
    output wire [3:0]                      M_AXIMM_96_ARCACHE,
    output wire [2:0]                      M_AXIMM_96_ARPROT,
    output wire [3:0]                      M_AXIMM_96_ARREGION,
    output wire [3:0]                      M_AXIMM_96_ARQOS,
    output wire                            M_AXIMM_96_ARVALID,
    input  wire                            M_AXIMM_96_ARREADY,
    input  wire [M_AXIMM_96_DATA_WIDTH-1:0]   M_AXIMM_96_RDATA,
    input  wire [1:0]                      M_AXIMM_96_RRESP,
    input  wire                            M_AXIMM_96_RLAST,
    input  wire                            M_AXIMM_96_RVALID,
    output wire                            M_AXIMM_96_RREADY,
    //AXI-MM pass-through interface 97
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_97_AWADDR,
    input wire [7:0]                      AP_AXIMM_97_AWLEN,
    input wire [2:0]                      AP_AXIMM_97_AWSIZE,
    input wire [1:0]                      AP_AXIMM_97_AWBURST,
    input wire [1:0]                      AP_AXIMM_97_AWLOCK,
    input wire [3:0]                      AP_AXIMM_97_AWCACHE,
    input wire [2:0]                      AP_AXIMM_97_AWPROT,
    input wire [3:0]                      AP_AXIMM_97_AWREGION,
    input wire [3:0]                      AP_AXIMM_97_AWQOS,
    input wire                            AP_AXIMM_97_AWVALID,
    output  wire                            AP_AXIMM_97_AWREADY,
    input wire [M_AXIMM_97_DATA_WIDTH-1:0]   AP_AXIMM_97_WDATA,
    input wire [M_AXIMM_97_DATA_WIDTH/8-1:0] AP_AXIMM_97_WSTRB,
    input wire                            AP_AXIMM_97_WLAST,
    input wire                            AP_AXIMM_97_WVALID,
    output  wire                            AP_AXIMM_97_WREADY,
    output  wire [1:0]                      AP_AXIMM_97_BRESP,
    output  wire                            AP_AXIMM_97_BVALID,
    input wire                            AP_AXIMM_97_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_97_ARADDR,
    input wire [7:0]                      AP_AXIMM_97_ARLEN,
    input wire [2:0]                      AP_AXIMM_97_ARSIZE,
    input wire [1:0]                      AP_AXIMM_97_ARBURST,
    input wire [1:0]                      AP_AXIMM_97_ARLOCK,
    input wire [3:0]                      AP_AXIMM_97_ARCACHE,
    input wire [2:0]                      AP_AXIMM_97_ARPROT,
    input wire [3:0]                      AP_AXIMM_97_ARREGION,
    input wire [3:0]                      AP_AXIMM_97_ARQOS,
    input wire                            AP_AXIMM_97_ARVALID,
    output  wire                            AP_AXIMM_97_ARREADY,
    output  wire [M_AXIMM_97_DATA_WIDTH-1:0]   AP_AXIMM_97_RDATA,
    output  wire [1:0]                      AP_AXIMM_97_RRESP,
    output  wire                            AP_AXIMM_97_RLAST,
    output  wire                            AP_AXIMM_97_RVALID,
    input  wire                            AP_AXIMM_97_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_97_AWADDR,
    output wire [7:0]                      M_AXIMM_97_AWLEN,
    output wire [2:0]                      M_AXIMM_97_AWSIZE,
    output wire [1:0]                      M_AXIMM_97_AWBURST,
    output wire [1:0]                      M_AXIMM_97_AWLOCK,
    output wire [3:0]                      M_AXIMM_97_AWCACHE,
    output wire [2:0]                      M_AXIMM_97_AWPROT,
    output wire [3:0]                      M_AXIMM_97_AWREGION,
    output wire [3:0]                      M_AXIMM_97_AWQOS,
    output wire                            M_AXIMM_97_AWVALID,
    input  wire                            M_AXIMM_97_AWREADY,
    output wire [M_AXIMM_97_DATA_WIDTH-1:0]   M_AXIMM_97_WDATA,
    output wire [M_AXIMM_97_DATA_WIDTH/8-1:0] M_AXIMM_97_WSTRB,
    output wire                            M_AXIMM_97_WLAST,
    output wire                            M_AXIMM_97_WVALID,
    input  wire                            M_AXIMM_97_WREADY,
    input  wire [1:0]                      M_AXIMM_97_BRESP,
    input  wire                            M_AXIMM_97_BVALID,
    output wire                            M_AXIMM_97_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_97_ARADDR,
    output wire [7:0]                      M_AXIMM_97_ARLEN,
    output wire [2:0]                      M_AXIMM_97_ARSIZE,
    output wire [1:0]                      M_AXIMM_97_ARBURST,
    output wire [1:0]                      M_AXIMM_97_ARLOCK,
    output wire [3:0]                      M_AXIMM_97_ARCACHE,
    output wire [2:0]                      M_AXIMM_97_ARPROT,
    output wire [3:0]                      M_AXIMM_97_ARREGION,
    output wire [3:0]                      M_AXIMM_97_ARQOS,
    output wire                            M_AXIMM_97_ARVALID,
    input  wire                            M_AXIMM_97_ARREADY,
    input  wire [M_AXIMM_97_DATA_WIDTH-1:0]   M_AXIMM_97_RDATA,
    input  wire [1:0]                      M_AXIMM_97_RRESP,
    input  wire                            M_AXIMM_97_RLAST,
    input  wire                            M_AXIMM_97_RVALID,
    output wire                            M_AXIMM_97_RREADY,
    //AXI-MM pass-through interface 98
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_98_AWADDR,
    input wire [7:0]                      AP_AXIMM_98_AWLEN,
    input wire [2:0]                      AP_AXIMM_98_AWSIZE,
    input wire [1:0]                      AP_AXIMM_98_AWBURST,
    input wire [1:0]                      AP_AXIMM_98_AWLOCK,
    input wire [3:0]                      AP_AXIMM_98_AWCACHE,
    input wire [2:0]                      AP_AXIMM_98_AWPROT,
    input wire [3:0]                      AP_AXIMM_98_AWREGION,
    input wire [3:0]                      AP_AXIMM_98_AWQOS,
    input wire                            AP_AXIMM_98_AWVALID,
    output  wire                            AP_AXIMM_98_AWREADY,
    input wire [M_AXIMM_98_DATA_WIDTH-1:0]   AP_AXIMM_98_WDATA,
    input wire [M_AXIMM_98_DATA_WIDTH/8-1:0] AP_AXIMM_98_WSTRB,
    input wire                            AP_AXIMM_98_WLAST,
    input wire                            AP_AXIMM_98_WVALID,
    output  wire                            AP_AXIMM_98_WREADY,
    output  wire [1:0]                      AP_AXIMM_98_BRESP,
    output  wire                            AP_AXIMM_98_BVALID,
    input wire                            AP_AXIMM_98_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_98_ARADDR,
    input wire [7:0]                      AP_AXIMM_98_ARLEN,
    input wire [2:0]                      AP_AXIMM_98_ARSIZE,
    input wire [1:0]                      AP_AXIMM_98_ARBURST,
    input wire [1:0]                      AP_AXIMM_98_ARLOCK,
    input wire [3:0]                      AP_AXIMM_98_ARCACHE,
    input wire [2:0]                      AP_AXIMM_98_ARPROT,
    input wire [3:0]                      AP_AXIMM_98_ARREGION,
    input wire [3:0]                      AP_AXIMM_98_ARQOS,
    input wire                            AP_AXIMM_98_ARVALID,
    output  wire                            AP_AXIMM_98_ARREADY,
    output  wire [M_AXIMM_98_DATA_WIDTH-1:0]   AP_AXIMM_98_RDATA,
    output  wire [1:0]                      AP_AXIMM_98_RRESP,
    output  wire                            AP_AXIMM_98_RLAST,
    output  wire                            AP_AXIMM_98_RVALID,
    input  wire                            AP_AXIMM_98_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_98_AWADDR,
    output wire [7:0]                      M_AXIMM_98_AWLEN,
    output wire [2:0]                      M_AXIMM_98_AWSIZE,
    output wire [1:0]                      M_AXIMM_98_AWBURST,
    output wire [1:0]                      M_AXIMM_98_AWLOCK,
    output wire [3:0]                      M_AXIMM_98_AWCACHE,
    output wire [2:0]                      M_AXIMM_98_AWPROT,
    output wire [3:0]                      M_AXIMM_98_AWREGION,
    output wire [3:0]                      M_AXIMM_98_AWQOS,
    output wire                            M_AXIMM_98_AWVALID,
    input  wire                            M_AXIMM_98_AWREADY,
    output wire [M_AXIMM_98_DATA_WIDTH-1:0]   M_AXIMM_98_WDATA,
    output wire [M_AXIMM_98_DATA_WIDTH/8-1:0] M_AXIMM_98_WSTRB,
    output wire                            M_AXIMM_98_WLAST,
    output wire                            M_AXIMM_98_WVALID,
    input  wire                            M_AXIMM_98_WREADY,
    input  wire [1:0]                      M_AXIMM_98_BRESP,
    input  wire                            M_AXIMM_98_BVALID,
    output wire                            M_AXIMM_98_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_98_ARADDR,
    output wire [7:0]                      M_AXIMM_98_ARLEN,
    output wire [2:0]                      M_AXIMM_98_ARSIZE,
    output wire [1:0]                      M_AXIMM_98_ARBURST,
    output wire [1:0]                      M_AXIMM_98_ARLOCK,
    output wire [3:0]                      M_AXIMM_98_ARCACHE,
    output wire [2:0]                      M_AXIMM_98_ARPROT,
    output wire [3:0]                      M_AXIMM_98_ARREGION,
    output wire [3:0]                      M_AXIMM_98_ARQOS,
    output wire                            M_AXIMM_98_ARVALID,
    input  wire                            M_AXIMM_98_ARREADY,
    input  wire [M_AXIMM_98_DATA_WIDTH-1:0]   M_AXIMM_98_RDATA,
    input  wire [1:0]                      M_AXIMM_98_RRESP,
    input  wire                            M_AXIMM_98_RLAST,
    input  wire                            M_AXIMM_98_RVALID,
    output wire                            M_AXIMM_98_RREADY,
    //AXI-MM pass-through interface 99
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_99_AWADDR,
    input wire [7:0]                      AP_AXIMM_99_AWLEN,
    input wire [2:0]                      AP_AXIMM_99_AWSIZE,
    input wire [1:0]                      AP_AXIMM_99_AWBURST,
    input wire [1:0]                      AP_AXIMM_99_AWLOCK,
    input wire [3:0]                      AP_AXIMM_99_AWCACHE,
    input wire [2:0]                      AP_AXIMM_99_AWPROT,
    input wire [3:0]                      AP_AXIMM_99_AWREGION,
    input wire [3:0]                      AP_AXIMM_99_AWQOS,
    input wire                            AP_AXIMM_99_AWVALID,
    output  wire                            AP_AXIMM_99_AWREADY,
    input wire [M_AXIMM_99_DATA_WIDTH-1:0]   AP_AXIMM_99_WDATA,
    input wire [M_AXIMM_99_DATA_WIDTH/8-1:0] AP_AXIMM_99_WSTRB,
    input wire                            AP_AXIMM_99_WLAST,
    input wire                            AP_AXIMM_99_WVALID,
    output  wire                            AP_AXIMM_99_WREADY,
    output  wire [1:0]                      AP_AXIMM_99_BRESP,
    output  wire                            AP_AXIMM_99_BVALID,
    input wire                            AP_AXIMM_99_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_99_ARADDR,
    input wire [7:0]                      AP_AXIMM_99_ARLEN,
    input wire [2:0]                      AP_AXIMM_99_ARSIZE,
    input wire [1:0]                      AP_AXIMM_99_ARBURST,
    input wire [1:0]                      AP_AXIMM_99_ARLOCK,
    input wire [3:0]                      AP_AXIMM_99_ARCACHE,
    input wire [2:0]                      AP_AXIMM_99_ARPROT,
    input wire [3:0]                      AP_AXIMM_99_ARREGION,
    input wire [3:0]                      AP_AXIMM_99_ARQOS,
    input wire                            AP_AXIMM_99_ARVALID,
    output  wire                            AP_AXIMM_99_ARREADY,
    output  wire [M_AXIMM_99_DATA_WIDTH-1:0]   AP_AXIMM_99_RDATA,
    output  wire [1:0]                      AP_AXIMM_99_RRESP,
    output  wire                            AP_AXIMM_99_RLAST,
    output  wire                            AP_AXIMM_99_RVALID,
    input  wire                            AP_AXIMM_99_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_99_AWADDR,
    output wire [7:0]                      M_AXIMM_99_AWLEN,
    output wire [2:0]                      M_AXIMM_99_AWSIZE,
    output wire [1:0]                      M_AXIMM_99_AWBURST,
    output wire [1:0]                      M_AXIMM_99_AWLOCK,
    output wire [3:0]                      M_AXIMM_99_AWCACHE,
    output wire [2:0]                      M_AXIMM_99_AWPROT,
    output wire [3:0]                      M_AXIMM_99_AWREGION,
    output wire [3:0]                      M_AXIMM_99_AWQOS,
    output wire                            M_AXIMM_99_AWVALID,
    input  wire                            M_AXIMM_99_AWREADY,
    output wire [M_AXIMM_99_DATA_WIDTH-1:0]   M_AXIMM_99_WDATA,
    output wire [M_AXIMM_99_DATA_WIDTH/8-1:0] M_AXIMM_99_WSTRB,
    output wire                            M_AXIMM_99_WLAST,
    output wire                            M_AXIMM_99_WVALID,
    input  wire                            M_AXIMM_99_WREADY,
    input  wire [1:0]                      M_AXIMM_99_BRESP,
    input  wire                            M_AXIMM_99_BVALID,
    output wire                            M_AXIMM_99_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_99_ARADDR,
    output wire [7:0]                      M_AXIMM_99_ARLEN,
    output wire [2:0]                      M_AXIMM_99_ARSIZE,
    output wire [1:0]                      M_AXIMM_99_ARBURST,
    output wire [1:0]                      M_AXIMM_99_ARLOCK,
    output wire [3:0]                      M_AXIMM_99_ARCACHE,
    output wire [2:0]                      M_AXIMM_99_ARPROT,
    output wire [3:0]                      M_AXIMM_99_ARREGION,
    output wire [3:0]                      M_AXIMM_99_ARQOS,
    output wire                            M_AXIMM_99_ARVALID,
    input  wire                            M_AXIMM_99_ARREADY,
    input  wire [M_AXIMM_99_DATA_WIDTH-1:0]   M_AXIMM_99_RDATA,
    input  wire [1:0]                      M_AXIMM_99_RRESP,
    input  wire                            M_AXIMM_99_RLAST,
    input  wire                            M_AXIMM_99_RVALID,
    output wire                            M_AXIMM_99_RREADY,
    //AXI-MM pass-through interface 100
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_100_AWADDR,
    input wire [7:0]                      AP_AXIMM_100_AWLEN,
    input wire [2:0]                      AP_AXIMM_100_AWSIZE,
    input wire [1:0]                      AP_AXIMM_100_AWBURST,
    input wire [1:0]                      AP_AXIMM_100_AWLOCK,
    input wire [3:0]                      AP_AXIMM_100_AWCACHE,
    input wire [2:0]                      AP_AXIMM_100_AWPROT,
    input wire [3:0]                      AP_AXIMM_100_AWREGION,
    input wire [3:0]                      AP_AXIMM_100_AWQOS,
    input wire                            AP_AXIMM_100_AWVALID,
    output  wire                            AP_AXIMM_100_AWREADY,
    input wire [M_AXIMM_100_DATA_WIDTH-1:0]   AP_AXIMM_100_WDATA,
    input wire [M_AXIMM_100_DATA_WIDTH/8-1:0] AP_AXIMM_100_WSTRB,
    input wire                            AP_AXIMM_100_WLAST,
    input wire                            AP_AXIMM_100_WVALID,
    output  wire                            AP_AXIMM_100_WREADY,
    output  wire [1:0]                      AP_AXIMM_100_BRESP,
    output  wire                            AP_AXIMM_100_BVALID,
    input wire                            AP_AXIMM_100_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_100_ARADDR,
    input wire [7:0]                      AP_AXIMM_100_ARLEN,
    input wire [2:0]                      AP_AXIMM_100_ARSIZE,
    input wire [1:0]                      AP_AXIMM_100_ARBURST,
    input wire [1:0]                      AP_AXIMM_100_ARLOCK,
    input wire [3:0]                      AP_AXIMM_100_ARCACHE,
    input wire [2:0]                      AP_AXIMM_100_ARPROT,
    input wire [3:0]                      AP_AXIMM_100_ARREGION,
    input wire [3:0]                      AP_AXIMM_100_ARQOS,
    input wire                            AP_AXIMM_100_ARVALID,
    output  wire                            AP_AXIMM_100_ARREADY,
    output  wire [M_AXIMM_100_DATA_WIDTH-1:0]   AP_AXIMM_100_RDATA,
    output  wire [1:0]                      AP_AXIMM_100_RRESP,
    output  wire                            AP_AXIMM_100_RLAST,
    output  wire                            AP_AXIMM_100_RVALID,
    input  wire                            AP_AXIMM_100_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_100_AWADDR,
    output wire [7:0]                      M_AXIMM_100_AWLEN,
    output wire [2:0]                      M_AXIMM_100_AWSIZE,
    output wire [1:0]                      M_AXIMM_100_AWBURST,
    output wire [1:0]                      M_AXIMM_100_AWLOCK,
    output wire [3:0]                      M_AXIMM_100_AWCACHE,
    output wire [2:0]                      M_AXIMM_100_AWPROT,
    output wire [3:0]                      M_AXIMM_100_AWREGION,
    output wire [3:0]                      M_AXIMM_100_AWQOS,
    output wire                            M_AXIMM_100_AWVALID,
    input  wire                            M_AXIMM_100_AWREADY,
    output wire [M_AXIMM_100_DATA_WIDTH-1:0]   M_AXIMM_100_WDATA,
    output wire [M_AXIMM_100_DATA_WIDTH/8-1:0] M_AXIMM_100_WSTRB,
    output wire                            M_AXIMM_100_WLAST,
    output wire                            M_AXIMM_100_WVALID,
    input  wire                            M_AXIMM_100_WREADY,
    input  wire [1:0]                      M_AXIMM_100_BRESP,
    input  wire                            M_AXIMM_100_BVALID,
    output wire                            M_AXIMM_100_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_100_ARADDR,
    output wire [7:0]                      M_AXIMM_100_ARLEN,
    output wire [2:0]                      M_AXIMM_100_ARSIZE,
    output wire [1:0]                      M_AXIMM_100_ARBURST,
    output wire [1:0]                      M_AXIMM_100_ARLOCK,
    output wire [3:0]                      M_AXIMM_100_ARCACHE,
    output wire [2:0]                      M_AXIMM_100_ARPROT,
    output wire [3:0]                      M_AXIMM_100_ARREGION,
    output wire [3:0]                      M_AXIMM_100_ARQOS,
    output wire                            M_AXIMM_100_ARVALID,
    input  wire                            M_AXIMM_100_ARREADY,
    input  wire [M_AXIMM_100_DATA_WIDTH-1:0]   M_AXIMM_100_RDATA,
    input  wire [1:0]                      M_AXIMM_100_RRESP,
    input  wire                            M_AXIMM_100_RLAST,
    input  wire                            M_AXIMM_100_RVALID,
    output wire                            M_AXIMM_100_RREADY,
    //AXI-MM pass-through interface 101
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_101_AWADDR,
    input wire [7:0]                      AP_AXIMM_101_AWLEN,
    input wire [2:0]                      AP_AXIMM_101_AWSIZE,
    input wire [1:0]                      AP_AXIMM_101_AWBURST,
    input wire [1:0]                      AP_AXIMM_101_AWLOCK,
    input wire [3:0]                      AP_AXIMM_101_AWCACHE,
    input wire [2:0]                      AP_AXIMM_101_AWPROT,
    input wire [3:0]                      AP_AXIMM_101_AWREGION,
    input wire [3:0]                      AP_AXIMM_101_AWQOS,
    input wire                            AP_AXIMM_101_AWVALID,
    output  wire                            AP_AXIMM_101_AWREADY,
    input wire [M_AXIMM_101_DATA_WIDTH-1:0]   AP_AXIMM_101_WDATA,
    input wire [M_AXIMM_101_DATA_WIDTH/8-1:0] AP_AXIMM_101_WSTRB,
    input wire                            AP_AXIMM_101_WLAST,
    input wire                            AP_AXIMM_101_WVALID,
    output  wire                            AP_AXIMM_101_WREADY,
    output  wire [1:0]                      AP_AXIMM_101_BRESP,
    output  wire                            AP_AXIMM_101_BVALID,
    input wire                            AP_AXIMM_101_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_101_ARADDR,
    input wire [7:0]                      AP_AXIMM_101_ARLEN,
    input wire [2:0]                      AP_AXIMM_101_ARSIZE,
    input wire [1:0]                      AP_AXIMM_101_ARBURST,
    input wire [1:0]                      AP_AXIMM_101_ARLOCK,
    input wire [3:0]                      AP_AXIMM_101_ARCACHE,
    input wire [2:0]                      AP_AXIMM_101_ARPROT,
    input wire [3:0]                      AP_AXIMM_101_ARREGION,
    input wire [3:0]                      AP_AXIMM_101_ARQOS,
    input wire                            AP_AXIMM_101_ARVALID,
    output  wire                            AP_AXIMM_101_ARREADY,
    output  wire [M_AXIMM_101_DATA_WIDTH-1:0]   AP_AXIMM_101_RDATA,
    output  wire [1:0]                      AP_AXIMM_101_RRESP,
    output  wire                            AP_AXIMM_101_RLAST,
    output  wire                            AP_AXIMM_101_RVALID,
    input  wire                            AP_AXIMM_101_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_101_AWADDR,
    output wire [7:0]                      M_AXIMM_101_AWLEN,
    output wire [2:0]                      M_AXIMM_101_AWSIZE,
    output wire [1:0]                      M_AXIMM_101_AWBURST,
    output wire [1:0]                      M_AXIMM_101_AWLOCK,
    output wire [3:0]                      M_AXIMM_101_AWCACHE,
    output wire [2:0]                      M_AXIMM_101_AWPROT,
    output wire [3:0]                      M_AXIMM_101_AWREGION,
    output wire [3:0]                      M_AXIMM_101_AWQOS,
    output wire                            M_AXIMM_101_AWVALID,
    input  wire                            M_AXIMM_101_AWREADY,
    output wire [M_AXIMM_101_DATA_WIDTH-1:0]   M_AXIMM_101_WDATA,
    output wire [M_AXIMM_101_DATA_WIDTH/8-1:0] M_AXIMM_101_WSTRB,
    output wire                            M_AXIMM_101_WLAST,
    output wire                            M_AXIMM_101_WVALID,
    input  wire                            M_AXIMM_101_WREADY,
    input  wire [1:0]                      M_AXIMM_101_BRESP,
    input  wire                            M_AXIMM_101_BVALID,
    output wire                            M_AXIMM_101_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_101_ARADDR,
    output wire [7:0]                      M_AXIMM_101_ARLEN,
    output wire [2:0]                      M_AXIMM_101_ARSIZE,
    output wire [1:0]                      M_AXIMM_101_ARBURST,
    output wire [1:0]                      M_AXIMM_101_ARLOCK,
    output wire [3:0]                      M_AXIMM_101_ARCACHE,
    output wire [2:0]                      M_AXIMM_101_ARPROT,
    output wire [3:0]                      M_AXIMM_101_ARREGION,
    output wire [3:0]                      M_AXIMM_101_ARQOS,
    output wire                            M_AXIMM_101_ARVALID,
    input  wire                            M_AXIMM_101_ARREADY,
    input  wire [M_AXIMM_101_DATA_WIDTH-1:0]   M_AXIMM_101_RDATA,
    input  wire [1:0]                      M_AXIMM_101_RRESP,
    input  wire                            M_AXIMM_101_RLAST,
    input  wire                            M_AXIMM_101_RVALID,
    output wire                            M_AXIMM_101_RREADY,
    //AXI-MM pass-through interface 102
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_102_AWADDR,
    input wire [7:0]                      AP_AXIMM_102_AWLEN,
    input wire [2:0]                      AP_AXIMM_102_AWSIZE,
    input wire [1:0]                      AP_AXIMM_102_AWBURST,
    input wire [1:0]                      AP_AXIMM_102_AWLOCK,
    input wire [3:0]                      AP_AXIMM_102_AWCACHE,
    input wire [2:0]                      AP_AXIMM_102_AWPROT,
    input wire [3:0]                      AP_AXIMM_102_AWREGION,
    input wire [3:0]                      AP_AXIMM_102_AWQOS,
    input wire                            AP_AXIMM_102_AWVALID,
    output  wire                            AP_AXIMM_102_AWREADY,
    input wire [M_AXIMM_102_DATA_WIDTH-1:0]   AP_AXIMM_102_WDATA,
    input wire [M_AXIMM_102_DATA_WIDTH/8-1:0] AP_AXIMM_102_WSTRB,
    input wire                            AP_AXIMM_102_WLAST,
    input wire                            AP_AXIMM_102_WVALID,
    output  wire                            AP_AXIMM_102_WREADY,
    output  wire [1:0]                      AP_AXIMM_102_BRESP,
    output  wire                            AP_AXIMM_102_BVALID,
    input wire                            AP_AXIMM_102_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_102_ARADDR,
    input wire [7:0]                      AP_AXIMM_102_ARLEN,
    input wire [2:0]                      AP_AXIMM_102_ARSIZE,
    input wire [1:0]                      AP_AXIMM_102_ARBURST,
    input wire [1:0]                      AP_AXIMM_102_ARLOCK,
    input wire [3:0]                      AP_AXIMM_102_ARCACHE,
    input wire [2:0]                      AP_AXIMM_102_ARPROT,
    input wire [3:0]                      AP_AXIMM_102_ARREGION,
    input wire [3:0]                      AP_AXIMM_102_ARQOS,
    input wire                            AP_AXIMM_102_ARVALID,
    output  wire                            AP_AXIMM_102_ARREADY,
    output  wire [M_AXIMM_102_DATA_WIDTH-1:0]   AP_AXIMM_102_RDATA,
    output  wire [1:0]                      AP_AXIMM_102_RRESP,
    output  wire                            AP_AXIMM_102_RLAST,
    output  wire                            AP_AXIMM_102_RVALID,
    input  wire                            AP_AXIMM_102_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_102_AWADDR,
    output wire [7:0]                      M_AXIMM_102_AWLEN,
    output wire [2:0]                      M_AXIMM_102_AWSIZE,
    output wire [1:0]                      M_AXIMM_102_AWBURST,
    output wire [1:0]                      M_AXIMM_102_AWLOCK,
    output wire [3:0]                      M_AXIMM_102_AWCACHE,
    output wire [2:0]                      M_AXIMM_102_AWPROT,
    output wire [3:0]                      M_AXIMM_102_AWREGION,
    output wire [3:0]                      M_AXIMM_102_AWQOS,
    output wire                            M_AXIMM_102_AWVALID,
    input  wire                            M_AXIMM_102_AWREADY,
    output wire [M_AXIMM_102_DATA_WIDTH-1:0]   M_AXIMM_102_WDATA,
    output wire [M_AXIMM_102_DATA_WIDTH/8-1:0] M_AXIMM_102_WSTRB,
    output wire                            M_AXIMM_102_WLAST,
    output wire                            M_AXIMM_102_WVALID,
    input  wire                            M_AXIMM_102_WREADY,
    input  wire [1:0]                      M_AXIMM_102_BRESP,
    input  wire                            M_AXIMM_102_BVALID,
    output wire                            M_AXIMM_102_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_102_ARADDR,
    output wire [7:0]                      M_AXIMM_102_ARLEN,
    output wire [2:0]                      M_AXIMM_102_ARSIZE,
    output wire [1:0]                      M_AXIMM_102_ARBURST,
    output wire [1:0]                      M_AXIMM_102_ARLOCK,
    output wire [3:0]                      M_AXIMM_102_ARCACHE,
    output wire [2:0]                      M_AXIMM_102_ARPROT,
    output wire [3:0]                      M_AXIMM_102_ARREGION,
    output wire [3:0]                      M_AXIMM_102_ARQOS,
    output wire                            M_AXIMM_102_ARVALID,
    input  wire                            M_AXIMM_102_ARREADY,
    input  wire [M_AXIMM_102_DATA_WIDTH-1:0]   M_AXIMM_102_RDATA,
    input  wire [1:0]                      M_AXIMM_102_RRESP,
    input  wire                            M_AXIMM_102_RLAST,
    input  wire                            M_AXIMM_102_RVALID,
    output wire                            M_AXIMM_102_RREADY,
    //AXI-MM pass-through interface 103
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_103_AWADDR,
    input wire [7:0]                      AP_AXIMM_103_AWLEN,
    input wire [2:0]                      AP_AXIMM_103_AWSIZE,
    input wire [1:0]                      AP_AXIMM_103_AWBURST,
    input wire [1:0]                      AP_AXIMM_103_AWLOCK,
    input wire [3:0]                      AP_AXIMM_103_AWCACHE,
    input wire [2:0]                      AP_AXIMM_103_AWPROT,
    input wire [3:0]                      AP_AXIMM_103_AWREGION,
    input wire [3:0]                      AP_AXIMM_103_AWQOS,
    input wire                            AP_AXIMM_103_AWVALID,
    output  wire                            AP_AXIMM_103_AWREADY,
    input wire [M_AXIMM_103_DATA_WIDTH-1:0]   AP_AXIMM_103_WDATA,
    input wire [M_AXIMM_103_DATA_WIDTH/8-1:0] AP_AXIMM_103_WSTRB,
    input wire                            AP_AXIMM_103_WLAST,
    input wire                            AP_AXIMM_103_WVALID,
    output  wire                            AP_AXIMM_103_WREADY,
    output  wire [1:0]                      AP_AXIMM_103_BRESP,
    output  wire                            AP_AXIMM_103_BVALID,
    input wire                            AP_AXIMM_103_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_103_ARADDR,
    input wire [7:0]                      AP_AXIMM_103_ARLEN,
    input wire [2:0]                      AP_AXIMM_103_ARSIZE,
    input wire [1:0]                      AP_AXIMM_103_ARBURST,
    input wire [1:0]                      AP_AXIMM_103_ARLOCK,
    input wire [3:0]                      AP_AXIMM_103_ARCACHE,
    input wire [2:0]                      AP_AXIMM_103_ARPROT,
    input wire [3:0]                      AP_AXIMM_103_ARREGION,
    input wire [3:0]                      AP_AXIMM_103_ARQOS,
    input wire                            AP_AXIMM_103_ARVALID,
    output  wire                            AP_AXIMM_103_ARREADY,
    output  wire [M_AXIMM_103_DATA_WIDTH-1:0]   AP_AXIMM_103_RDATA,
    output  wire [1:0]                      AP_AXIMM_103_RRESP,
    output  wire                            AP_AXIMM_103_RLAST,
    output  wire                            AP_AXIMM_103_RVALID,
    input  wire                            AP_AXIMM_103_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_103_AWADDR,
    output wire [7:0]                      M_AXIMM_103_AWLEN,
    output wire [2:0]                      M_AXIMM_103_AWSIZE,
    output wire [1:0]                      M_AXIMM_103_AWBURST,
    output wire [1:0]                      M_AXIMM_103_AWLOCK,
    output wire [3:0]                      M_AXIMM_103_AWCACHE,
    output wire [2:0]                      M_AXIMM_103_AWPROT,
    output wire [3:0]                      M_AXIMM_103_AWREGION,
    output wire [3:0]                      M_AXIMM_103_AWQOS,
    output wire                            M_AXIMM_103_AWVALID,
    input  wire                            M_AXIMM_103_AWREADY,
    output wire [M_AXIMM_103_DATA_WIDTH-1:0]   M_AXIMM_103_WDATA,
    output wire [M_AXIMM_103_DATA_WIDTH/8-1:0] M_AXIMM_103_WSTRB,
    output wire                            M_AXIMM_103_WLAST,
    output wire                            M_AXIMM_103_WVALID,
    input  wire                            M_AXIMM_103_WREADY,
    input  wire [1:0]                      M_AXIMM_103_BRESP,
    input  wire                            M_AXIMM_103_BVALID,
    output wire                            M_AXIMM_103_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_103_ARADDR,
    output wire [7:0]                      M_AXIMM_103_ARLEN,
    output wire [2:0]                      M_AXIMM_103_ARSIZE,
    output wire [1:0]                      M_AXIMM_103_ARBURST,
    output wire [1:0]                      M_AXIMM_103_ARLOCK,
    output wire [3:0]                      M_AXIMM_103_ARCACHE,
    output wire [2:0]                      M_AXIMM_103_ARPROT,
    output wire [3:0]                      M_AXIMM_103_ARREGION,
    output wire [3:0]                      M_AXIMM_103_ARQOS,
    output wire                            M_AXIMM_103_ARVALID,
    input  wire                            M_AXIMM_103_ARREADY,
    input  wire [M_AXIMM_103_DATA_WIDTH-1:0]   M_AXIMM_103_RDATA,
    input  wire [1:0]                      M_AXIMM_103_RRESP,
    input  wire                            M_AXIMM_103_RLAST,
    input  wire                            M_AXIMM_103_RVALID,
    output wire                            M_AXIMM_103_RREADY,
    //AXI-MM pass-through interface 104
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_104_AWADDR,
    input wire [7:0]                      AP_AXIMM_104_AWLEN,
    input wire [2:0]                      AP_AXIMM_104_AWSIZE,
    input wire [1:0]                      AP_AXIMM_104_AWBURST,
    input wire [1:0]                      AP_AXIMM_104_AWLOCK,
    input wire [3:0]                      AP_AXIMM_104_AWCACHE,
    input wire [2:0]                      AP_AXIMM_104_AWPROT,
    input wire [3:0]                      AP_AXIMM_104_AWREGION,
    input wire [3:0]                      AP_AXIMM_104_AWQOS,
    input wire                            AP_AXIMM_104_AWVALID,
    output  wire                            AP_AXIMM_104_AWREADY,
    input wire [M_AXIMM_104_DATA_WIDTH-1:0]   AP_AXIMM_104_WDATA,
    input wire [M_AXIMM_104_DATA_WIDTH/8-1:0] AP_AXIMM_104_WSTRB,
    input wire                            AP_AXIMM_104_WLAST,
    input wire                            AP_AXIMM_104_WVALID,
    output  wire                            AP_AXIMM_104_WREADY,
    output  wire [1:0]                      AP_AXIMM_104_BRESP,
    output  wire                            AP_AXIMM_104_BVALID,
    input wire                            AP_AXIMM_104_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_104_ARADDR,
    input wire [7:0]                      AP_AXIMM_104_ARLEN,
    input wire [2:0]                      AP_AXIMM_104_ARSIZE,
    input wire [1:0]                      AP_AXIMM_104_ARBURST,
    input wire [1:0]                      AP_AXIMM_104_ARLOCK,
    input wire [3:0]                      AP_AXIMM_104_ARCACHE,
    input wire [2:0]                      AP_AXIMM_104_ARPROT,
    input wire [3:0]                      AP_AXIMM_104_ARREGION,
    input wire [3:0]                      AP_AXIMM_104_ARQOS,
    input wire                            AP_AXIMM_104_ARVALID,
    output  wire                            AP_AXIMM_104_ARREADY,
    output  wire [M_AXIMM_104_DATA_WIDTH-1:0]   AP_AXIMM_104_RDATA,
    output  wire [1:0]                      AP_AXIMM_104_RRESP,
    output  wire                            AP_AXIMM_104_RLAST,
    output  wire                            AP_AXIMM_104_RVALID,
    input  wire                            AP_AXIMM_104_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_104_AWADDR,
    output wire [7:0]                      M_AXIMM_104_AWLEN,
    output wire [2:0]                      M_AXIMM_104_AWSIZE,
    output wire [1:0]                      M_AXIMM_104_AWBURST,
    output wire [1:0]                      M_AXIMM_104_AWLOCK,
    output wire [3:0]                      M_AXIMM_104_AWCACHE,
    output wire [2:0]                      M_AXIMM_104_AWPROT,
    output wire [3:0]                      M_AXIMM_104_AWREGION,
    output wire [3:0]                      M_AXIMM_104_AWQOS,
    output wire                            M_AXIMM_104_AWVALID,
    input  wire                            M_AXIMM_104_AWREADY,
    output wire [M_AXIMM_104_DATA_WIDTH-1:0]   M_AXIMM_104_WDATA,
    output wire [M_AXIMM_104_DATA_WIDTH/8-1:0] M_AXIMM_104_WSTRB,
    output wire                            M_AXIMM_104_WLAST,
    output wire                            M_AXIMM_104_WVALID,
    input  wire                            M_AXIMM_104_WREADY,
    input  wire [1:0]                      M_AXIMM_104_BRESP,
    input  wire                            M_AXIMM_104_BVALID,
    output wire                            M_AXIMM_104_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_104_ARADDR,
    output wire [7:0]                      M_AXIMM_104_ARLEN,
    output wire [2:0]                      M_AXIMM_104_ARSIZE,
    output wire [1:0]                      M_AXIMM_104_ARBURST,
    output wire [1:0]                      M_AXIMM_104_ARLOCK,
    output wire [3:0]                      M_AXIMM_104_ARCACHE,
    output wire [2:0]                      M_AXIMM_104_ARPROT,
    output wire [3:0]                      M_AXIMM_104_ARREGION,
    output wire [3:0]                      M_AXIMM_104_ARQOS,
    output wire                            M_AXIMM_104_ARVALID,
    input  wire                            M_AXIMM_104_ARREADY,
    input  wire [M_AXIMM_104_DATA_WIDTH-1:0]   M_AXIMM_104_RDATA,
    input  wire [1:0]                      M_AXIMM_104_RRESP,
    input  wire                            M_AXIMM_104_RLAST,
    input  wire                            M_AXIMM_104_RVALID,
    output wire                            M_AXIMM_104_RREADY,
    //AXI-MM pass-through interface 105
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_105_AWADDR,
    input wire [7:0]                      AP_AXIMM_105_AWLEN,
    input wire [2:0]                      AP_AXIMM_105_AWSIZE,
    input wire [1:0]                      AP_AXIMM_105_AWBURST,
    input wire [1:0]                      AP_AXIMM_105_AWLOCK,
    input wire [3:0]                      AP_AXIMM_105_AWCACHE,
    input wire [2:0]                      AP_AXIMM_105_AWPROT,
    input wire [3:0]                      AP_AXIMM_105_AWREGION,
    input wire [3:0]                      AP_AXIMM_105_AWQOS,
    input wire                            AP_AXIMM_105_AWVALID,
    output  wire                            AP_AXIMM_105_AWREADY,
    input wire [M_AXIMM_105_DATA_WIDTH-1:0]   AP_AXIMM_105_WDATA,
    input wire [M_AXIMM_105_DATA_WIDTH/8-1:0] AP_AXIMM_105_WSTRB,
    input wire                            AP_AXIMM_105_WLAST,
    input wire                            AP_AXIMM_105_WVALID,
    output  wire                            AP_AXIMM_105_WREADY,
    output  wire [1:0]                      AP_AXIMM_105_BRESP,
    output  wire                            AP_AXIMM_105_BVALID,
    input wire                            AP_AXIMM_105_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_105_ARADDR,
    input wire [7:0]                      AP_AXIMM_105_ARLEN,
    input wire [2:0]                      AP_AXIMM_105_ARSIZE,
    input wire [1:0]                      AP_AXIMM_105_ARBURST,
    input wire [1:0]                      AP_AXIMM_105_ARLOCK,
    input wire [3:0]                      AP_AXIMM_105_ARCACHE,
    input wire [2:0]                      AP_AXIMM_105_ARPROT,
    input wire [3:0]                      AP_AXIMM_105_ARREGION,
    input wire [3:0]                      AP_AXIMM_105_ARQOS,
    input wire                            AP_AXIMM_105_ARVALID,
    output  wire                            AP_AXIMM_105_ARREADY,
    output  wire [M_AXIMM_105_DATA_WIDTH-1:0]   AP_AXIMM_105_RDATA,
    output  wire [1:0]                      AP_AXIMM_105_RRESP,
    output  wire                            AP_AXIMM_105_RLAST,
    output  wire                            AP_AXIMM_105_RVALID,
    input  wire                            AP_AXIMM_105_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_105_AWADDR,
    output wire [7:0]                      M_AXIMM_105_AWLEN,
    output wire [2:0]                      M_AXIMM_105_AWSIZE,
    output wire [1:0]                      M_AXIMM_105_AWBURST,
    output wire [1:0]                      M_AXIMM_105_AWLOCK,
    output wire [3:0]                      M_AXIMM_105_AWCACHE,
    output wire [2:0]                      M_AXIMM_105_AWPROT,
    output wire [3:0]                      M_AXIMM_105_AWREGION,
    output wire [3:0]                      M_AXIMM_105_AWQOS,
    output wire                            M_AXIMM_105_AWVALID,
    input  wire                            M_AXIMM_105_AWREADY,
    output wire [M_AXIMM_105_DATA_WIDTH-1:0]   M_AXIMM_105_WDATA,
    output wire [M_AXIMM_105_DATA_WIDTH/8-1:0] M_AXIMM_105_WSTRB,
    output wire                            M_AXIMM_105_WLAST,
    output wire                            M_AXIMM_105_WVALID,
    input  wire                            M_AXIMM_105_WREADY,
    input  wire [1:0]                      M_AXIMM_105_BRESP,
    input  wire                            M_AXIMM_105_BVALID,
    output wire                            M_AXIMM_105_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_105_ARADDR,
    output wire [7:0]                      M_AXIMM_105_ARLEN,
    output wire [2:0]                      M_AXIMM_105_ARSIZE,
    output wire [1:0]                      M_AXIMM_105_ARBURST,
    output wire [1:0]                      M_AXIMM_105_ARLOCK,
    output wire [3:0]                      M_AXIMM_105_ARCACHE,
    output wire [2:0]                      M_AXIMM_105_ARPROT,
    output wire [3:0]                      M_AXIMM_105_ARREGION,
    output wire [3:0]                      M_AXIMM_105_ARQOS,
    output wire                            M_AXIMM_105_ARVALID,
    input  wire                            M_AXIMM_105_ARREADY,
    input  wire [M_AXIMM_105_DATA_WIDTH-1:0]   M_AXIMM_105_RDATA,
    input  wire [1:0]                      M_AXIMM_105_RRESP,
    input  wire                            M_AXIMM_105_RLAST,
    input  wire                            M_AXIMM_105_RVALID,
    output wire                            M_AXIMM_105_RREADY,
    //AXI-MM pass-through interface 106
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_106_AWADDR,
    input wire [7:0]                      AP_AXIMM_106_AWLEN,
    input wire [2:0]                      AP_AXIMM_106_AWSIZE,
    input wire [1:0]                      AP_AXIMM_106_AWBURST,
    input wire [1:0]                      AP_AXIMM_106_AWLOCK,
    input wire [3:0]                      AP_AXIMM_106_AWCACHE,
    input wire [2:0]                      AP_AXIMM_106_AWPROT,
    input wire [3:0]                      AP_AXIMM_106_AWREGION,
    input wire [3:0]                      AP_AXIMM_106_AWQOS,
    input wire                            AP_AXIMM_106_AWVALID,
    output  wire                            AP_AXIMM_106_AWREADY,
    input wire [M_AXIMM_106_DATA_WIDTH-1:0]   AP_AXIMM_106_WDATA,
    input wire [M_AXIMM_106_DATA_WIDTH/8-1:0] AP_AXIMM_106_WSTRB,
    input wire                            AP_AXIMM_106_WLAST,
    input wire                            AP_AXIMM_106_WVALID,
    output  wire                            AP_AXIMM_106_WREADY,
    output  wire [1:0]                      AP_AXIMM_106_BRESP,
    output  wire                            AP_AXIMM_106_BVALID,
    input wire                            AP_AXIMM_106_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_106_ARADDR,
    input wire [7:0]                      AP_AXIMM_106_ARLEN,
    input wire [2:0]                      AP_AXIMM_106_ARSIZE,
    input wire [1:0]                      AP_AXIMM_106_ARBURST,
    input wire [1:0]                      AP_AXIMM_106_ARLOCK,
    input wire [3:0]                      AP_AXIMM_106_ARCACHE,
    input wire [2:0]                      AP_AXIMM_106_ARPROT,
    input wire [3:0]                      AP_AXIMM_106_ARREGION,
    input wire [3:0]                      AP_AXIMM_106_ARQOS,
    input wire                            AP_AXIMM_106_ARVALID,
    output  wire                            AP_AXIMM_106_ARREADY,
    output  wire [M_AXIMM_106_DATA_WIDTH-1:0]   AP_AXIMM_106_RDATA,
    output  wire [1:0]                      AP_AXIMM_106_RRESP,
    output  wire                            AP_AXIMM_106_RLAST,
    output  wire                            AP_AXIMM_106_RVALID,
    input  wire                            AP_AXIMM_106_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_106_AWADDR,
    output wire [7:0]                      M_AXIMM_106_AWLEN,
    output wire [2:0]                      M_AXIMM_106_AWSIZE,
    output wire [1:0]                      M_AXIMM_106_AWBURST,
    output wire [1:0]                      M_AXIMM_106_AWLOCK,
    output wire [3:0]                      M_AXIMM_106_AWCACHE,
    output wire [2:0]                      M_AXIMM_106_AWPROT,
    output wire [3:0]                      M_AXIMM_106_AWREGION,
    output wire [3:0]                      M_AXIMM_106_AWQOS,
    output wire                            M_AXIMM_106_AWVALID,
    input  wire                            M_AXIMM_106_AWREADY,
    output wire [M_AXIMM_106_DATA_WIDTH-1:0]   M_AXIMM_106_WDATA,
    output wire [M_AXIMM_106_DATA_WIDTH/8-1:0] M_AXIMM_106_WSTRB,
    output wire                            M_AXIMM_106_WLAST,
    output wire                            M_AXIMM_106_WVALID,
    input  wire                            M_AXIMM_106_WREADY,
    input  wire [1:0]                      M_AXIMM_106_BRESP,
    input  wire                            M_AXIMM_106_BVALID,
    output wire                            M_AXIMM_106_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_106_ARADDR,
    output wire [7:0]                      M_AXIMM_106_ARLEN,
    output wire [2:0]                      M_AXIMM_106_ARSIZE,
    output wire [1:0]                      M_AXIMM_106_ARBURST,
    output wire [1:0]                      M_AXIMM_106_ARLOCK,
    output wire [3:0]                      M_AXIMM_106_ARCACHE,
    output wire [2:0]                      M_AXIMM_106_ARPROT,
    output wire [3:0]                      M_AXIMM_106_ARREGION,
    output wire [3:0]                      M_AXIMM_106_ARQOS,
    output wire                            M_AXIMM_106_ARVALID,
    input  wire                            M_AXIMM_106_ARREADY,
    input  wire [M_AXIMM_106_DATA_WIDTH-1:0]   M_AXIMM_106_RDATA,
    input  wire [1:0]                      M_AXIMM_106_RRESP,
    input  wire                            M_AXIMM_106_RLAST,
    input  wire                            M_AXIMM_106_RVALID,
    output wire                            M_AXIMM_106_RREADY,
    //AXI-MM pass-through interface 107
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_107_AWADDR,
    input wire [7:0]                      AP_AXIMM_107_AWLEN,
    input wire [2:0]                      AP_AXIMM_107_AWSIZE,
    input wire [1:0]                      AP_AXIMM_107_AWBURST,
    input wire [1:0]                      AP_AXIMM_107_AWLOCK,
    input wire [3:0]                      AP_AXIMM_107_AWCACHE,
    input wire [2:0]                      AP_AXIMM_107_AWPROT,
    input wire [3:0]                      AP_AXIMM_107_AWREGION,
    input wire [3:0]                      AP_AXIMM_107_AWQOS,
    input wire                            AP_AXIMM_107_AWVALID,
    output  wire                            AP_AXIMM_107_AWREADY,
    input wire [M_AXIMM_107_DATA_WIDTH-1:0]   AP_AXIMM_107_WDATA,
    input wire [M_AXIMM_107_DATA_WIDTH/8-1:0] AP_AXIMM_107_WSTRB,
    input wire                            AP_AXIMM_107_WLAST,
    input wire                            AP_AXIMM_107_WVALID,
    output  wire                            AP_AXIMM_107_WREADY,
    output  wire [1:0]                      AP_AXIMM_107_BRESP,
    output  wire                            AP_AXIMM_107_BVALID,
    input wire                            AP_AXIMM_107_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_107_ARADDR,
    input wire [7:0]                      AP_AXIMM_107_ARLEN,
    input wire [2:0]                      AP_AXIMM_107_ARSIZE,
    input wire [1:0]                      AP_AXIMM_107_ARBURST,
    input wire [1:0]                      AP_AXIMM_107_ARLOCK,
    input wire [3:0]                      AP_AXIMM_107_ARCACHE,
    input wire [2:0]                      AP_AXIMM_107_ARPROT,
    input wire [3:0]                      AP_AXIMM_107_ARREGION,
    input wire [3:0]                      AP_AXIMM_107_ARQOS,
    input wire                            AP_AXIMM_107_ARVALID,
    output  wire                            AP_AXIMM_107_ARREADY,
    output  wire [M_AXIMM_107_DATA_WIDTH-1:0]   AP_AXIMM_107_RDATA,
    output  wire [1:0]                      AP_AXIMM_107_RRESP,
    output  wire                            AP_AXIMM_107_RLAST,
    output  wire                            AP_AXIMM_107_RVALID,
    input  wire                            AP_AXIMM_107_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_107_AWADDR,
    output wire [7:0]                      M_AXIMM_107_AWLEN,
    output wire [2:0]                      M_AXIMM_107_AWSIZE,
    output wire [1:0]                      M_AXIMM_107_AWBURST,
    output wire [1:0]                      M_AXIMM_107_AWLOCK,
    output wire [3:0]                      M_AXIMM_107_AWCACHE,
    output wire [2:0]                      M_AXIMM_107_AWPROT,
    output wire [3:0]                      M_AXIMM_107_AWREGION,
    output wire [3:0]                      M_AXIMM_107_AWQOS,
    output wire                            M_AXIMM_107_AWVALID,
    input  wire                            M_AXIMM_107_AWREADY,
    output wire [M_AXIMM_107_DATA_WIDTH-1:0]   M_AXIMM_107_WDATA,
    output wire [M_AXIMM_107_DATA_WIDTH/8-1:0] M_AXIMM_107_WSTRB,
    output wire                            M_AXIMM_107_WLAST,
    output wire                            M_AXIMM_107_WVALID,
    input  wire                            M_AXIMM_107_WREADY,
    input  wire [1:0]                      M_AXIMM_107_BRESP,
    input  wire                            M_AXIMM_107_BVALID,
    output wire                            M_AXIMM_107_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_107_ARADDR,
    output wire [7:0]                      M_AXIMM_107_ARLEN,
    output wire [2:0]                      M_AXIMM_107_ARSIZE,
    output wire [1:0]                      M_AXIMM_107_ARBURST,
    output wire [1:0]                      M_AXIMM_107_ARLOCK,
    output wire [3:0]                      M_AXIMM_107_ARCACHE,
    output wire [2:0]                      M_AXIMM_107_ARPROT,
    output wire [3:0]                      M_AXIMM_107_ARREGION,
    output wire [3:0]                      M_AXIMM_107_ARQOS,
    output wire                            M_AXIMM_107_ARVALID,
    input  wire                            M_AXIMM_107_ARREADY,
    input  wire [M_AXIMM_107_DATA_WIDTH-1:0]   M_AXIMM_107_RDATA,
    input  wire [1:0]                      M_AXIMM_107_RRESP,
    input  wire                            M_AXIMM_107_RLAST,
    input  wire                            M_AXIMM_107_RVALID,
    output wire                            M_AXIMM_107_RREADY,
    //AXI-MM pass-through interface 108
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_108_AWADDR,
    input wire [7:0]                      AP_AXIMM_108_AWLEN,
    input wire [2:0]                      AP_AXIMM_108_AWSIZE,
    input wire [1:0]                      AP_AXIMM_108_AWBURST,
    input wire [1:0]                      AP_AXIMM_108_AWLOCK,
    input wire [3:0]                      AP_AXIMM_108_AWCACHE,
    input wire [2:0]                      AP_AXIMM_108_AWPROT,
    input wire [3:0]                      AP_AXIMM_108_AWREGION,
    input wire [3:0]                      AP_AXIMM_108_AWQOS,
    input wire                            AP_AXIMM_108_AWVALID,
    output  wire                            AP_AXIMM_108_AWREADY,
    input wire [M_AXIMM_108_DATA_WIDTH-1:0]   AP_AXIMM_108_WDATA,
    input wire [M_AXIMM_108_DATA_WIDTH/8-1:0] AP_AXIMM_108_WSTRB,
    input wire                            AP_AXIMM_108_WLAST,
    input wire                            AP_AXIMM_108_WVALID,
    output  wire                            AP_AXIMM_108_WREADY,
    output  wire [1:0]                      AP_AXIMM_108_BRESP,
    output  wire                            AP_AXIMM_108_BVALID,
    input wire                            AP_AXIMM_108_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_108_ARADDR,
    input wire [7:0]                      AP_AXIMM_108_ARLEN,
    input wire [2:0]                      AP_AXIMM_108_ARSIZE,
    input wire [1:0]                      AP_AXIMM_108_ARBURST,
    input wire [1:0]                      AP_AXIMM_108_ARLOCK,
    input wire [3:0]                      AP_AXIMM_108_ARCACHE,
    input wire [2:0]                      AP_AXIMM_108_ARPROT,
    input wire [3:0]                      AP_AXIMM_108_ARREGION,
    input wire [3:0]                      AP_AXIMM_108_ARQOS,
    input wire                            AP_AXIMM_108_ARVALID,
    output  wire                            AP_AXIMM_108_ARREADY,
    output  wire [M_AXIMM_108_DATA_WIDTH-1:0]   AP_AXIMM_108_RDATA,
    output  wire [1:0]                      AP_AXIMM_108_RRESP,
    output  wire                            AP_AXIMM_108_RLAST,
    output  wire                            AP_AXIMM_108_RVALID,
    input  wire                            AP_AXIMM_108_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_108_AWADDR,
    output wire [7:0]                      M_AXIMM_108_AWLEN,
    output wire [2:0]                      M_AXIMM_108_AWSIZE,
    output wire [1:0]                      M_AXIMM_108_AWBURST,
    output wire [1:0]                      M_AXIMM_108_AWLOCK,
    output wire [3:0]                      M_AXIMM_108_AWCACHE,
    output wire [2:0]                      M_AXIMM_108_AWPROT,
    output wire [3:0]                      M_AXIMM_108_AWREGION,
    output wire [3:0]                      M_AXIMM_108_AWQOS,
    output wire                            M_AXIMM_108_AWVALID,
    input  wire                            M_AXIMM_108_AWREADY,
    output wire [M_AXIMM_108_DATA_WIDTH-1:0]   M_AXIMM_108_WDATA,
    output wire [M_AXIMM_108_DATA_WIDTH/8-1:0] M_AXIMM_108_WSTRB,
    output wire                            M_AXIMM_108_WLAST,
    output wire                            M_AXIMM_108_WVALID,
    input  wire                            M_AXIMM_108_WREADY,
    input  wire [1:0]                      M_AXIMM_108_BRESP,
    input  wire                            M_AXIMM_108_BVALID,
    output wire                            M_AXIMM_108_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_108_ARADDR,
    output wire [7:0]                      M_AXIMM_108_ARLEN,
    output wire [2:0]                      M_AXIMM_108_ARSIZE,
    output wire [1:0]                      M_AXIMM_108_ARBURST,
    output wire [1:0]                      M_AXIMM_108_ARLOCK,
    output wire [3:0]                      M_AXIMM_108_ARCACHE,
    output wire [2:0]                      M_AXIMM_108_ARPROT,
    output wire [3:0]                      M_AXIMM_108_ARREGION,
    output wire [3:0]                      M_AXIMM_108_ARQOS,
    output wire                            M_AXIMM_108_ARVALID,
    input  wire                            M_AXIMM_108_ARREADY,
    input  wire [M_AXIMM_108_DATA_WIDTH-1:0]   M_AXIMM_108_RDATA,
    input  wire [1:0]                      M_AXIMM_108_RRESP,
    input  wire                            M_AXIMM_108_RLAST,
    input  wire                            M_AXIMM_108_RVALID,
    output wire                            M_AXIMM_108_RREADY,
    //AXI-MM pass-through interface 109
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_109_AWADDR,
    input wire [7:0]                      AP_AXIMM_109_AWLEN,
    input wire [2:0]                      AP_AXIMM_109_AWSIZE,
    input wire [1:0]                      AP_AXIMM_109_AWBURST,
    input wire [1:0]                      AP_AXIMM_109_AWLOCK,
    input wire [3:0]                      AP_AXIMM_109_AWCACHE,
    input wire [2:0]                      AP_AXIMM_109_AWPROT,
    input wire [3:0]                      AP_AXIMM_109_AWREGION,
    input wire [3:0]                      AP_AXIMM_109_AWQOS,
    input wire                            AP_AXIMM_109_AWVALID,
    output  wire                            AP_AXIMM_109_AWREADY,
    input wire [M_AXIMM_109_DATA_WIDTH-1:0]   AP_AXIMM_109_WDATA,
    input wire [M_AXIMM_109_DATA_WIDTH/8-1:0] AP_AXIMM_109_WSTRB,
    input wire                            AP_AXIMM_109_WLAST,
    input wire                            AP_AXIMM_109_WVALID,
    output  wire                            AP_AXIMM_109_WREADY,
    output  wire [1:0]                      AP_AXIMM_109_BRESP,
    output  wire                            AP_AXIMM_109_BVALID,
    input wire                            AP_AXIMM_109_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_109_ARADDR,
    input wire [7:0]                      AP_AXIMM_109_ARLEN,
    input wire [2:0]                      AP_AXIMM_109_ARSIZE,
    input wire [1:0]                      AP_AXIMM_109_ARBURST,
    input wire [1:0]                      AP_AXIMM_109_ARLOCK,
    input wire [3:0]                      AP_AXIMM_109_ARCACHE,
    input wire [2:0]                      AP_AXIMM_109_ARPROT,
    input wire [3:0]                      AP_AXIMM_109_ARREGION,
    input wire [3:0]                      AP_AXIMM_109_ARQOS,
    input wire                            AP_AXIMM_109_ARVALID,
    output  wire                            AP_AXIMM_109_ARREADY,
    output  wire [M_AXIMM_109_DATA_WIDTH-1:0]   AP_AXIMM_109_RDATA,
    output  wire [1:0]                      AP_AXIMM_109_RRESP,
    output  wire                            AP_AXIMM_109_RLAST,
    output  wire                            AP_AXIMM_109_RVALID,
    input  wire                            AP_AXIMM_109_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_109_AWADDR,
    output wire [7:0]                      M_AXIMM_109_AWLEN,
    output wire [2:0]                      M_AXIMM_109_AWSIZE,
    output wire [1:0]                      M_AXIMM_109_AWBURST,
    output wire [1:0]                      M_AXIMM_109_AWLOCK,
    output wire [3:0]                      M_AXIMM_109_AWCACHE,
    output wire [2:0]                      M_AXIMM_109_AWPROT,
    output wire [3:0]                      M_AXIMM_109_AWREGION,
    output wire [3:0]                      M_AXIMM_109_AWQOS,
    output wire                            M_AXIMM_109_AWVALID,
    input  wire                            M_AXIMM_109_AWREADY,
    output wire [M_AXIMM_109_DATA_WIDTH-1:0]   M_AXIMM_109_WDATA,
    output wire [M_AXIMM_109_DATA_WIDTH/8-1:0] M_AXIMM_109_WSTRB,
    output wire                            M_AXIMM_109_WLAST,
    output wire                            M_AXIMM_109_WVALID,
    input  wire                            M_AXIMM_109_WREADY,
    input  wire [1:0]                      M_AXIMM_109_BRESP,
    input  wire                            M_AXIMM_109_BVALID,
    output wire                            M_AXIMM_109_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_109_ARADDR,
    output wire [7:0]                      M_AXIMM_109_ARLEN,
    output wire [2:0]                      M_AXIMM_109_ARSIZE,
    output wire [1:0]                      M_AXIMM_109_ARBURST,
    output wire [1:0]                      M_AXIMM_109_ARLOCK,
    output wire [3:0]                      M_AXIMM_109_ARCACHE,
    output wire [2:0]                      M_AXIMM_109_ARPROT,
    output wire [3:0]                      M_AXIMM_109_ARREGION,
    output wire [3:0]                      M_AXIMM_109_ARQOS,
    output wire                            M_AXIMM_109_ARVALID,
    input  wire                            M_AXIMM_109_ARREADY,
    input  wire [M_AXIMM_109_DATA_WIDTH-1:0]   M_AXIMM_109_RDATA,
    input  wire [1:0]                      M_AXIMM_109_RRESP,
    input  wire                            M_AXIMM_109_RLAST,
    input  wire                            M_AXIMM_109_RVALID,
    output wire                            M_AXIMM_109_RREADY,
    //AXI-MM pass-through interface 110
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_110_AWADDR,
    input wire [7:0]                      AP_AXIMM_110_AWLEN,
    input wire [2:0]                      AP_AXIMM_110_AWSIZE,
    input wire [1:0]                      AP_AXIMM_110_AWBURST,
    input wire [1:0]                      AP_AXIMM_110_AWLOCK,
    input wire [3:0]                      AP_AXIMM_110_AWCACHE,
    input wire [2:0]                      AP_AXIMM_110_AWPROT,
    input wire [3:0]                      AP_AXIMM_110_AWREGION,
    input wire [3:0]                      AP_AXIMM_110_AWQOS,
    input wire                            AP_AXIMM_110_AWVALID,
    output  wire                            AP_AXIMM_110_AWREADY,
    input wire [M_AXIMM_110_DATA_WIDTH-1:0]   AP_AXIMM_110_WDATA,
    input wire [M_AXIMM_110_DATA_WIDTH/8-1:0] AP_AXIMM_110_WSTRB,
    input wire                            AP_AXIMM_110_WLAST,
    input wire                            AP_AXIMM_110_WVALID,
    output  wire                            AP_AXIMM_110_WREADY,
    output  wire [1:0]                      AP_AXIMM_110_BRESP,
    output  wire                            AP_AXIMM_110_BVALID,
    input wire                            AP_AXIMM_110_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_110_ARADDR,
    input wire [7:0]                      AP_AXIMM_110_ARLEN,
    input wire [2:0]                      AP_AXIMM_110_ARSIZE,
    input wire [1:0]                      AP_AXIMM_110_ARBURST,
    input wire [1:0]                      AP_AXIMM_110_ARLOCK,
    input wire [3:0]                      AP_AXIMM_110_ARCACHE,
    input wire [2:0]                      AP_AXIMM_110_ARPROT,
    input wire [3:0]                      AP_AXIMM_110_ARREGION,
    input wire [3:0]                      AP_AXIMM_110_ARQOS,
    input wire                            AP_AXIMM_110_ARVALID,
    output  wire                            AP_AXIMM_110_ARREADY,
    output  wire [M_AXIMM_110_DATA_WIDTH-1:0]   AP_AXIMM_110_RDATA,
    output  wire [1:0]                      AP_AXIMM_110_RRESP,
    output  wire                            AP_AXIMM_110_RLAST,
    output  wire                            AP_AXIMM_110_RVALID,
    input  wire                            AP_AXIMM_110_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_110_AWADDR,
    output wire [7:0]                      M_AXIMM_110_AWLEN,
    output wire [2:0]                      M_AXIMM_110_AWSIZE,
    output wire [1:0]                      M_AXIMM_110_AWBURST,
    output wire [1:0]                      M_AXIMM_110_AWLOCK,
    output wire [3:0]                      M_AXIMM_110_AWCACHE,
    output wire [2:0]                      M_AXIMM_110_AWPROT,
    output wire [3:0]                      M_AXIMM_110_AWREGION,
    output wire [3:0]                      M_AXIMM_110_AWQOS,
    output wire                            M_AXIMM_110_AWVALID,
    input  wire                            M_AXIMM_110_AWREADY,
    output wire [M_AXIMM_110_DATA_WIDTH-1:0]   M_AXIMM_110_WDATA,
    output wire [M_AXIMM_110_DATA_WIDTH/8-1:0] M_AXIMM_110_WSTRB,
    output wire                            M_AXIMM_110_WLAST,
    output wire                            M_AXIMM_110_WVALID,
    input  wire                            M_AXIMM_110_WREADY,
    input  wire [1:0]                      M_AXIMM_110_BRESP,
    input  wire                            M_AXIMM_110_BVALID,
    output wire                            M_AXIMM_110_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_110_ARADDR,
    output wire [7:0]                      M_AXIMM_110_ARLEN,
    output wire [2:0]                      M_AXIMM_110_ARSIZE,
    output wire [1:0]                      M_AXIMM_110_ARBURST,
    output wire [1:0]                      M_AXIMM_110_ARLOCK,
    output wire [3:0]                      M_AXIMM_110_ARCACHE,
    output wire [2:0]                      M_AXIMM_110_ARPROT,
    output wire [3:0]                      M_AXIMM_110_ARREGION,
    output wire [3:0]                      M_AXIMM_110_ARQOS,
    output wire                            M_AXIMM_110_ARVALID,
    input  wire                            M_AXIMM_110_ARREADY,
    input  wire [M_AXIMM_110_DATA_WIDTH-1:0]   M_AXIMM_110_RDATA,
    input  wire [1:0]                      M_AXIMM_110_RRESP,
    input  wire                            M_AXIMM_110_RLAST,
    input  wire                            M_AXIMM_110_RVALID,
    output wire                            M_AXIMM_110_RREADY,
    //AXI-MM pass-through interface 111
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_111_AWADDR,
    input wire [7:0]                      AP_AXIMM_111_AWLEN,
    input wire [2:0]                      AP_AXIMM_111_AWSIZE,
    input wire [1:0]                      AP_AXIMM_111_AWBURST,
    input wire [1:0]                      AP_AXIMM_111_AWLOCK,
    input wire [3:0]                      AP_AXIMM_111_AWCACHE,
    input wire [2:0]                      AP_AXIMM_111_AWPROT,
    input wire [3:0]                      AP_AXIMM_111_AWREGION,
    input wire [3:0]                      AP_AXIMM_111_AWQOS,
    input wire                            AP_AXIMM_111_AWVALID,
    output  wire                            AP_AXIMM_111_AWREADY,
    input wire [M_AXIMM_111_DATA_WIDTH-1:0]   AP_AXIMM_111_WDATA,
    input wire [M_AXIMM_111_DATA_WIDTH/8-1:0] AP_AXIMM_111_WSTRB,
    input wire                            AP_AXIMM_111_WLAST,
    input wire                            AP_AXIMM_111_WVALID,
    output  wire                            AP_AXIMM_111_WREADY,
    output  wire [1:0]                      AP_AXIMM_111_BRESP,
    output  wire                            AP_AXIMM_111_BVALID,
    input wire                            AP_AXIMM_111_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_111_ARADDR,
    input wire [7:0]                      AP_AXIMM_111_ARLEN,
    input wire [2:0]                      AP_AXIMM_111_ARSIZE,
    input wire [1:0]                      AP_AXIMM_111_ARBURST,
    input wire [1:0]                      AP_AXIMM_111_ARLOCK,
    input wire [3:0]                      AP_AXIMM_111_ARCACHE,
    input wire [2:0]                      AP_AXIMM_111_ARPROT,
    input wire [3:0]                      AP_AXIMM_111_ARREGION,
    input wire [3:0]                      AP_AXIMM_111_ARQOS,
    input wire                            AP_AXIMM_111_ARVALID,
    output  wire                            AP_AXIMM_111_ARREADY,
    output  wire [M_AXIMM_111_DATA_WIDTH-1:0]   AP_AXIMM_111_RDATA,
    output  wire [1:0]                      AP_AXIMM_111_RRESP,
    output  wire                            AP_AXIMM_111_RLAST,
    output  wire                            AP_AXIMM_111_RVALID,
    input  wire                            AP_AXIMM_111_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_111_AWADDR,
    output wire [7:0]                      M_AXIMM_111_AWLEN,
    output wire [2:0]                      M_AXIMM_111_AWSIZE,
    output wire [1:0]                      M_AXIMM_111_AWBURST,
    output wire [1:0]                      M_AXIMM_111_AWLOCK,
    output wire [3:0]                      M_AXIMM_111_AWCACHE,
    output wire [2:0]                      M_AXIMM_111_AWPROT,
    output wire [3:0]                      M_AXIMM_111_AWREGION,
    output wire [3:0]                      M_AXIMM_111_AWQOS,
    output wire                            M_AXIMM_111_AWVALID,
    input  wire                            M_AXIMM_111_AWREADY,
    output wire [M_AXIMM_111_DATA_WIDTH-1:0]   M_AXIMM_111_WDATA,
    output wire [M_AXIMM_111_DATA_WIDTH/8-1:0] M_AXIMM_111_WSTRB,
    output wire                            M_AXIMM_111_WLAST,
    output wire                            M_AXIMM_111_WVALID,
    input  wire                            M_AXIMM_111_WREADY,
    input  wire [1:0]                      M_AXIMM_111_BRESP,
    input  wire                            M_AXIMM_111_BVALID,
    output wire                            M_AXIMM_111_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_111_ARADDR,
    output wire [7:0]                      M_AXIMM_111_ARLEN,
    output wire [2:0]                      M_AXIMM_111_ARSIZE,
    output wire [1:0]                      M_AXIMM_111_ARBURST,
    output wire [1:0]                      M_AXIMM_111_ARLOCK,
    output wire [3:0]                      M_AXIMM_111_ARCACHE,
    output wire [2:0]                      M_AXIMM_111_ARPROT,
    output wire [3:0]                      M_AXIMM_111_ARREGION,
    output wire [3:0]                      M_AXIMM_111_ARQOS,
    output wire                            M_AXIMM_111_ARVALID,
    input  wire                            M_AXIMM_111_ARREADY,
    input  wire [M_AXIMM_111_DATA_WIDTH-1:0]   M_AXIMM_111_RDATA,
    input  wire [1:0]                      M_AXIMM_111_RRESP,
    input  wire                            M_AXIMM_111_RLAST,
    input  wire                            M_AXIMM_111_RVALID,
    output wire                            M_AXIMM_111_RREADY,
    //AXI-MM pass-through interface 112
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_112_AWADDR,
    input wire [7:0]                      AP_AXIMM_112_AWLEN,
    input wire [2:0]                      AP_AXIMM_112_AWSIZE,
    input wire [1:0]                      AP_AXIMM_112_AWBURST,
    input wire [1:0]                      AP_AXIMM_112_AWLOCK,
    input wire [3:0]                      AP_AXIMM_112_AWCACHE,
    input wire [2:0]                      AP_AXIMM_112_AWPROT,
    input wire [3:0]                      AP_AXIMM_112_AWREGION,
    input wire [3:0]                      AP_AXIMM_112_AWQOS,
    input wire                            AP_AXIMM_112_AWVALID,
    output  wire                            AP_AXIMM_112_AWREADY,
    input wire [M_AXIMM_112_DATA_WIDTH-1:0]   AP_AXIMM_112_WDATA,
    input wire [M_AXIMM_112_DATA_WIDTH/8-1:0] AP_AXIMM_112_WSTRB,
    input wire                            AP_AXIMM_112_WLAST,
    input wire                            AP_AXIMM_112_WVALID,
    output  wire                            AP_AXIMM_112_WREADY,
    output  wire [1:0]                      AP_AXIMM_112_BRESP,
    output  wire                            AP_AXIMM_112_BVALID,
    input wire                            AP_AXIMM_112_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_112_ARADDR,
    input wire [7:0]                      AP_AXIMM_112_ARLEN,
    input wire [2:0]                      AP_AXIMM_112_ARSIZE,
    input wire [1:0]                      AP_AXIMM_112_ARBURST,
    input wire [1:0]                      AP_AXIMM_112_ARLOCK,
    input wire [3:0]                      AP_AXIMM_112_ARCACHE,
    input wire [2:0]                      AP_AXIMM_112_ARPROT,
    input wire [3:0]                      AP_AXIMM_112_ARREGION,
    input wire [3:0]                      AP_AXIMM_112_ARQOS,
    input wire                            AP_AXIMM_112_ARVALID,
    output  wire                            AP_AXIMM_112_ARREADY,
    output  wire [M_AXIMM_112_DATA_WIDTH-1:0]   AP_AXIMM_112_RDATA,
    output  wire [1:0]                      AP_AXIMM_112_RRESP,
    output  wire                            AP_AXIMM_112_RLAST,
    output  wire                            AP_AXIMM_112_RVALID,
    input  wire                            AP_AXIMM_112_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_112_AWADDR,
    output wire [7:0]                      M_AXIMM_112_AWLEN,
    output wire [2:0]                      M_AXIMM_112_AWSIZE,
    output wire [1:0]                      M_AXIMM_112_AWBURST,
    output wire [1:0]                      M_AXIMM_112_AWLOCK,
    output wire [3:0]                      M_AXIMM_112_AWCACHE,
    output wire [2:0]                      M_AXIMM_112_AWPROT,
    output wire [3:0]                      M_AXIMM_112_AWREGION,
    output wire [3:0]                      M_AXIMM_112_AWQOS,
    output wire                            M_AXIMM_112_AWVALID,
    input  wire                            M_AXIMM_112_AWREADY,
    output wire [M_AXIMM_112_DATA_WIDTH-1:0]   M_AXIMM_112_WDATA,
    output wire [M_AXIMM_112_DATA_WIDTH/8-1:0] M_AXIMM_112_WSTRB,
    output wire                            M_AXIMM_112_WLAST,
    output wire                            M_AXIMM_112_WVALID,
    input  wire                            M_AXIMM_112_WREADY,
    input  wire [1:0]                      M_AXIMM_112_BRESP,
    input  wire                            M_AXIMM_112_BVALID,
    output wire                            M_AXIMM_112_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_112_ARADDR,
    output wire [7:0]                      M_AXIMM_112_ARLEN,
    output wire [2:0]                      M_AXIMM_112_ARSIZE,
    output wire [1:0]                      M_AXIMM_112_ARBURST,
    output wire [1:0]                      M_AXIMM_112_ARLOCK,
    output wire [3:0]                      M_AXIMM_112_ARCACHE,
    output wire [2:0]                      M_AXIMM_112_ARPROT,
    output wire [3:0]                      M_AXIMM_112_ARREGION,
    output wire [3:0]                      M_AXIMM_112_ARQOS,
    output wire                            M_AXIMM_112_ARVALID,
    input  wire                            M_AXIMM_112_ARREADY,
    input  wire [M_AXIMM_112_DATA_WIDTH-1:0]   M_AXIMM_112_RDATA,
    input  wire [1:0]                      M_AXIMM_112_RRESP,
    input  wire                            M_AXIMM_112_RLAST,
    input  wire                            M_AXIMM_112_RVALID,
    output wire                            M_AXIMM_112_RREADY,
    //AXI-MM pass-through interface 113
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_113_AWADDR,
    input wire [7:0]                      AP_AXIMM_113_AWLEN,
    input wire [2:0]                      AP_AXIMM_113_AWSIZE,
    input wire [1:0]                      AP_AXIMM_113_AWBURST,
    input wire [1:0]                      AP_AXIMM_113_AWLOCK,
    input wire [3:0]                      AP_AXIMM_113_AWCACHE,
    input wire [2:0]                      AP_AXIMM_113_AWPROT,
    input wire [3:0]                      AP_AXIMM_113_AWREGION,
    input wire [3:0]                      AP_AXIMM_113_AWQOS,
    input wire                            AP_AXIMM_113_AWVALID,
    output  wire                            AP_AXIMM_113_AWREADY,
    input wire [M_AXIMM_113_DATA_WIDTH-1:0]   AP_AXIMM_113_WDATA,
    input wire [M_AXIMM_113_DATA_WIDTH/8-1:0] AP_AXIMM_113_WSTRB,
    input wire                            AP_AXIMM_113_WLAST,
    input wire                            AP_AXIMM_113_WVALID,
    output  wire                            AP_AXIMM_113_WREADY,
    output  wire [1:0]                      AP_AXIMM_113_BRESP,
    output  wire                            AP_AXIMM_113_BVALID,
    input wire                            AP_AXIMM_113_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_113_ARADDR,
    input wire [7:0]                      AP_AXIMM_113_ARLEN,
    input wire [2:0]                      AP_AXIMM_113_ARSIZE,
    input wire [1:0]                      AP_AXIMM_113_ARBURST,
    input wire [1:0]                      AP_AXIMM_113_ARLOCK,
    input wire [3:0]                      AP_AXIMM_113_ARCACHE,
    input wire [2:0]                      AP_AXIMM_113_ARPROT,
    input wire [3:0]                      AP_AXIMM_113_ARREGION,
    input wire [3:0]                      AP_AXIMM_113_ARQOS,
    input wire                            AP_AXIMM_113_ARVALID,
    output  wire                            AP_AXIMM_113_ARREADY,
    output  wire [M_AXIMM_113_DATA_WIDTH-1:0]   AP_AXIMM_113_RDATA,
    output  wire [1:0]                      AP_AXIMM_113_RRESP,
    output  wire                            AP_AXIMM_113_RLAST,
    output  wire                            AP_AXIMM_113_RVALID,
    input  wire                            AP_AXIMM_113_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_113_AWADDR,
    output wire [7:0]                      M_AXIMM_113_AWLEN,
    output wire [2:0]                      M_AXIMM_113_AWSIZE,
    output wire [1:0]                      M_AXIMM_113_AWBURST,
    output wire [1:0]                      M_AXIMM_113_AWLOCK,
    output wire [3:0]                      M_AXIMM_113_AWCACHE,
    output wire [2:0]                      M_AXIMM_113_AWPROT,
    output wire [3:0]                      M_AXIMM_113_AWREGION,
    output wire [3:0]                      M_AXIMM_113_AWQOS,
    output wire                            M_AXIMM_113_AWVALID,
    input  wire                            M_AXIMM_113_AWREADY,
    output wire [M_AXIMM_113_DATA_WIDTH-1:0]   M_AXIMM_113_WDATA,
    output wire [M_AXIMM_113_DATA_WIDTH/8-1:0] M_AXIMM_113_WSTRB,
    output wire                            M_AXIMM_113_WLAST,
    output wire                            M_AXIMM_113_WVALID,
    input  wire                            M_AXIMM_113_WREADY,
    input  wire [1:0]                      M_AXIMM_113_BRESP,
    input  wire                            M_AXIMM_113_BVALID,
    output wire                            M_AXIMM_113_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_113_ARADDR,
    output wire [7:0]                      M_AXIMM_113_ARLEN,
    output wire [2:0]                      M_AXIMM_113_ARSIZE,
    output wire [1:0]                      M_AXIMM_113_ARBURST,
    output wire [1:0]                      M_AXIMM_113_ARLOCK,
    output wire [3:0]                      M_AXIMM_113_ARCACHE,
    output wire [2:0]                      M_AXIMM_113_ARPROT,
    output wire [3:0]                      M_AXIMM_113_ARREGION,
    output wire [3:0]                      M_AXIMM_113_ARQOS,
    output wire                            M_AXIMM_113_ARVALID,
    input  wire                            M_AXIMM_113_ARREADY,
    input  wire [M_AXIMM_113_DATA_WIDTH-1:0]   M_AXIMM_113_RDATA,
    input  wire [1:0]                      M_AXIMM_113_RRESP,
    input  wire                            M_AXIMM_113_RLAST,
    input  wire                            M_AXIMM_113_RVALID,
    output wire                            M_AXIMM_113_RREADY,
    //AXI-MM pass-through interface 114
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_114_AWADDR,
    input wire [7:0]                      AP_AXIMM_114_AWLEN,
    input wire [2:0]                      AP_AXIMM_114_AWSIZE,
    input wire [1:0]                      AP_AXIMM_114_AWBURST,
    input wire [1:0]                      AP_AXIMM_114_AWLOCK,
    input wire [3:0]                      AP_AXIMM_114_AWCACHE,
    input wire [2:0]                      AP_AXIMM_114_AWPROT,
    input wire [3:0]                      AP_AXIMM_114_AWREGION,
    input wire [3:0]                      AP_AXIMM_114_AWQOS,
    input wire                            AP_AXIMM_114_AWVALID,
    output  wire                            AP_AXIMM_114_AWREADY,
    input wire [M_AXIMM_114_DATA_WIDTH-1:0]   AP_AXIMM_114_WDATA,
    input wire [M_AXIMM_114_DATA_WIDTH/8-1:0] AP_AXIMM_114_WSTRB,
    input wire                            AP_AXIMM_114_WLAST,
    input wire                            AP_AXIMM_114_WVALID,
    output  wire                            AP_AXIMM_114_WREADY,
    output  wire [1:0]                      AP_AXIMM_114_BRESP,
    output  wire                            AP_AXIMM_114_BVALID,
    input wire                            AP_AXIMM_114_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_114_ARADDR,
    input wire [7:0]                      AP_AXIMM_114_ARLEN,
    input wire [2:0]                      AP_AXIMM_114_ARSIZE,
    input wire [1:0]                      AP_AXIMM_114_ARBURST,
    input wire [1:0]                      AP_AXIMM_114_ARLOCK,
    input wire [3:0]                      AP_AXIMM_114_ARCACHE,
    input wire [2:0]                      AP_AXIMM_114_ARPROT,
    input wire [3:0]                      AP_AXIMM_114_ARREGION,
    input wire [3:0]                      AP_AXIMM_114_ARQOS,
    input wire                            AP_AXIMM_114_ARVALID,
    output  wire                            AP_AXIMM_114_ARREADY,
    output  wire [M_AXIMM_114_DATA_WIDTH-1:0]   AP_AXIMM_114_RDATA,
    output  wire [1:0]                      AP_AXIMM_114_RRESP,
    output  wire                            AP_AXIMM_114_RLAST,
    output  wire                            AP_AXIMM_114_RVALID,
    input  wire                            AP_AXIMM_114_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_114_AWADDR,
    output wire [7:0]                      M_AXIMM_114_AWLEN,
    output wire [2:0]                      M_AXIMM_114_AWSIZE,
    output wire [1:0]                      M_AXIMM_114_AWBURST,
    output wire [1:0]                      M_AXIMM_114_AWLOCK,
    output wire [3:0]                      M_AXIMM_114_AWCACHE,
    output wire [2:0]                      M_AXIMM_114_AWPROT,
    output wire [3:0]                      M_AXIMM_114_AWREGION,
    output wire [3:0]                      M_AXIMM_114_AWQOS,
    output wire                            M_AXIMM_114_AWVALID,
    input  wire                            M_AXIMM_114_AWREADY,
    output wire [M_AXIMM_114_DATA_WIDTH-1:0]   M_AXIMM_114_WDATA,
    output wire [M_AXIMM_114_DATA_WIDTH/8-1:0] M_AXIMM_114_WSTRB,
    output wire                            M_AXIMM_114_WLAST,
    output wire                            M_AXIMM_114_WVALID,
    input  wire                            M_AXIMM_114_WREADY,
    input  wire [1:0]                      M_AXIMM_114_BRESP,
    input  wire                            M_AXIMM_114_BVALID,
    output wire                            M_AXIMM_114_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_114_ARADDR,
    output wire [7:0]                      M_AXIMM_114_ARLEN,
    output wire [2:0]                      M_AXIMM_114_ARSIZE,
    output wire [1:0]                      M_AXIMM_114_ARBURST,
    output wire [1:0]                      M_AXIMM_114_ARLOCK,
    output wire [3:0]                      M_AXIMM_114_ARCACHE,
    output wire [2:0]                      M_AXIMM_114_ARPROT,
    output wire [3:0]                      M_AXIMM_114_ARREGION,
    output wire [3:0]                      M_AXIMM_114_ARQOS,
    output wire                            M_AXIMM_114_ARVALID,
    input  wire                            M_AXIMM_114_ARREADY,
    input  wire [M_AXIMM_114_DATA_WIDTH-1:0]   M_AXIMM_114_RDATA,
    input  wire [1:0]                      M_AXIMM_114_RRESP,
    input  wire                            M_AXIMM_114_RLAST,
    input  wire                            M_AXIMM_114_RVALID,
    output wire                            M_AXIMM_114_RREADY,
    //AXI-MM pass-through interface 115
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_115_AWADDR,
    input wire [7:0]                      AP_AXIMM_115_AWLEN,
    input wire [2:0]                      AP_AXIMM_115_AWSIZE,
    input wire [1:0]                      AP_AXIMM_115_AWBURST,
    input wire [1:0]                      AP_AXIMM_115_AWLOCK,
    input wire [3:0]                      AP_AXIMM_115_AWCACHE,
    input wire [2:0]                      AP_AXIMM_115_AWPROT,
    input wire [3:0]                      AP_AXIMM_115_AWREGION,
    input wire [3:0]                      AP_AXIMM_115_AWQOS,
    input wire                            AP_AXIMM_115_AWVALID,
    output  wire                            AP_AXIMM_115_AWREADY,
    input wire [M_AXIMM_115_DATA_WIDTH-1:0]   AP_AXIMM_115_WDATA,
    input wire [M_AXIMM_115_DATA_WIDTH/8-1:0] AP_AXIMM_115_WSTRB,
    input wire                            AP_AXIMM_115_WLAST,
    input wire                            AP_AXIMM_115_WVALID,
    output  wire                            AP_AXIMM_115_WREADY,
    output  wire [1:0]                      AP_AXIMM_115_BRESP,
    output  wire                            AP_AXIMM_115_BVALID,
    input wire                            AP_AXIMM_115_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_115_ARADDR,
    input wire [7:0]                      AP_AXIMM_115_ARLEN,
    input wire [2:0]                      AP_AXIMM_115_ARSIZE,
    input wire [1:0]                      AP_AXIMM_115_ARBURST,
    input wire [1:0]                      AP_AXIMM_115_ARLOCK,
    input wire [3:0]                      AP_AXIMM_115_ARCACHE,
    input wire [2:0]                      AP_AXIMM_115_ARPROT,
    input wire [3:0]                      AP_AXIMM_115_ARREGION,
    input wire [3:0]                      AP_AXIMM_115_ARQOS,
    input wire                            AP_AXIMM_115_ARVALID,
    output  wire                            AP_AXIMM_115_ARREADY,
    output  wire [M_AXIMM_115_DATA_WIDTH-1:0]   AP_AXIMM_115_RDATA,
    output  wire [1:0]                      AP_AXIMM_115_RRESP,
    output  wire                            AP_AXIMM_115_RLAST,
    output  wire                            AP_AXIMM_115_RVALID,
    input  wire                            AP_AXIMM_115_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_115_AWADDR,
    output wire [7:0]                      M_AXIMM_115_AWLEN,
    output wire [2:0]                      M_AXIMM_115_AWSIZE,
    output wire [1:0]                      M_AXIMM_115_AWBURST,
    output wire [1:0]                      M_AXIMM_115_AWLOCK,
    output wire [3:0]                      M_AXIMM_115_AWCACHE,
    output wire [2:0]                      M_AXIMM_115_AWPROT,
    output wire [3:0]                      M_AXIMM_115_AWREGION,
    output wire [3:0]                      M_AXIMM_115_AWQOS,
    output wire                            M_AXIMM_115_AWVALID,
    input  wire                            M_AXIMM_115_AWREADY,
    output wire [M_AXIMM_115_DATA_WIDTH-1:0]   M_AXIMM_115_WDATA,
    output wire [M_AXIMM_115_DATA_WIDTH/8-1:0] M_AXIMM_115_WSTRB,
    output wire                            M_AXIMM_115_WLAST,
    output wire                            M_AXIMM_115_WVALID,
    input  wire                            M_AXIMM_115_WREADY,
    input  wire [1:0]                      M_AXIMM_115_BRESP,
    input  wire                            M_AXIMM_115_BVALID,
    output wire                            M_AXIMM_115_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_115_ARADDR,
    output wire [7:0]                      M_AXIMM_115_ARLEN,
    output wire [2:0]                      M_AXIMM_115_ARSIZE,
    output wire [1:0]                      M_AXIMM_115_ARBURST,
    output wire [1:0]                      M_AXIMM_115_ARLOCK,
    output wire [3:0]                      M_AXIMM_115_ARCACHE,
    output wire [2:0]                      M_AXIMM_115_ARPROT,
    output wire [3:0]                      M_AXIMM_115_ARREGION,
    output wire [3:0]                      M_AXIMM_115_ARQOS,
    output wire                            M_AXIMM_115_ARVALID,
    input  wire                            M_AXIMM_115_ARREADY,
    input  wire [M_AXIMM_115_DATA_WIDTH-1:0]   M_AXIMM_115_RDATA,
    input  wire [1:0]                      M_AXIMM_115_RRESP,
    input  wire                            M_AXIMM_115_RLAST,
    input  wire                            M_AXIMM_115_RVALID,
    output wire                            M_AXIMM_115_RREADY,
    //AXI-MM pass-through interface 116
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_116_AWADDR,
    input wire [7:0]                      AP_AXIMM_116_AWLEN,
    input wire [2:0]                      AP_AXIMM_116_AWSIZE,
    input wire [1:0]                      AP_AXIMM_116_AWBURST,
    input wire [1:0]                      AP_AXIMM_116_AWLOCK,
    input wire [3:0]                      AP_AXIMM_116_AWCACHE,
    input wire [2:0]                      AP_AXIMM_116_AWPROT,
    input wire [3:0]                      AP_AXIMM_116_AWREGION,
    input wire [3:0]                      AP_AXIMM_116_AWQOS,
    input wire                            AP_AXIMM_116_AWVALID,
    output  wire                            AP_AXIMM_116_AWREADY,
    input wire [M_AXIMM_116_DATA_WIDTH-1:0]   AP_AXIMM_116_WDATA,
    input wire [M_AXIMM_116_DATA_WIDTH/8-1:0] AP_AXIMM_116_WSTRB,
    input wire                            AP_AXIMM_116_WLAST,
    input wire                            AP_AXIMM_116_WVALID,
    output  wire                            AP_AXIMM_116_WREADY,
    output  wire [1:0]                      AP_AXIMM_116_BRESP,
    output  wire                            AP_AXIMM_116_BVALID,
    input wire                            AP_AXIMM_116_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_116_ARADDR,
    input wire [7:0]                      AP_AXIMM_116_ARLEN,
    input wire [2:0]                      AP_AXIMM_116_ARSIZE,
    input wire [1:0]                      AP_AXIMM_116_ARBURST,
    input wire [1:0]                      AP_AXIMM_116_ARLOCK,
    input wire [3:0]                      AP_AXIMM_116_ARCACHE,
    input wire [2:0]                      AP_AXIMM_116_ARPROT,
    input wire [3:0]                      AP_AXIMM_116_ARREGION,
    input wire [3:0]                      AP_AXIMM_116_ARQOS,
    input wire                            AP_AXIMM_116_ARVALID,
    output  wire                            AP_AXIMM_116_ARREADY,
    output  wire [M_AXIMM_116_DATA_WIDTH-1:0]   AP_AXIMM_116_RDATA,
    output  wire [1:0]                      AP_AXIMM_116_RRESP,
    output  wire                            AP_AXIMM_116_RLAST,
    output  wire                            AP_AXIMM_116_RVALID,
    input  wire                            AP_AXIMM_116_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_116_AWADDR,
    output wire [7:0]                      M_AXIMM_116_AWLEN,
    output wire [2:0]                      M_AXIMM_116_AWSIZE,
    output wire [1:0]                      M_AXIMM_116_AWBURST,
    output wire [1:0]                      M_AXIMM_116_AWLOCK,
    output wire [3:0]                      M_AXIMM_116_AWCACHE,
    output wire [2:0]                      M_AXIMM_116_AWPROT,
    output wire [3:0]                      M_AXIMM_116_AWREGION,
    output wire [3:0]                      M_AXIMM_116_AWQOS,
    output wire                            M_AXIMM_116_AWVALID,
    input  wire                            M_AXIMM_116_AWREADY,
    output wire [M_AXIMM_116_DATA_WIDTH-1:0]   M_AXIMM_116_WDATA,
    output wire [M_AXIMM_116_DATA_WIDTH/8-1:0] M_AXIMM_116_WSTRB,
    output wire                            M_AXIMM_116_WLAST,
    output wire                            M_AXIMM_116_WVALID,
    input  wire                            M_AXIMM_116_WREADY,
    input  wire [1:0]                      M_AXIMM_116_BRESP,
    input  wire                            M_AXIMM_116_BVALID,
    output wire                            M_AXIMM_116_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_116_ARADDR,
    output wire [7:0]                      M_AXIMM_116_ARLEN,
    output wire [2:0]                      M_AXIMM_116_ARSIZE,
    output wire [1:0]                      M_AXIMM_116_ARBURST,
    output wire [1:0]                      M_AXIMM_116_ARLOCK,
    output wire [3:0]                      M_AXIMM_116_ARCACHE,
    output wire [2:0]                      M_AXIMM_116_ARPROT,
    output wire [3:0]                      M_AXIMM_116_ARREGION,
    output wire [3:0]                      M_AXIMM_116_ARQOS,
    output wire                            M_AXIMM_116_ARVALID,
    input  wire                            M_AXIMM_116_ARREADY,
    input  wire [M_AXIMM_116_DATA_WIDTH-1:0]   M_AXIMM_116_RDATA,
    input  wire [1:0]                      M_AXIMM_116_RRESP,
    input  wire                            M_AXIMM_116_RLAST,
    input  wire                            M_AXIMM_116_RVALID,
    output wire                            M_AXIMM_116_RREADY,
    //AXI-MM pass-through interface 117
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_117_AWADDR,
    input wire [7:0]                      AP_AXIMM_117_AWLEN,
    input wire [2:0]                      AP_AXIMM_117_AWSIZE,
    input wire [1:0]                      AP_AXIMM_117_AWBURST,
    input wire [1:0]                      AP_AXIMM_117_AWLOCK,
    input wire [3:0]                      AP_AXIMM_117_AWCACHE,
    input wire [2:0]                      AP_AXIMM_117_AWPROT,
    input wire [3:0]                      AP_AXIMM_117_AWREGION,
    input wire [3:0]                      AP_AXIMM_117_AWQOS,
    input wire                            AP_AXIMM_117_AWVALID,
    output  wire                            AP_AXIMM_117_AWREADY,
    input wire [M_AXIMM_117_DATA_WIDTH-1:0]   AP_AXIMM_117_WDATA,
    input wire [M_AXIMM_117_DATA_WIDTH/8-1:0] AP_AXIMM_117_WSTRB,
    input wire                            AP_AXIMM_117_WLAST,
    input wire                            AP_AXIMM_117_WVALID,
    output  wire                            AP_AXIMM_117_WREADY,
    output  wire [1:0]                      AP_AXIMM_117_BRESP,
    output  wire                            AP_AXIMM_117_BVALID,
    input wire                            AP_AXIMM_117_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_117_ARADDR,
    input wire [7:0]                      AP_AXIMM_117_ARLEN,
    input wire [2:0]                      AP_AXIMM_117_ARSIZE,
    input wire [1:0]                      AP_AXIMM_117_ARBURST,
    input wire [1:0]                      AP_AXIMM_117_ARLOCK,
    input wire [3:0]                      AP_AXIMM_117_ARCACHE,
    input wire [2:0]                      AP_AXIMM_117_ARPROT,
    input wire [3:0]                      AP_AXIMM_117_ARREGION,
    input wire [3:0]                      AP_AXIMM_117_ARQOS,
    input wire                            AP_AXIMM_117_ARVALID,
    output  wire                            AP_AXIMM_117_ARREADY,
    output  wire [M_AXIMM_117_DATA_WIDTH-1:0]   AP_AXIMM_117_RDATA,
    output  wire [1:0]                      AP_AXIMM_117_RRESP,
    output  wire                            AP_AXIMM_117_RLAST,
    output  wire                            AP_AXIMM_117_RVALID,
    input  wire                            AP_AXIMM_117_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_117_AWADDR,
    output wire [7:0]                      M_AXIMM_117_AWLEN,
    output wire [2:0]                      M_AXIMM_117_AWSIZE,
    output wire [1:0]                      M_AXIMM_117_AWBURST,
    output wire [1:0]                      M_AXIMM_117_AWLOCK,
    output wire [3:0]                      M_AXIMM_117_AWCACHE,
    output wire [2:0]                      M_AXIMM_117_AWPROT,
    output wire [3:0]                      M_AXIMM_117_AWREGION,
    output wire [3:0]                      M_AXIMM_117_AWQOS,
    output wire                            M_AXIMM_117_AWVALID,
    input  wire                            M_AXIMM_117_AWREADY,
    output wire [M_AXIMM_117_DATA_WIDTH-1:0]   M_AXIMM_117_WDATA,
    output wire [M_AXIMM_117_DATA_WIDTH/8-1:0] M_AXIMM_117_WSTRB,
    output wire                            M_AXIMM_117_WLAST,
    output wire                            M_AXIMM_117_WVALID,
    input  wire                            M_AXIMM_117_WREADY,
    input  wire [1:0]                      M_AXIMM_117_BRESP,
    input  wire                            M_AXIMM_117_BVALID,
    output wire                            M_AXIMM_117_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_117_ARADDR,
    output wire [7:0]                      M_AXIMM_117_ARLEN,
    output wire [2:0]                      M_AXIMM_117_ARSIZE,
    output wire [1:0]                      M_AXIMM_117_ARBURST,
    output wire [1:0]                      M_AXIMM_117_ARLOCK,
    output wire [3:0]                      M_AXIMM_117_ARCACHE,
    output wire [2:0]                      M_AXIMM_117_ARPROT,
    output wire [3:0]                      M_AXIMM_117_ARREGION,
    output wire [3:0]                      M_AXIMM_117_ARQOS,
    output wire                            M_AXIMM_117_ARVALID,
    input  wire                            M_AXIMM_117_ARREADY,
    input  wire [M_AXIMM_117_DATA_WIDTH-1:0]   M_AXIMM_117_RDATA,
    input  wire [1:0]                      M_AXIMM_117_RRESP,
    input  wire                            M_AXIMM_117_RLAST,
    input  wire                            M_AXIMM_117_RVALID,
    output wire                            M_AXIMM_117_RREADY,
    //AXI-MM pass-through interface 118
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_118_AWADDR,
    input wire [7:0]                      AP_AXIMM_118_AWLEN,
    input wire [2:0]                      AP_AXIMM_118_AWSIZE,
    input wire [1:0]                      AP_AXIMM_118_AWBURST,
    input wire [1:0]                      AP_AXIMM_118_AWLOCK,
    input wire [3:0]                      AP_AXIMM_118_AWCACHE,
    input wire [2:0]                      AP_AXIMM_118_AWPROT,
    input wire [3:0]                      AP_AXIMM_118_AWREGION,
    input wire [3:0]                      AP_AXIMM_118_AWQOS,
    input wire                            AP_AXIMM_118_AWVALID,
    output  wire                            AP_AXIMM_118_AWREADY,
    input wire [M_AXIMM_118_DATA_WIDTH-1:0]   AP_AXIMM_118_WDATA,
    input wire [M_AXIMM_118_DATA_WIDTH/8-1:0] AP_AXIMM_118_WSTRB,
    input wire                            AP_AXIMM_118_WLAST,
    input wire                            AP_AXIMM_118_WVALID,
    output  wire                            AP_AXIMM_118_WREADY,
    output  wire [1:0]                      AP_AXIMM_118_BRESP,
    output  wire                            AP_AXIMM_118_BVALID,
    input wire                            AP_AXIMM_118_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_118_ARADDR,
    input wire [7:0]                      AP_AXIMM_118_ARLEN,
    input wire [2:0]                      AP_AXIMM_118_ARSIZE,
    input wire [1:0]                      AP_AXIMM_118_ARBURST,
    input wire [1:0]                      AP_AXIMM_118_ARLOCK,
    input wire [3:0]                      AP_AXIMM_118_ARCACHE,
    input wire [2:0]                      AP_AXIMM_118_ARPROT,
    input wire [3:0]                      AP_AXIMM_118_ARREGION,
    input wire [3:0]                      AP_AXIMM_118_ARQOS,
    input wire                            AP_AXIMM_118_ARVALID,
    output  wire                            AP_AXIMM_118_ARREADY,
    output  wire [M_AXIMM_118_DATA_WIDTH-1:0]   AP_AXIMM_118_RDATA,
    output  wire [1:0]                      AP_AXIMM_118_RRESP,
    output  wire                            AP_AXIMM_118_RLAST,
    output  wire                            AP_AXIMM_118_RVALID,
    input  wire                            AP_AXIMM_118_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_118_AWADDR,
    output wire [7:0]                      M_AXIMM_118_AWLEN,
    output wire [2:0]                      M_AXIMM_118_AWSIZE,
    output wire [1:0]                      M_AXIMM_118_AWBURST,
    output wire [1:0]                      M_AXIMM_118_AWLOCK,
    output wire [3:0]                      M_AXIMM_118_AWCACHE,
    output wire [2:0]                      M_AXIMM_118_AWPROT,
    output wire [3:0]                      M_AXIMM_118_AWREGION,
    output wire [3:0]                      M_AXIMM_118_AWQOS,
    output wire                            M_AXIMM_118_AWVALID,
    input  wire                            M_AXIMM_118_AWREADY,
    output wire [M_AXIMM_118_DATA_WIDTH-1:0]   M_AXIMM_118_WDATA,
    output wire [M_AXIMM_118_DATA_WIDTH/8-1:0] M_AXIMM_118_WSTRB,
    output wire                            M_AXIMM_118_WLAST,
    output wire                            M_AXIMM_118_WVALID,
    input  wire                            M_AXIMM_118_WREADY,
    input  wire [1:0]                      M_AXIMM_118_BRESP,
    input  wire                            M_AXIMM_118_BVALID,
    output wire                            M_AXIMM_118_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_118_ARADDR,
    output wire [7:0]                      M_AXIMM_118_ARLEN,
    output wire [2:0]                      M_AXIMM_118_ARSIZE,
    output wire [1:0]                      M_AXIMM_118_ARBURST,
    output wire [1:0]                      M_AXIMM_118_ARLOCK,
    output wire [3:0]                      M_AXIMM_118_ARCACHE,
    output wire [2:0]                      M_AXIMM_118_ARPROT,
    output wire [3:0]                      M_AXIMM_118_ARREGION,
    output wire [3:0]                      M_AXIMM_118_ARQOS,
    output wire                            M_AXIMM_118_ARVALID,
    input  wire                            M_AXIMM_118_ARREADY,
    input  wire [M_AXIMM_118_DATA_WIDTH-1:0]   M_AXIMM_118_RDATA,
    input  wire [1:0]                      M_AXIMM_118_RRESP,
    input  wire                            M_AXIMM_118_RLAST,
    input  wire                            M_AXIMM_118_RVALID,
    output wire                            M_AXIMM_118_RREADY,
    //AXI-MM pass-through interface 119
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_119_AWADDR,
    input wire [7:0]                      AP_AXIMM_119_AWLEN,
    input wire [2:0]                      AP_AXIMM_119_AWSIZE,
    input wire [1:0]                      AP_AXIMM_119_AWBURST,
    input wire [1:0]                      AP_AXIMM_119_AWLOCK,
    input wire [3:0]                      AP_AXIMM_119_AWCACHE,
    input wire [2:0]                      AP_AXIMM_119_AWPROT,
    input wire [3:0]                      AP_AXIMM_119_AWREGION,
    input wire [3:0]                      AP_AXIMM_119_AWQOS,
    input wire                            AP_AXIMM_119_AWVALID,
    output  wire                            AP_AXIMM_119_AWREADY,
    input wire [M_AXIMM_119_DATA_WIDTH-1:0]   AP_AXIMM_119_WDATA,
    input wire [M_AXIMM_119_DATA_WIDTH/8-1:0] AP_AXIMM_119_WSTRB,
    input wire                            AP_AXIMM_119_WLAST,
    input wire                            AP_AXIMM_119_WVALID,
    output  wire                            AP_AXIMM_119_WREADY,
    output  wire [1:0]                      AP_AXIMM_119_BRESP,
    output  wire                            AP_AXIMM_119_BVALID,
    input wire                            AP_AXIMM_119_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_119_ARADDR,
    input wire [7:0]                      AP_AXIMM_119_ARLEN,
    input wire [2:0]                      AP_AXIMM_119_ARSIZE,
    input wire [1:0]                      AP_AXIMM_119_ARBURST,
    input wire [1:0]                      AP_AXIMM_119_ARLOCK,
    input wire [3:0]                      AP_AXIMM_119_ARCACHE,
    input wire [2:0]                      AP_AXIMM_119_ARPROT,
    input wire [3:0]                      AP_AXIMM_119_ARREGION,
    input wire [3:0]                      AP_AXIMM_119_ARQOS,
    input wire                            AP_AXIMM_119_ARVALID,
    output  wire                            AP_AXIMM_119_ARREADY,
    output  wire [M_AXIMM_119_DATA_WIDTH-1:0]   AP_AXIMM_119_RDATA,
    output  wire [1:0]                      AP_AXIMM_119_RRESP,
    output  wire                            AP_AXIMM_119_RLAST,
    output  wire                            AP_AXIMM_119_RVALID,
    input  wire                            AP_AXIMM_119_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_119_AWADDR,
    output wire [7:0]                      M_AXIMM_119_AWLEN,
    output wire [2:0]                      M_AXIMM_119_AWSIZE,
    output wire [1:0]                      M_AXIMM_119_AWBURST,
    output wire [1:0]                      M_AXIMM_119_AWLOCK,
    output wire [3:0]                      M_AXIMM_119_AWCACHE,
    output wire [2:0]                      M_AXIMM_119_AWPROT,
    output wire [3:0]                      M_AXIMM_119_AWREGION,
    output wire [3:0]                      M_AXIMM_119_AWQOS,
    output wire                            M_AXIMM_119_AWVALID,
    input  wire                            M_AXIMM_119_AWREADY,
    output wire [M_AXIMM_119_DATA_WIDTH-1:0]   M_AXIMM_119_WDATA,
    output wire [M_AXIMM_119_DATA_WIDTH/8-1:0] M_AXIMM_119_WSTRB,
    output wire                            M_AXIMM_119_WLAST,
    output wire                            M_AXIMM_119_WVALID,
    input  wire                            M_AXIMM_119_WREADY,
    input  wire [1:0]                      M_AXIMM_119_BRESP,
    input  wire                            M_AXIMM_119_BVALID,
    output wire                            M_AXIMM_119_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_119_ARADDR,
    output wire [7:0]                      M_AXIMM_119_ARLEN,
    output wire [2:0]                      M_AXIMM_119_ARSIZE,
    output wire [1:0]                      M_AXIMM_119_ARBURST,
    output wire [1:0]                      M_AXIMM_119_ARLOCK,
    output wire [3:0]                      M_AXIMM_119_ARCACHE,
    output wire [2:0]                      M_AXIMM_119_ARPROT,
    output wire [3:0]                      M_AXIMM_119_ARREGION,
    output wire [3:0]                      M_AXIMM_119_ARQOS,
    output wire                            M_AXIMM_119_ARVALID,
    input  wire                            M_AXIMM_119_ARREADY,
    input  wire [M_AXIMM_119_DATA_WIDTH-1:0]   M_AXIMM_119_RDATA,
    input  wire [1:0]                      M_AXIMM_119_RRESP,
    input  wire                            M_AXIMM_119_RLAST,
    input  wire                            M_AXIMM_119_RVALID,
    output wire                            M_AXIMM_119_RREADY,
    //AXI-MM pass-through interface 120
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_120_AWADDR,
    input wire [7:0]                      AP_AXIMM_120_AWLEN,
    input wire [2:0]                      AP_AXIMM_120_AWSIZE,
    input wire [1:0]                      AP_AXIMM_120_AWBURST,
    input wire [1:0]                      AP_AXIMM_120_AWLOCK,
    input wire [3:0]                      AP_AXIMM_120_AWCACHE,
    input wire [2:0]                      AP_AXIMM_120_AWPROT,
    input wire [3:0]                      AP_AXIMM_120_AWREGION,
    input wire [3:0]                      AP_AXIMM_120_AWQOS,
    input wire                            AP_AXIMM_120_AWVALID,
    output  wire                            AP_AXIMM_120_AWREADY,
    input wire [M_AXIMM_120_DATA_WIDTH-1:0]   AP_AXIMM_120_WDATA,
    input wire [M_AXIMM_120_DATA_WIDTH/8-1:0] AP_AXIMM_120_WSTRB,
    input wire                            AP_AXIMM_120_WLAST,
    input wire                            AP_AXIMM_120_WVALID,
    output  wire                            AP_AXIMM_120_WREADY,
    output  wire [1:0]                      AP_AXIMM_120_BRESP,
    output  wire                            AP_AXIMM_120_BVALID,
    input wire                            AP_AXIMM_120_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_120_ARADDR,
    input wire [7:0]                      AP_AXIMM_120_ARLEN,
    input wire [2:0]                      AP_AXIMM_120_ARSIZE,
    input wire [1:0]                      AP_AXIMM_120_ARBURST,
    input wire [1:0]                      AP_AXIMM_120_ARLOCK,
    input wire [3:0]                      AP_AXIMM_120_ARCACHE,
    input wire [2:0]                      AP_AXIMM_120_ARPROT,
    input wire [3:0]                      AP_AXIMM_120_ARREGION,
    input wire [3:0]                      AP_AXIMM_120_ARQOS,
    input wire                            AP_AXIMM_120_ARVALID,
    output  wire                            AP_AXIMM_120_ARREADY,
    output  wire [M_AXIMM_120_DATA_WIDTH-1:0]   AP_AXIMM_120_RDATA,
    output  wire [1:0]                      AP_AXIMM_120_RRESP,
    output  wire                            AP_AXIMM_120_RLAST,
    output  wire                            AP_AXIMM_120_RVALID,
    input  wire                            AP_AXIMM_120_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_120_AWADDR,
    output wire [7:0]                      M_AXIMM_120_AWLEN,
    output wire [2:0]                      M_AXIMM_120_AWSIZE,
    output wire [1:0]                      M_AXIMM_120_AWBURST,
    output wire [1:0]                      M_AXIMM_120_AWLOCK,
    output wire [3:0]                      M_AXIMM_120_AWCACHE,
    output wire [2:0]                      M_AXIMM_120_AWPROT,
    output wire [3:0]                      M_AXIMM_120_AWREGION,
    output wire [3:0]                      M_AXIMM_120_AWQOS,
    output wire                            M_AXIMM_120_AWVALID,
    input  wire                            M_AXIMM_120_AWREADY,
    output wire [M_AXIMM_120_DATA_WIDTH-1:0]   M_AXIMM_120_WDATA,
    output wire [M_AXIMM_120_DATA_WIDTH/8-1:0] M_AXIMM_120_WSTRB,
    output wire                            M_AXIMM_120_WLAST,
    output wire                            M_AXIMM_120_WVALID,
    input  wire                            M_AXIMM_120_WREADY,
    input  wire [1:0]                      M_AXIMM_120_BRESP,
    input  wire                            M_AXIMM_120_BVALID,
    output wire                            M_AXIMM_120_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_120_ARADDR,
    output wire [7:0]                      M_AXIMM_120_ARLEN,
    output wire [2:0]                      M_AXIMM_120_ARSIZE,
    output wire [1:0]                      M_AXIMM_120_ARBURST,
    output wire [1:0]                      M_AXIMM_120_ARLOCK,
    output wire [3:0]                      M_AXIMM_120_ARCACHE,
    output wire [2:0]                      M_AXIMM_120_ARPROT,
    output wire [3:0]                      M_AXIMM_120_ARREGION,
    output wire [3:0]                      M_AXIMM_120_ARQOS,
    output wire                            M_AXIMM_120_ARVALID,
    input  wire                            M_AXIMM_120_ARREADY,
    input  wire [M_AXIMM_120_DATA_WIDTH-1:0]   M_AXIMM_120_RDATA,
    input  wire [1:0]                      M_AXIMM_120_RRESP,
    input  wire                            M_AXIMM_120_RLAST,
    input  wire                            M_AXIMM_120_RVALID,
    output wire                            M_AXIMM_120_RREADY,
    //AXI-MM pass-through interface 121
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_121_AWADDR,
    input wire [7:0]                      AP_AXIMM_121_AWLEN,
    input wire [2:0]                      AP_AXIMM_121_AWSIZE,
    input wire [1:0]                      AP_AXIMM_121_AWBURST,
    input wire [1:0]                      AP_AXIMM_121_AWLOCK,
    input wire [3:0]                      AP_AXIMM_121_AWCACHE,
    input wire [2:0]                      AP_AXIMM_121_AWPROT,
    input wire [3:0]                      AP_AXIMM_121_AWREGION,
    input wire [3:0]                      AP_AXIMM_121_AWQOS,
    input wire                            AP_AXIMM_121_AWVALID,
    output  wire                            AP_AXIMM_121_AWREADY,
    input wire [M_AXIMM_121_DATA_WIDTH-1:0]   AP_AXIMM_121_WDATA,
    input wire [M_AXIMM_121_DATA_WIDTH/8-1:0] AP_AXIMM_121_WSTRB,
    input wire                            AP_AXIMM_121_WLAST,
    input wire                            AP_AXIMM_121_WVALID,
    output  wire                            AP_AXIMM_121_WREADY,
    output  wire [1:0]                      AP_AXIMM_121_BRESP,
    output  wire                            AP_AXIMM_121_BVALID,
    input wire                            AP_AXIMM_121_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_121_ARADDR,
    input wire [7:0]                      AP_AXIMM_121_ARLEN,
    input wire [2:0]                      AP_AXIMM_121_ARSIZE,
    input wire [1:0]                      AP_AXIMM_121_ARBURST,
    input wire [1:0]                      AP_AXIMM_121_ARLOCK,
    input wire [3:0]                      AP_AXIMM_121_ARCACHE,
    input wire [2:0]                      AP_AXIMM_121_ARPROT,
    input wire [3:0]                      AP_AXIMM_121_ARREGION,
    input wire [3:0]                      AP_AXIMM_121_ARQOS,
    input wire                            AP_AXIMM_121_ARVALID,
    output  wire                            AP_AXIMM_121_ARREADY,
    output  wire [M_AXIMM_121_DATA_WIDTH-1:0]   AP_AXIMM_121_RDATA,
    output  wire [1:0]                      AP_AXIMM_121_RRESP,
    output  wire                            AP_AXIMM_121_RLAST,
    output  wire                            AP_AXIMM_121_RVALID,
    input  wire                            AP_AXIMM_121_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_121_AWADDR,
    output wire [7:0]                      M_AXIMM_121_AWLEN,
    output wire [2:0]                      M_AXIMM_121_AWSIZE,
    output wire [1:0]                      M_AXIMM_121_AWBURST,
    output wire [1:0]                      M_AXIMM_121_AWLOCK,
    output wire [3:0]                      M_AXIMM_121_AWCACHE,
    output wire [2:0]                      M_AXIMM_121_AWPROT,
    output wire [3:0]                      M_AXIMM_121_AWREGION,
    output wire [3:0]                      M_AXIMM_121_AWQOS,
    output wire                            M_AXIMM_121_AWVALID,
    input  wire                            M_AXIMM_121_AWREADY,
    output wire [M_AXIMM_121_DATA_WIDTH-1:0]   M_AXIMM_121_WDATA,
    output wire [M_AXIMM_121_DATA_WIDTH/8-1:0] M_AXIMM_121_WSTRB,
    output wire                            M_AXIMM_121_WLAST,
    output wire                            M_AXIMM_121_WVALID,
    input  wire                            M_AXIMM_121_WREADY,
    input  wire [1:0]                      M_AXIMM_121_BRESP,
    input  wire                            M_AXIMM_121_BVALID,
    output wire                            M_AXIMM_121_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_121_ARADDR,
    output wire [7:0]                      M_AXIMM_121_ARLEN,
    output wire [2:0]                      M_AXIMM_121_ARSIZE,
    output wire [1:0]                      M_AXIMM_121_ARBURST,
    output wire [1:0]                      M_AXIMM_121_ARLOCK,
    output wire [3:0]                      M_AXIMM_121_ARCACHE,
    output wire [2:0]                      M_AXIMM_121_ARPROT,
    output wire [3:0]                      M_AXIMM_121_ARREGION,
    output wire [3:0]                      M_AXIMM_121_ARQOS,
    output wire                            M_AXIMM_121_ARVALID,
    input  wire                            M_AXIMM_121_ARREADY,
    input  wire [M_AXIMM_121_DATA_WIDTH-1:0]   M_AXIMM_121_RDATA,
    input  wire [1:0]                      M_AXIMM_121_RRESP,
    input  wire                            M_AXIMM_121_RLAST,
    input  wire                            M_AXIMM_121_RVALID,
    output wire                            M_AXIMM_121_RREADY,
    //AXI-MM pass-through interface 122
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_122_AWADDR,
    input wire [7:0]                      AP_AXIMM_122_AWLEN,
    input wire [2:0]                      AP_AXIMM_122_AWSIZE,
    input wire [1:0]                      AP_AXIMM_122_AWBURST,
    input wire [1:0]                      AP_AXIMM_122_AWLOCK,
    input wire [3:0]                      AP_AXIMM_122_AWCACHE,
    input wire [2:0]                      AP_AXIMM_122_AWPROT,
    input wire [3:0]                      AP_AXIMM_122_AWREGION,
    input wire [3:0]                      AP_AXIMM_122_AWQOS,
    input wire                            AP_AXIMM_122_AWVALID,
    output  wire                            AP_AXIMM_122_AWREADY,
    input wire [M_AXIMM_122_DATA_WIDTH-1:0]   AP_AXIMM_122_WDATA,
    input wire [M_AXIMM_122_DATA_WIDTH/8-1:0] AP_AXIMM_122_WSTRB,
    input wire                            AP_AXIMM_122_WLAST,
    input wire                            AP_AXIMM_122_WVALID,
    output  wire                            AP_AXIMM_122_WREADY,
    output  wire [1:0]                      AP_AXIMM_122_BRESP,
    output  wire                            AP_AXIMM_122_BVALID,
    input wire                            AP_AXIMM_122_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_122_ARADDR,
    input wire [7:0]                      AP_AXIMM_122_ARLEN,
    input wire [2:0]                      AP_AXIMM_122_ARSIZE,
    input wire [1:0]                      AP_AXIMM_122_ARBURST,
    input wire [1:0]                      AP_AXIMM_122_ARLOCK,
    input wire [3:0]                      AP_AXIMM_122_ARCACHE,
    input wire [2:0]                      AP_AXIMM_122_ARPROT,
    input wire [3:0]                      AP_AXIMM_122_ARREGION,
    input wire [3:0]                      AP_AXIMM_122_ARQOS,
    input wire                            AP_AXIMM_122_ARVALID,
    output  wire                            AP_AXIMM_122_ARREADY,
    output  wire [M_AXIMM_122_DATA_WIDTH-1:0]   AP_AXIMM_122_RDATA,
    output  wire [1:0]                      AP_AXIMM_122_RRESP,
    output  wire                            AP_AXIMM_122_RLAST,
    output  wire                            AP_AXIMM_122_RVALID,
    input  wire                            AP_AXIMM_122_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_122_AWADDR,
    output wire [7:0]                      M_AXIMM_122_AWLEN,
    output wire [2:0]                      M_AXIMM_122_AWSIZE,
    output wire [1:0]                      M_AXIMM_122_AWBURST,
    output wire [1:0]                      M_AXIMM_122_AWLOCK,
    output wire [3:0]                      M_AXIMM_122_AWCACHE,
    output wire [2:0]                      M_AXIMM_122_AWPROT,
    output wire [3:0]                      M_AXIMM_122_AWREGION,
    output wire [3:0]                      M_AXIMM_122_AWQOS,
    output wire                            M_AXIMM_122_AWVALID,
    input  wire                            M_AXIMM_122_AWREADY,
    output wire [M_AXIMM_122_DATA_WIDTH-1:0]   M_AXIMM_122_WDATA,
    output wire [M_AXIMM_122_DATA_WIDTH/8-1:0] M_AXIMM_122_WSTRB,
    output wire                            M_AXIMM_122_WLAST,
    output wire                            M_AXIMM_122_WVALID,
    input  wire                            M_AXIMM_122_WREADY,
    input  wire [1:0]                      M_AXIMM_122_BRESP,
    input  wire                            M_AXIMM_122_BVALID,
    output wire                            M_AXIMM_122_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_122_ARADDR,
    output wire [7:0]                      M_AXIMM_122_ARLEN,
    output wire [2:0]                      M_AXIMM_122_ARSIZE,
    output wire [1:0]                      M_AXIMM_122_ARBURST,
    output wire [1:0]                      M_AXIMM_122_ARLOCK,
    output wire [3:0]                      M_AXIMM_122_ARCACHE,
    output wire [2:0]                      M_AXIMM_122_ARPROT,
    output wire [3:0]                      M_AXIMM_122_ARREGION,
    output wire [3:0]                      M_AXIMM_122_ARQOS,
    output wire                            M_AXIMM_122_ARVALID,
    input  wire                            M_AXIMM_122_ARREADY,
    input  wire [M_AXIMM_122_DATA_WIDTH-1:0]   M_AXIMM_122_RDATA,
    input  wire [1:0]                      M_AXIMM_122_RRESP,
    input  wire                            M_AXIMM_122_RLAST,
    input  wire                            M_AXIMM_122_RVALID,
    output wire                            M_AXIMM_122_RREADY,
    //AXI-MM pass-through interface 123
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_123_AWADDR,
    input wire [7:0]                      AP_AXIMM_123_AWLEN,
    input wire [2:0]                      AP_AXIMM_123_AWSIZE,
    input wire [1:0]                      AP_AXIMM_123_AWBURST,
    input wire [1:0]                      AP_AXIMM_123_AWLOCK,
    input wire [3:0]                      AP_AXIMM_123_AWCACHE,
    input wire [2:0]                      AP_AXIMM_123_AWPROT,
    input wire [3:0]                      AP_AXIMM_123_AWREGION,
    input wire [3:0]                      AP_AXIMM_123_AWQOS,
    input wire                            AP_AXIMM_123_AWVALID,
    output  wire                            AP_AXIMM_123_AWREADY,
    input wire [M_AXIMM_123_DATA_WIDTH-1:0]   AP_AXIMM_123_WDATA,
    input wire [M_AXIMM_123_DATA_WIDTH/8-1:0] AP_AXIMM_123_WSTRB,
    input wire                            AP_AXIMM_123_WLAST,
    input wire                            AP_AXIMM_123_WVALID,
    output  wire                            AP_AXIMM_123_WREADY,
    output  wire [1:0]                      AP_AXIMM_123_BRESP,
    output  wire                            AP_AXIMM_123_BVALID,
    input wire                            AP_AXIMM_123_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_123_ARADDR,
    input wire [7:0]                      AP_AXIMM_123_ARLEN,
    input wire [2:0]                      AP_AXIMM_123_ARSIZE,
    input wire [1:0]                      AP_AXIMM_123_ARBURST,
    input wire [1:0]                      AP_AXIMM_123_ARLOCK,
    input wire [3:0]                      AP_AXIMM_123_ARCACHE,
    input wire [2:0]                      AP_AXIMM_123_ARPROT,
    input wire [3:0]                      AP_AXIMM_123_ARREGION,
    input wire [3:0]                      AP_AXIMM_123_ARQOS,
    input wire                            AP_AXIMM_123_ARVALID,
    output  wire                            AP_AXIMM_123_ARREADY,
    output  wire [M_AXIMM_123_DATA_WIDTH-1:0]   AP_AXIMM_123_RDATA,
    output  wire [1:0]                      AP_AXIMM_123_RRESP,
    output  wire                            AP_AXIMM_123_RLAST,
    output  wire                            AP_AXIMM_123_RVALID,
    input  wire                            AP_AXIMM_123_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_123_AWADDR,
    output wire [7:0]                      M_AXIMM_123_AWLEN,
    output wire [2:0]                      M_AXIMM_123_AWSIZE,
    output wire [1:0]                      M_AXIMM_123_AWBURST,
    output wire [1:0]                      M_AXIMM_123_AWLOCK,
    output wire [3:0]                      M_AXIMM_123_AWCACHE,
    output wire [2:0]                      M_AXIMM_123_AWPROT,
    output wire [3:0]                      M_AXIMM_123_AWREGION,
    output wire [3:0]                      M_AXIMM_123_AWQOS,
    output wire                            M_AXIMM_123_AWVALID,
    input  wire                            M_AXIMM_123_AWREADY,
    output wire [M_AXIMM_123_DATA_WIDTH-1:0]   M_AXIMM_123_WDATA,
    output wire [M_AXIMM_123_DATA_WIDTH/8-1:0] M_AXIMM_123_WSTRB,
    output wire                            M_AXIMM_123_WLAST,
    output wire                            M_AXIMM_123_WVALID,
    input  wire                            M_AXIMM_123_WREADY,
    input  wire [1:0]                      M_AXIMM_123_BRESP,
    input  wire                            M_AXIMM_123_BVALID,
    output wire                            M_AXIMM_123_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_123_ARADDR,
    output wire [7:0]                      M_AXIMM_123_ARLEN,
    output wire [2:0]                      M_AXIMM_123_ARSIZE,
    output wire [1:0]                      M_AXIMM_123_ARBURST,
    output wire [1:0]                      M_AXIMM_123_ARLOCK,
    output wire [3:0]                      M_AXIMM_123_ARCACHE,
    output wire [2:0]                      M_AXIMM_123_ARPROT,
    output wire [3:0]                      M_AXIMM_123_ARREGION,
    output wire [3:0]                      M_AXIMM_123_ARQOS,
    output wire                            M_AXIMM_123_ARVALID,
    input  wire                            M_AXIMM_123_ARREADY,
    input  wire [M_AXIMM_123_DATA_WIDTH-1:0]   M_AXIMM_123_RDATA,
    input  wire [1:0]                      M_AXIMM_123_RRESP,
    input  wire                            M_AXIMM_123_RLAST,
    input  wire                            M_AXIMM_123_RVALID,
    output wire                            M_AXIMM_123_RREADY,
    //AXI-MM pass-through interface 124
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_124_AWADDR,
    input wire [7:0]                      AP_AXIMM_124_AWLEN,
    input wire [2:0]                      AP_AXIMM_124_AWSIZE,
    input wire [1:0]                      AP_AXIMM_124_AWBURST,
    input wire [1:0]                      AP_AXIMM_124_AWLOCK,
    input wire [3:0]                      AP_AXIMM_124_AWCACHE,
    input wire [2:0]                      AP_AXIMM_124_AWPROT,
    input wire [3:0]                      AP_AXIMM_124_AWREGION,
    input wire [3:0]                      AP_AXIMM_124_AWQOS,
    input wire                            AP_AXIMM_124_AWVALID,
    output  wire                            AP_AXIMM_124_AWREADY,
    input wire [M_AXIMM_124_DATA_WIDTH-1:0]   AP_AXIMM_124_WDATA,
    input wire [M_AXIMM_124_DATA_WIDTH/8-1:0] AP_AXIMM_124_WSTRB,
    input wire                            AP_AXIMM_124_WLAST,
    input wire                            AP_AXIMM_124_WVALID,
    output  wire                            AP_AXIMM_124_WREADY,
    output  wire [1:0]                      AP_AXIMM_124_BRESP,
    output  wire                            AP_AXIMM_124_BVALID,
    input wire                            AP_AXIMM_124_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_124_ARADDR,
    input wire [7:0]                      AP_AXIMM_124_ARLEN,
    input wire [2:0]                      AP_AXIMM_124_ARSIZE,
    input wire [1:0]                      AP_AXIMM_124_ARBURST,
    input wire [1:0]                      AP_AXIMM_124_ARLOCK,
    input wire [3:0]                      AP_AXIMM_124_ARCACHE,
    input wire [2:0]                      AP_AXIMM_124_ARPROT,
    input wire [3:0]                      AP_AXIMM_124_ARREGION,
    input wire [3:0]                      AP_AXIMM_124_ARQOS,
    input wire                            AP_AXIMM_124_ARVALID,
    output  wire                            AP_AXIMM_124_ARREADY,
    output  wire [M_AXIMM_124_DATA_WIDTH-1:0]   AP_AXIMM_124_RDATA,
    output  wire [1:0]                      AP_AXIMM_124_RRESP,
    output  wire                            AP_AXIMM_124_RLAST,
    output  wire                            AP_AXIMM_124_RVALID,
    input  wire                            AP_AXIMM_124_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_124_AWADDR,
    output wire [7:0]                      M_AXIMM_124_AWLEN,
    output wire [2:0]                      M_AXIMM_124_AWSIZE,
    output wire [1:0]                      M_AXIMM_124_AWBURST,
    output wire [1:0]                      M_AXIMM_124_AWLOCK,
    output wire [3:0]                      M_AXIMM_124_AWCACHE,
    output wire [2:0]                      M_AXIMM_124_AWPROT,
    output wire [3:0]                      M_AXIMM_124_AWREGION,
    output wire [3:0]                      M_AXIMM_124_AWQOS,
    output wire                            M_AXIMM_124_AWVALID,
    input  wire                            M_AXIMM_124_AWREADY,
    output wire [M_AXIMM_124_DATA_WIDTH-1:0]   M_AXIMM_124_WDATA,
    output wire [M_AXIMM_124_DATA_WIDTH/8-1:0] M_AXIMM_124_WSTRB,
    output wire                            M_AXIMM_124_WLAST,
    output wire                            M_AXIMM_124_WVALID,
    input  wire                            M_AXIMM_124_WREADY,
    input  wire [1:0]                      M_AXIMM_124_BRESP,
    input  wire                            M_AXIMM_124_BVALID,
    output wire                            M_AXIMM_124_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_124_ARADDR,
    output wire [7:0]                      M_AXIMM_124_ARLEN,
    output wire [2:0]                      M_AXIMM_124_ARSIZE,
    output wire [1:0]                      M_AXIMM_124_ARBURST,
    output wire [1:0]                      M_AXIMM_124_ARLOCK,
    output wire [3:0]                      M_AXIMM_124_ARCACHE,
    output wire [2:0]                      M_AXIMM_124_ARPROT,
    output wire [3:0]                      M_AXIMM_124_ARREGION,
    output wire [3:0]                      M_AXIMM_124_ARQOS,
    output wire                            M_AXIMM_124_ARVALID,
    input  wire                            M_AXIMM_124_ARREADY,
    input  wire [M_AXIMM_124_DATA_WIDTH-1:0]   M_AXIMM_124_RDATA,
    input  wire [1:0]                      M_AXIMM_124_RRESP,
    input  wire                            M_AXIMM_124_RLAST,
    input  wire                            M_AXIMM_124_RVALID,
    output wire                            M_AXIMM_124_RREADY,
    //AXI-MM pass-through interface 125
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_125_AWADDR,
    input wire [7:0]                      AP_AXIMM_125_AWLEN,
    input wire [2:0]                      AP_AXIMM_125_AWSIZE,
    input wire [1:0]                      AP_AXIMM_125_AWBURST,
    input wire [1:0]                      AP_AXIMM_125_AWLOCK,
    input wire [3:0]                      AP_AXIMM_125_AWCACHE,
    input wire [2:0]                      AP_AXIMM_125_AWPROT,
    input wire [3:0]                      AP_AXIMM_125_AWREGION,
    input wire [3:0]                      AP_AXIMM_125_AWQOS,
    input wire                            AP_AXIMM_125_AWVALID,
    output  wire                            AP_AXIMM_125_AWREADY,
    input wire [M_AXIMM_125_DATA_WIDTH-1:0]   AP_AXIMM_125_WDATA,
    input wire [M_AXIMM_125_DATA_WIDTH/8-1:0] AP_AXIMM_125_WSTRB,
    input wire                            AP_AXIMM_125_WLAST,
    input wire                            AP_AXIMM_125_WVALID,
    output  wire                            AP_AXIMM_125_WREADY,
    output  wire [1:0]                      AP_AXIMM_125_BRESP,
    output  wire                            AP_AXIMM_125_BVALID,
    input wire                            AP_AXIMM_125_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_125_ARADDR,
    input wire [7:0]                      AP_AXIMM_125_ARLEN,
    input wire [2:0]                      AP_AXIMM_125_ARSIZE,
    input wire [1:0]                      AP_AXIMM_125_ARBURST,
    input wire [1:0]                      AP_AXIMM_125_ARLOCK,
    input wire [3:0]                      AP_AXIMM_125_ARCACHE,
    input wire [2:0]                      AP_AXIMM_125_ARPROT,
    input wire [3:0]                      AP_AXIMM_125_ARREGION,
    input wire [3:0]                      AP_AXIMM_125_ARQOS,
    input wire                            AP_AXIMM_125_ARVALID,
    output  wire                            AP_AXIMM_125_ARREADY,
    output  wire [M_AXIMM_125_DATA_WIDTH-1:0]   AP_AXIMM_125_RDATA,
    output  wire [1:0]                      AP_AXIMM_125_RRESP,
    output  wire                            AP_AXIMM_125_RLAST,
    output  wire                            AP_AXIMM_125_RVALID,
    input  wire                            AP_AXIMM_125_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_125_AWADDR,
    output wire [7:0]                      M_AXIMM_125_AWLEN,
    output wire [2:0]                      M_AXIMM_125_AWSIZE,
    output wire [1:0]                      M_AXIMM_125_AWBURST,
    output wire [1:0]                      M_AXIMM_125_AWLOCK,
    output wire [3:0]                      M_AXIMM_125_AWCACHE,
    output wire [2:0]                      M_AXIMM_125_AWPROT,
    output wire [3:0]                      M_AXIMM_125_AWREGION,
    output wire [3:0]                      M_AXIMM_125_AWQOS,
    output wire                            M_AXIMM_125_AWVALID,
    input  wire                            M_AXIMM_125_AWREADY,
    output wire [M_AXIMM_125_DATA_WIDTH-1:0]   M_AXIMM_125_WDATA,
    output wire [M_AXIMM_125_DATA_WIDTH/8-1:0] M_AXIMM_125_WSTRB,
    output wire                            M_AXIMM_125_WLAST,
    output wire                            M_AXIMM_125_WVALID,
    input  wire                            M_AXIMM_125_WREADY,
    input  wire [1:0]                      M_AXIMM_125_BRESP,
    input  wire                            M_AXIMM_125_BVALID,
    output wire                            M_AXIMM_125_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_125_ARADDR,
    output wire [7:0]                      M_AXIMM_125_ARLEN,
    output wire [2:0]                      M_AXIMM_125_ARSIZE,
    output wire [1:0]                      M_AXIMM_125_ARBURST,
    output wire [1:0]                      M_AXIMM_125_ARLOCK,
    output wire [3:0]                      M_AXIMM_125_ARCACHE,
    output wire [2:0]                      M_AXIMM_125_ARPROT,
    output wire [3:0]                      M_AXIMM_125_ARREGION,
    output wire [3:0]                      M_AXIMM_125_ARQOS,
    output wire                            M_AXIMM_125_ARVALID,
    input  wire                            M_AXIMM_125_ARREADY,
    input  wire [M_AXIMM_125_DATA_WIDTH-1:0]   M_AXIMM_125_RDATA,
    input  wire [1:0]                      M_AXIMM_125_RRESP,
    input  wire                            M_AXIMM_125_RLAST,
    input  wire                            M_AXIMM_125_RVALID,
    output wire                            M_AXIMM_125_RREADY,
    //AXI-MM pass-through interface 126
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_126_AWADDR,
    input wire [7:0]                      AP_AXIMM_126_AWLEN,
    input wire [2:0]                      AP_AXIMM_126_AWSIZE,
    input wire [1:0]                      AP_AXIMM_126_AWBURST,
    input wire [1:0]                      AP_AXIMM_126_AWLOCK,
    input wire [3:0]                      AP_AXIMM_126_AWCACHE,
    input wire [2:0]                      AP_AXIMM_126_AWPROT,
    input wire [3:0]                      AP_AXIMM_126_AWREGION,
    input wire [3:0]                      AP_AXIMM_126_AWQOS,
    input wire                            AP_AXIMM_126_AWVALID,
    output  wire                            AP_AXIMM_126_AWREADY,
    input wire [M_AXIMM_126_DATA_WIDTH-1:0]   AP_AXIMM_126_WDATA,
    input wire [M_AXIMM_126_DATA_WIDTH/8-1:0] AP_AXIMM_126_WSTRB,
    input wire                            AP_AXIMM_126_WLAST,
    input wire                            AP_AXIMM_126_WVALID,
    output  wire                            AP_AXIMM_126_WREADY,
    output  wire [1:0]                      AP_AXIMM_126_BRESP,
    output  wire                            AP_AXIMM_126_BVALID,
    input wire                            AP_AXIMM_126_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_126_ARADDR,
    input wire [7:0]                      AP_AXIMM_126_ARLEN,
    input wire [2:0]                      AP_AXIMM_126_ARSIZE,
    input wire [1:0]                      AP_AXIMM_126_ARBURST,
    input wire [1:0]                      AP_AXIMM_126_ARLOCK,
    input wire [3:0]                      AP_AXIMM_126_ARCACHE,
    input wire [2:0]                      AP_AXIMM_126_ARPROT,
    input wire [3:0]                      AP_AXIMM_126_ARREGION,
    input wire [3:0]                      AP_AXIMM_126_ARQOS,
    input wire                            AP_AXIMM_126_ARVALID,
    output  wire                            AP_AXIMM_126_ARREADY,
    output  wire [M_AXIMM_126_DATA_WIDTH-1:0]   AP_AXIMM_126_RDATA,
    output  wire [1:0]                      AP_AXIMM_126_RRESP,
    output  wire                            AP_AXIMM_126_RLAST,
    output  wire                            AP_AXIMM_126_RVALID,
    input  wire                            AP_AXIMM_126_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_126_AWADDR,
    output wire [7:0]                      M_AXIMM_126_AWLEN,
    output wire [2:0]                      M_AXIMM_126_AWSIZE,
    output wire [1:0]                      M_AXIMM_126_AWBURST,
    output wire [1:0]                      M_AXIMM_126_AWLOCK,
    output wire [3:0]                      M_AXIMM_126_AWCACHE,
    output wire [2:0]                      M_AXIMM_126_AWPROT,
    output wire [3:0]                      M_AXIMM_126_AWREGION,
    output wire [3:0]                      M_AXIMM_126_AWQOS,
    output wire                            M_AXIMM_126_AWVALID,
    input  wire                            M_AXIMM_126_AWREADY,
    output wire [M_AXIMM_126_DATA_WIDTH-1:0]   M_AXIMM_126_WDATA,
    output wire [M_AXIMM_126_DATA_WIDTH/8-1:0] M_AXIMM_126_WSTRB,
    output wire                            M_AXIMM_126_WLAST,
    output wire                            M_AXIMM_126_WVALID,
    input  wire                            M_AXIMM_126_WREADY,
    input  wire [1:0]                      M_AXIMM_126_BRESP,
    input  wire                            M_AXIMM_126_BVALID,
    output wire                            M_AXIMM_126_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_126_ARADDR,
    output wire [7:0]                      M_AXIMM_126_ARLEN,
    output wire [2:0]                      M_AXIMM_126_ARSIZE,
    output wire [1:0]                      M_AXIMM_126_ARBURST,
    output wire [1:0]                      M_AXIMM_126_ARLOCK,
    output wire [3:0]                      M_AXIMM_126_ARCACHE,
    output wire [2:0]                      M_AXIMM_126_ARPROT,
    output wire [3:0]                      M_AXIMM_126_ARREGION,
    output wire [3:0]                      M_AXIMM_126_ARQOS,
    output wire                            M_AXIMM_126_ARVALID,
    input  wire                            M_AXIMM_126_ARREADY,
    input  wire [M_AXIMM_126_DATA_WIDTH-1:0]   M_AXIMM_126_RDATA,
    input  wire [1:0]                      M_AXIMM_126_RRESP,
    input  wire                            M_AXIMM_126_RLAST,
    input  wire                            M_AXIMM_126_RVALID,
    output wire                            M_AXIMM_126_RREADY,
    //AXI-MM pass-through interface 127
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_127_AWADDR,
    input wire [7:0]                      AP_AXIMM_127_AWLEN,
    input wire [2:0]                      AP_AXIMM_127_AWSIZE,
    input wire [1:0]                      AP_AXIMM_127_AWBURST,
    input wire [1:0]                      AP_AXIMM_127_AWLOCK,
    input wire [3:0]                      AP_AXIMM_127_AWCACHE,
    input wire [2:0]                      AP_AXIMM_127_AWPROT,
    input wire [3:0]                      AP_AXIMM_127_AWREGION,
    input wire [3:0]                      AP_AXIMM_127_AWQOS,
    input wire                            AP_AXIMM_127_AWVALID,
    output  wire                            AP_AXIMM_127_AWREADY,
    input wire [M_AXIMM_127_DATA_WIDTH-1:0]   AP_AXIMM_127_WDATA,
    input wire [M_AXIMM_127_DATA_WIDTH/8-1:0] AP_AXIMM_127_WSTRB,
    input wire                            AP_AXIMM_127_WLAST,
    input wire                            AP_AXIMM_127_WVALID,
    output  wire                            AP_AXIMM_127_WREADY,
    output  wire [1:0]                      AP_AXIMM_127_BRESP,
    output  wire                            AP_AXIMM_127_BVALID,
    input wire                            AP_AXIMM_127_BREADY,
    input wire [M_AXIMM_ADDR_WIDTH-1:0]   AP_AXIMM_127_ARADDR,
    input wire [7:0]                      AP_AXIMM_127_ARLEN,
    input wire [2:0]                      AP_AXIMM_127_ARSIZE,
    input wire [1:0]                      AP_AXIMM_127_ARBURST,
    input wire [1:0]                      AP_AXIMM_127_ARLOCK,
    input wire [3:0]                      AP_AXIMM_127_ARCACHE,
    input wire [2:0]                      AP_AXIMM_127_ARPROT,
    input wire [3:0]                      AP_AXIMM_127_ARREGION,
    input wire [3:0]                      AP_AXIMM_127_ARQOS,
    input wire                            AP_AXIMM_127_ARVALID,
    output  wire                            AP_AXIMM_127_ARREADY,
    output  wire [M_AXIMM_127_DATA_WIDTH-1:0]   AP_AXIMM_127_RDATA,
    output  wire [1:0]                      AP_AXIMM_127_RRESP,
    output  wire                            AP_AXIMM_127_RLAST,
    output  wire                            AP_AXIMM_127_RVALID,
    input  wire                            AP_AXIMM_127_RREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_127_AWADDR,
    output wire [7:0]                      M_AXIMM_127_AWLEN,
    output wire [2:0]                      M_AXIMM_127_AWSIZE,
    output wire [1:0]                      M_AXIMM_127_AWBURST,
    output wire [1:0]                      M_AXIMM_127_AWLOCK,
    output wire [3:0]                      M_AXIMM_127_AWCACHE,
    output wire [2:0]                      M_AXIMM_127_AWPROT,
    output wire [3:0]                      M_AXIMM_127_AWREGION,
    output wire [3:0]                      M_AXIMM_127_AWQOS,
    output wire                            M_AXIMM_127_AWVALID,
    input  wire                            M_AXIMM_127_AWREADY,
    output wire [M_AXIMM_127_DATA_WIDTH-1:0]   M_AXIMM_127_WDATA,
    output wire [M_AXIMM_127_DATA_WIDTH/8-1:0] M_AXIMM_127_WSTRB,
    output wire                            M_AXIMM_127_WLAST,
    output wire                            M_AXIMM_127_WVALID,
    input  wire                            M_AXIMM_127_WREADY,
    input  wire [1:0]                      M_AXIMM_127_BRESP,
    input  wire                            M_AXIMM_127_BVALID,
    output wire                            M_AXIMM_127_BREADY,
    output wire [M_AXIMM_ADDR_WIDTH-1:0]   M_AXIMM_127_ARADDR,
    output wire [7:0]                      M_AXIMM_127_ARLEN,
    output wire [2:0]                      M_AXIMM_127_ARSIZE,
    output wire [1:0]                      M_AXIMM_127_ARBURST,
    output wire [1:0]                      M_AXIMM_127_ARLOCK,
    output wire [3:0]                      M_AXIMM_127_ARCACHE,
    output wire [2:0]                      M_AXIMM_127_ARPROT,
    output wire [3:0]                      M_AXIMM_127_ARREGION,
    output wire [3:0]                      M_AXIMM_127_ARQOS,
    output wire                            M_AXIMM_127_ARVALID,
    input  wire                            M_AXIMM_127_ARREADY,
    input  wire [M_AXIMM_127_DATA_WIDTH-1:0]   M_AXIMM_127_RDATA,
    input  wire [1:0]                      M_AXIMM_127_RRESP,
    input  wire                            M_AXIMM_127_RLAST,
    input  wire                            M_AXIMM_127_RVALID,
    output wire                            M_AXIMM_127_RREADY
    );

    localparam C_MAX_BIT_WIDTH = 1024;
    localparam C_MAX_AXIMMs = 128;
    localparam [(C_MAX_AXIMMs*32)-1:0] M_AXIMM_BIT_ARRAY = {M_AXIMM_127_DATA_WIDTH,M_AXIMM_126_DATA_WIDTH,M_AXIMM_125_DATA_WIDTH,M_AXIMM_124_DATA_WIDTH,M_AXIMM_123_DATA_WIDTH,M_AXIMM_122_DATA_WIDTH,M_AXIMM_121_DATA_WIDTH,M_AXIMM_120_DATA_WIDTH,M_AXIMM_119_DATA_WIDTH,M_AXIMM_118_DATA_WIDTH,M_AXIMM_117_DATA_WIDTH,M_AXIMM_116_DATA_WIDTH,M_AXIMM_115_DATA_WIDTH,M_AXIMM_114_DATA_WIDTH,M_AXIMM_113_DATA_WIDTH,M_AXIMM_112_DATA_WIDTH,M_AXIMM_111_DATA_WIDTH,M_AXIMM_110_DATA_WIDTH,M_AXIMM_109_DATA_WIDTH,M_AXIMM_108_DATA_WIDTH,M_AXIMM_107_DATA_WIDTH,M_AXIMM_106_DATA_WIDTH,M_AXIMM_105_DATA_WIDTH,M_AXIMM_104_DATA_WIDTH,M_AXIMM_103_DATA_WIDTH,M_AXIMM_102_DATA_WIDTH,M_AXIMM_101_DATA_WIDTH,M_AXIMM_100_DATA_WIDTH,M_AXIMM_99_DATA_WIDTH,M_AXIMM_98_DATA_WIDTH,M_AXIMM_97_DATA_WIDTH,M_AXIMM_96_DATA_WIDTH,M_AXIMM_95_DATA_WIDTH,M_AXIMM_94_DATA_WIDTH,M_AXIMM_93_DATA_WIDTH,M_AXIMM_92_DATA_WIDTH,M_AXIMM_91_DATA_WIDTH,M_AXIMM_90_DATA_WIDTH,M_AXIMM_89_DATA_WIDTH,M_AXIMM_88_DATA_WIDTH,M_AXIMM_87_DATA_WIDTH,M_AXIMM_86_DATA_WIDTH,M_AXIMM_85_DATA_WIDTH,M_AXIMM_84_DATA_WIDTH,M_AXIMM_83_DATA_WIDTH,M_AXIMM_82_DATA_WIDTH,M_AXIMM_81_DATA_WIDTH,M_AXIMM_80_DATA_WIDTH,M_AXIMM_79_DATA_WIDTH,M_AXIMM_78_DATA_WIDTH,M_AXIMM_77_DATA_WIDTH,M_AXIMM_76_DATA_WIDTH,M_AXIMM_75_DATA_WIDTH,M_AXIMM_74_DATA_WIDTH,M_AXIMM_73_DATA_WIDTH,M_AXIMM_72_DATA_WIDTH,M_AXIMM_71_DATA_WIDTH,M_AXIMM_70_DATA_WIDTH,M_AXIMM_69_DATA_WIDTH,M_AXIMM_68_DATA_WIDTH,M_AXIMM_67_DATA_WIDTH,M_AXIMM_66_DATA_WIDTH,M_AXIMM_65_DATA_WIDTH,M_AXIMM_64_DATA_WIDTH,M_AXIMM_63_DATA_WIDTH,M_AXIMM_62_DATA_WIDTH,M_AXIMM_61_DATA_WIDTH,M_AXIMM_60_DATA_WIDTH,M_AXIMM_59_DATA_WIDTH,M_AXIMM_58_DATA_WIDTH,M_AXIMM_57_DATA_WIDTH,M_AXIMM_56_DATA_WIDTH,M_AXIMM_55_DATA_WIDTH,M_AXIMM_54_DATA_WIDTH,M_AXIMM_53_DATA_WIDTH,M_AXIMM_52_DATA_WIDTH,M_AXIMM_51_DATA_WIDTH,M_AXIMM_50_DATA_WIDTH,M_AXIMM_49_DATA_WIDTH,M_AXIMM_48_DATA_WIDTH,M_AXIMM_47_DATA_WIDTH,M_AXIMM_46_DATA_WIDTH,M_AXIMM_45_DATA_WIDTH,M_AXIMM_44_DATA_WIDTH,M_AXIMM_43_DATA_WIDTH,M_AXIMM_42_DATA_WIDTH,M_AXIMM_41_DATA_WIDTH,M_AXIMM_40_DATA_WIDTH,M_AXIMM_39_DATA_WIDTH,M_AXIMM_38_DATA_WIDTH,M_AXIMM_37_DATA_WIDTH,M_AXIMM_36_DATA_WIDTH,M_AXIMM_35_DATA_WIDTH,M_AXIMM_34_DATA_WIDTH,M_AXIMM_33_DATA_WIDTH,M_AXIMM_32_DATA_WIDTH,M_AXIMM_31_DATA_WIDTH,M_AXIMM_30_DATA_WIDTH,M_AXIMM_29_DATA_WIDTH,M_AXIMM_28_DATA_WIDTH,M_AXIMM_27_DATA_WIDTH,M_AXIMM_26_DATA_WIDTH,M_AXIMM_25_DATA_WIDTH,M_AXIMM_24_DATA_WIDTH,M_AXIMM_23_DATA_WIDTH,M_AXIMM_22_DATA_WIDTH,M_AXIMM_21_DATA_WIDTH,M_AXIMM_20_DATA_WIDTH,M_AXIMM_19_DATA_WIDTH,M_AXIMM_18_DATA_WIDTH,M_AXIMM_17_DATA_WIDTH,M_AXIMM_16_DATA_WIDTH,M_AXIMM_15_DATA_WIDTH,M_AXIMM_14_DATA_WIDTH,M_AXIMM_13_DATA_WIDTH,M_AXIMM_12_DATA_WIDTH,M_AXIMM_11_DATA_WIDTH,M_AXIMM_10_DATA_WIDTH,M_AXIMM_9_DATA_WIDTH,M_AXIMM_8_DATA_WIDTH,M_AXIMM_7_DATA_WIDTH,M_AXIMM_6_DATA_WIDTH,M_AXIMM_5_DATA_WIDTH,M_AXIMM_4_DATA_WIDTH,M_AXIMM_3_DATA_WIDTH,M_AXIMM_2_DATA_WIDTH,M_AXIMM_1_DATA_WIDTH,M_AXIMM_0_DATA_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_ARUSER_ARRAY = {M_AXIMM_127_ARUSER_WIDTH,M_AXIMM_126_ARUSER_WIDTH,M_AXIMM_125_ARUSER_WIDTH,M_AXIMM_124_ARUSER_WIDTH,M_AXIMM_123_ARUSER_WIDTH,M_AXIMM_122_ARUSER_WIDTH,M_AXIMM_121_ARUSER_WIDTH,M_AXIMM_120_ARUSER_WIDTH,M_AXIMM_119_ARUSER_WIDTH,M_AXIMM_118_ARUSER_WIDTH,M_AXIMM_117_ARUSER_WIDTH,M_AXIMM_116_ARUSER_WIDTH,M_AXIMM_115_ARUSER_WIDTH,M_AXIMM_114_ARUSER_WIDTH,M_AXIMM_113_ARUSER_WIDTH,M_AXIMM_112_ARUSER_WIDTH,M_AXIMM_111_ARUSER_WIDTH,M_AXIMM_110_ARUSER_WIDTH,M_AXIMM_109_ARUSER_WIDTH,M_AXIMM_108_ARUSER_WIDTH,M_AXIMM_107_ARUSER_WIDTH,M_AXIMM_106_ARUSER_WIDTH,M_AXIMM_105_ARUSER_WIDTH,M_AXIMM_104_ARUSER_WIDTH,M_AXIMM_103_ARUSER_WIDTH,M_AXIMM_102_ARUSER_WIDTH,M_AXIMM_101_ARUSER_WIDTH,M_AXIMM_100_ARUSER_WIDTH,M_AXIMM_99_ARUSER_WIDTH,M_AXIMM_98_ARUSER_WIDTH,M_AXIMM_97_ARUSER_WIDTH,M_AXIMM_96_ARUSER_WIDTH,M_AXIMM_95_ARUSER_WIDTH,M_AXIMM_94_ARUSER_WIDTH,M_AXIMM_93_ARUSER_WIDTH,M_AXIMM_92_ARUSER_WIDTH,M_AXIMM_91_ARUSER_WIDTH,M_AXIMM_90_ARUSER_WIDTH,M_AXIMM_89_ARUSER_WIDTH,M_AXIMM_88_ARUSER_WIDTH,M_AXIMM_87_ARUSER_WIDTH,M_AXIMM_86_ARUSER_WIDTH,M_AXIMM_85_ARUSER_WIDTH,M_AXIMM_84_ARUSER_WIDTH,M_AXIMM_83_ARUSER_WIDTH,M_AXIMM_82_ARUSER_WIDTH,M_AXIMM_81_ARUSER_WIDTH,M_AXIMM_80_ARUSER_WIDTH,M_AXIMM_79_ARUSER_WIDTH,M_AXIMM_78_ARUSER_WIDTH,M_AXIMM_77_ARUSER_WIDTH,M_AXIMM_76_ARUSER_WIDTH,M_AXIMM_75_ARUSER_WIDTH,M_AXIMM_74_ARUSER_WIDTH,M_AXIMM_73_ARUSER_WIDTH,M_AXIMM_72_ARUSER_WIDTH,M_AXIMM_71_ARUSER_WIDTH,M_AXIMM_70_ARUSER_WIDTH,M_AXIMM_69_ARUSER_WIDTH,M_AXIMM_68_ARUSER_WIDTH,M_AXIMM_67_ARUSER_WIDTH,M_AXIMM_66_ARUSER_WIDTH,M_AXIMM_65_ARUSER_WIDTH,M_AXIMM_64_ARUSER_WIDTH,M_AXIMM_63_ARUSER_WIDTH,M_AXIMM_62_ARUSER_WIDTH,M_AXIMM_61_ARUSER_WIDTH,M_AXIMM_60_ARUSER_WIDTH,M_AXIMM_59_ARUSER_WIDTH,M_AXIMM_58_ARUSER_WIDTH,M_AXIMM_57_ARUSER_WIDTH,M_AXIMM_56_ARUSER_WIDTH,M_AXIMM_55_ARUSER_WIDTH,M_AXIMM_54_ARUSER_WIDTH,M_AXIMM_53_ARUSER_WIDTH,M_AXIMM_52_ARUSER_WIDTH,M_AXIMM_51_ARUSER_WIDTH,M_AXIMM_50_ARUSER_WIDTH,M_AXIMM_49_ARUSER_WIDTH,M_AXIMM_48_ARUSER_WIDTH,M_AXIMM_47_ARUSER_WIDTH,M_AXIMM_46_ARUSER_WIDTH,M_AXIMM_45_ARUSER_WIDTH,M_AXIMM_44_ARUSER_WIDTH,M_AXIMM_43_ARUSER_WIDTH,M_AXIMM_42_ARUSER_WIDTH,M_AXIMM_41_ARUSER_WIDTH,M_AXIMM_40_ARUSER_WIDTH,M_AXIMM_39_ARUSER_WIDTH,M_AXIMM_38_ARUSER_WIDTH,M_AXIMM_37_ARUSER_WIDTH,M_AXIMM_36_ARUSER_WIDTH,M_AXIMM_35_ARUSER_WIDTH,M_AXIMM_34_ARUSER_WIDTH,M_AXIMM_33_ARUSER_WIDTH,M_AXIMM_32_ARUSER_WIDTH,M_AXIMM_31_ARUSER_WIDTH,M_AXIMM_30_ARUSER_WIDTH,M_AXIMM_29_ARUSER_WIDTH,M_AXIMM_28_ARUSER_WIDTH,M_AXIMM_27_ARUSER_WIDTH,M_AXIMM_26_ARUSER_WIDTH,M_AXIMM_25_ARUSER_WIDTH,M_AXIMM_24_ARUSER_WIDTH,M_AXIMM_23_ARUSER_WIDTH,M_AXIMM_22_ARUSER_WIDTH,M_AXIMM_21_ARUSER_WIDTH,M_AXIMM_20_ARUSER_WIDTH,M_AXIMM_19_ARUSER_WIDTH,M_AXIMM_18_ARUSER_WIDTH,M_AXIMM_17_ARUSER_WIDTH,M_AXIMM_16_ARUSER_WIDTH,M_AXIMM_15_ARUSER_WIDTH,M_AXIMM_14_ARUSER_WIDTH,M_AXIMM_13_ARUSER_WIDTH,M_AXIMM_12_ARUSER_WIDTH,M_AXIMM_11_ARUSER_WIDTH,M_AXIMM_10_ARUSER_WIDTH,M_AXIMM_9_ARUSER_WIDTH,M_AXIMM_8_ARUSER_WIDTH,M_AXIMM_7_ARUSER_WIDTH,M_AXIMM_6_ARUSER_WIDTH,M_AXIMM_5_ARUSER_WIDTH,M_AXIMM_4_ARUSER_WIDTH,M_AXIMM_3_ARUSER_WIDTH,M_AXIMM_2_ARUSER_WIDTH,M_AXIMM_1_ARUSER_WIDTH,M_AXIMM_0_ARUSER_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_AWUSER_ARRAY = {M_AXIMM_127_AWUSER_WIDTH,M_AXIMM_126_AWUSER_WIDTH,M_AXIMM_125_AWUSER_WIDTH,M_AXIMM_124_AWUSER_WIDTH,M_AXIMM_123_AWUSER_WIDTH,M_AXIMM_122_AWUSER_WIDTH,M_AXIMM_121_AWUSER_WIDTH,M_AXIMM_120_AWUSER_WIDTH,M_AXIMM_119_AWUSER_WIDTH,M_AXIMM_118_AWUSER_WIDTH,M_AXIMM_117_AWUSER_WIDTH,M_AXIMM_116_AWUSER_WIDTH,M_AXIMM_115_AWUSER_WIDTH,M_AXIMM_114_AWUSER_WIDTH,M_AXIMM_113_AWUSER_WIDTH,M_AXIMM_112_AWUSER_WIDTH,M_AXIMM_111_AWUSER_WIDTH,M_AXIMM_110_AWUSER_WIDTH,M_AXIMM_109_AWUSER_WIDTH,M_AXIMM_108_AWUSER_WIDTH,M_AXIMM_107_AWUSER_WIDTH,M_AXIMM_106_AWUSER_WIDTH,M_AXIMM_105_AWUSER_WIDTH,M_AXIMM_104_AWUSER_WIDTH,M_AXIMM_103_AWUSER_WIDTH,M_AXIMM_102_AWUSER_WIDTH,M_AXIMM_101_AWUSER_WIDTH,M_AXIMM_100_AWUSER_WIDTH,M_AXIMM_99_AWUSER_WIDTH,M_AXIMM_98_AWUSER_WIDTH,M_AXIMM_97_AWUSER_WIDTH,M_AXIMM_96_AWUSER_WIDTH,M_AXIMM_95_AWUSER_WIDTH,M_AXIMM_94_AWUSER_WIDTH,M_AXIMM_93_AWUSER_WIDTH,M_AXIMM_92_AWUSER_WIDTH,M_AXIMM_91_AWUSER_WIDTH,M_AXIMM_90_AWUSER_WIDTH,M_AXIMM_89_AWUSER_WIDTH,M_AXIMM_88_AWUSER_WIDTH,M_AXIMM_87_AWUSER_WIDTH,M_AXIMM_86_AWUSER_WIDTH,M_AXIMM_85_AWUSER_WIDTH,M_AXIMM_84_AWUSER_WIDTH,M_AXIMM_83_AWUSER_WIDTH,M_AXIMM_82_AWUSER_WIDTH,M_AXIMM_81_AWUSER_WIDTH,M_AXIMM_80_AWUSER_WIDTH,M_AXIMM_79_AWUSER_WIDTH,M_AXIMM_78_AWUSER_WIDTH,M_AXIMM_77_AWUSER_WIDTH,M_AXIMM_76_AWUSER_WIDTH,M_AXIMM_75_AWUSER_WIDTH,M_AXIMM_74_AWUSER_WIDTH,M_AXIMM_73_AWUSER_WIDTH,M_AXIMM_72_AWUSER_WIDTH,M_AXIMM_71_AWUSER_WIDTH,M_AXIMM_70_AWUSER_WIDTH,M_AXIMM_69_AWUSER_WIDTH,M_AXIMM_68_AWUSER_WIDTH,M_AXIMM_67_AWUSER_WIDTH,M_AXIMM_66_AWUSER_WIDTH,M_AXIMM_65_AWUSER_WIDTH,M_AXIMM_64_AWUSER_WIDTH,M_AXIMM_63_AWUSER_WIDTH,M_AXIMM_62_AWUSER_WIDTH,M_AXIMM_61_AWUSER_WIDTH,M_AXIMM_60_AWUSER_WIDTH,M_AXIMM_59_AWUSER_WIDTH,M_AXIMM_58_AWUSER_WIDTH,M_AXIMM_57_AWUSER_WIDTH,M_AXIMM_56_AWUSER_WIDTH,M_AXIMM_55_AWUSER_WIDTH,M_AXIMM_54_AWUSER_WIDTH,M_AXIMM_53_AWUSER_WIDTH,M_AXIMM_52_AWUSER_WIDTH,M_AXIMM_51_AWUSER_WIDTH,M_AXIMM_50_AWUSER_WIDTH,M_AXIMM_49_AWUSER_WIDTH,M_AXIMM_48_AWUSER_WIDTH,M_AXIMM_47_AWUSER_WIDTH,M_AXIMM_46_AWUSER_WIDTH,M_AXIMM_45_AWUSER_WIDTH,M_AXIMM_44_AWUSER_WIDTH,M_AXIMM_43_AWUSER_WIDTH,M_AXIMM_42_AWUSER_WIDTH,M_AXIMM_41_AWUSER_WIDTH,M_AXIMM_40_AWUSER_WIDTH,M_AXIMM_39_AWUSER_WIDTH,M_AXIMM_38_AWUSER_WIDTH,M_AXIMM_37_AWUSER_WIDTH,M_AXIMM_36_AWUSER_WIDTH,M_AXIMM_35_AWUSER_WIDTH,M_AXIMM_34_AWUSER_WIDTH,M_AXIMM_33_AWUSER_WIDTH,M_AXIMM_32_AWUSER_WIDTH,M_AXIMM_31_AWUSER_WIDTH,M_AXIMM_30_AWUSER_WIDTH,M_AXIMM_29_AWUSER_WIDTH,M_AXIMM_28_AWUSER_WIDTH,M_AXIMM_27_AWUSER_WIDTH,M_AXIMM_26_AWUSER_WIDTH,M_AXIMM_25_AWUSER_WIDTH,M_AXIMM_24_AWUSER_WIDTH,M_AXIMM_23_AWUSER_WIDTH,M_AXIMM_22_AWUSER_WIDTH,M_AXIMM_21_AWUSER_WIDTH,M_AXIMM_20_AWUSER_WIDTH,M_AXIMM_19_AWUSER_WIDTH,M_AXIMM_18_AWUSER_WIDTH,M_AXIMM_17_AWUSER_WIDTH,M_AXIMM_16_AWUSER_WIDTH,M_AXIMM_15_AWUSER_WIDTH,M_AXIMM_14_AWUSER_WIDTH,M_AXIMM_13_AWUSER_WIDTH,M_AXIMM_12_AWUSER_WIDTH,M_AXIMM_11_AWUSER_WIDTH,M_AXIMM_10_AWUSER_WIDTH,M_AXIMM_9_AWUSER_WIDTH,M_AXIMM_8_AWUSER_WIDTH,M_AXIMM_7_AWUSER_WIDTH,M_AXIMM_6_AWUSER_WIDTH,M_AXIMM_5_AWUSER_WIDTH,M_AXIMM_4_AWUSER_WIDTH,M_AXIMM_3_AWUSER_WIDTH,M_AXIMM_2_AWUSER_WIDTH,M_AXIMM_1_AWUSER_WIDTH,M_AXIMM_0_AWUSER_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_BUSER_ARRAY = {M_AXIMM_127_BUSER_WIDTH,M_AXIMM_126_BUSER_WIDTH,M_AXIMM_125_BUSER_WIDTH,M_AXIMM_124_BUSER_WIDTH,M_AXIMM_123_BUSER_WIDTH,M_AXIMM_122_BUSER_WIDTH,M_AXIMM_121_BUSER_WIDTH,M_AXIMM_120_BUSER_WIDTH,M_AXIMM_119_BUSER_WIDTH,M_AXIMM_118_BUSER_WIDTH,M_AXIMM_117_BUSER_WIDTH,M_AXIMM_116_BUSER_WIDTH,M_AXIMM_115_BUSER_WIDTH,M_AXIMM_114_BUSER_WIDTH,M_AXIMM_113_BUSER_WIDTH,M_AXIMM_112_BUSER_WIDTH,M_AXIMM_111_BUSER_WIDTH,M_AXIMM_110_BUSER_WIDTH,M_AXIMM_109_BUSER_WIDTH,M_AXIMM_108_BUSER_WIDTH,M_AXIMM_107_BUSER_WIDTH,M_AXIMM_106_BUSER_WIDTH,M_AXIMM_105_BUSER_WIDTH,M_AXIMM_104_BUSER_WIDTH,M_AXIMM_103_BUSER_WIDTH,M_AXIMM_102_BUSER_WIDTH,M_AXIMM_101_BUSER_WIDTH,M_AXIMM_100_BUSER_WIDTH,M_AXIMM_99_BUSER_WIDTH,M_AXIMM_98_BUSER_WIDTH,M_AXIMM_97_BUSER_WIDTH,M_AXIMM_96_BUSER_WIDTH,M_AXIMM_95_BUSER_WIDTH,M_AXIMM_94_BUSER_WIDTH,M_AXIMM_93_BUSER_WIDTH,M_AXIMM_92_BUSER_WIDTH,M_AXIMM_91_BUSER_WIDTH,M_AXIMM_90_BUSER_WIDTH,M_AXIMM_89_BUSER_WIDTH,M_AXIMM_88_BUSER_WIDTH,M_AXIMM_87_BUSER_WIDTH,M_AXIMM_86_BUSER_WIDTH,M_AXIMM_85_BUSER_WIDTH,M_AXIMM_84_BUSER_WIDTH,M_AXIMM_83_BUSER_WIDTH,M_AXIMM_82_BUSER_WIDTH,M_AXIMM_81_BUSER_WIDTH,M_AXIMM_80_BUSER_WIDTH,M_AXIMM_79_BUSER_WIDTH,M_AXIMM_78_BUSER_WIDTH,M_AXIMM_77_BUSER_WIDTH,M_AXIMM_76_BUSER_WIDTH,M_AXIMM_75_BUSER_WIDTH,M_AXIMM_74_BUSER_WIDTH,M_AXIMM_73_BUSER_WIDTH,M_AXIMM_72_BUSER_WIDTH,M_AXIMM_71_BUSER_WIDTH,M_AXIMM_70_BUSER_WIDTH,M_AXIMM_69_BUSER_WIDTH,M_AXIMM_68_BUSER_WIDTH,M_AXIMM_67_BUSER_WIDTH,M_AXIMM_66_BUSER_WIDTH,M_AXIMM_65_BUSER_WIDTH,M_AXIMM_64_BUSER_WIDTH,M_AXIMM_63_BUSER_WIDTH,M_AXIMM_62_BUSER_WIDTH,M_AXIMM_61_BUSER_WIDTH,M_AXIMM_60_BUSER_WIDTH,M_AXIMM_59_BUSER_WIDTH,M_AXIMM_58_BUSER_WIDTH,M_AXIMM_57_BUSER_WIDTH,M_AXIMM_56_BUSER_WIDTH,M_AXIMM_55_BUSER_WIDTH,M_AXIMM_54_BUSER_WIDTH,M_AXIMM_53_BUSER_WIDTH,M_AXIMM_52_BUSER_WIDTH,M_AXIMM_51_BUSER_WIDTH,M_AXIMM_50_BUSER_WIDTH,M_AXIMM_49_BUSER_WIDTH,M_AXIMM_48_BUSER_WIDTH,M_AXIMM_47_BUSER_WIDTH,M_AXIMM_46_BUSER_WIDTH,M_AXIMM_45_BUSER_WIDTH,M_AXIMM_44_BUSER_WIDTH,M_AXIMM_43_BUSER_WIDTH,M_AXIMM_42_BUSER_WIDTH,M_AXIMM_41_BUSER_WIDTH,M_AXIMM_40_BUSER_WIDTH,M_AXIMM_39_BUSER_WIDTH,M_AXIMM_38_BUSER_WIDTH,M_AXIMM_37_BUSER_WIDTH,M_AXIMM_36_BUSER_WIDTH,M_AXIMM_35_BUSER_WIDTH,M_AXIMM_34_BUSER_WIDTH,M_AXIMM_33_BUSER_WIDTH,M_AXIMM_32_BUSER_WIDTH,M_AXIMM_31_BUSER_WIDTH,M_AXIMM_30_BUSER_WIDTH,M_AXIMM_29_BUSER_WIDTH,M_AXIMM_28_BUSER_WIDTH,M_AXIMM_27_BUSER_WIDTH,M_AXIMM_26_BUSER_WIDTH,M_AXIMM_25_BUSER_WIDTH,M_AXIMM_24_BUSER_WIDTH,M_AXIMM_23_BUSER_WIDTH,M_AXIMM_22_BUSER_WIDTH,M_AXIMM_21_BUSER_WIDTH,M_AXIMM_20_BUSER_WIDTH,M_AXIMM_19_BUSER_WIDTH,M_AXIMM_18_BUSER_WIDTH,M_AXIMM_17_BUSER_WIDTH,M_AXIMM_16_BUSER_WIDTH,M_AXIMM_15_BUSER_WIDTH,M_AXIMM_14_BUSER_WIDTH,M_AXIMM_13_BUSER_WIDTH,M_AXIMM_12_BUSER_WIDTH,M_AXIMM_11_BUSER_WIDTH,M_AXIMM_10_BUSER_WIDTH,M_AXIMM_9_BUSER_WIDTH,M_AXIMM_8_BUSER_WIDTH,M_AXIMM_7_BUSER_WIDTH,M_AXIMM_6_BUSER_WIDTH,M_AXIMM_5_BUSER_WIDTH,M_AXIMM_4_BUSER_WIDTH,M_AXIMM_3_BUSER_WIDTH,M_AXIMM_2_BUSER_WIDTH,M_AXIMM_1_BUSER_WIDTH,M_AXIMM_0_BUSER_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_RUSER_ARRAY = {M_AXIMM_127_RUSER_WIDTH,M_AXIMM_126_RUSER_WIDTH,M_AXIMM_125_RUSER_WIDTH,M_AXIMM_124_RUSER_WIDTH,M_AXIMM_123_RUSER_WIDTH,M_AXIMM_122_RUSER_WIDTH,M_AXIMM_121_RUSER_WIDTH,M_AXIMM_120_RUSER_WIDTH,M_AXIMM_119_RUSER_WIDTH,M_AXIMM_118_RUSER_WIDTH,M_AXIMM_117_RUSER_WIDTH,M_AXIMM_116_RUSER_WIDTH,M_AXIMM_115_RUSER_WIDTH,M_AXIMM_114_RUSER_WIDTH,M_AXIMM_113_RUSER_WIDTH,M_AXIMM_112_RUSER_WIDTH,M_AXIMM_111_RUSER_WIDTH,M_AXIMM_110_RUSER_WIDTH,M_AXIMM_109_RUSER_WIDTH,M_AXIMM_108_RUSER_WIDTH,M_AXIMM_107_RUSER_WIDTH,M_AXIMM_106_RUSER_WIDTH,M_AXIMM_105_RUSER_WIDTH,M_AXIMM_104_RUSER_WIDTH,M_AXIMM_103_RUSER_WIDTH,M_AXIMM_102_RUSER_WIDTH,M_AXIMM_101_RUSER_WIDTH,M_AXIMM_100_RUSER_WIDTH,M_AXIMM_99_RUSER_WIDTH,M_AXIMM_98_RUSER_WIDTH,M_AXIMM_97_RUSER_WIDTH,M_AXIMM_96_RUSER_WIDTH,M_AXIMM_95_RUSER_WIDTH,M_AXIMM_94_RUSER_WIDTH,M_AXIMM_93_RUSER_WIDTH,M_AXIMM_92_RUSER_WIDTH,M_AXIMM_91_RUSER_WIDTH,M_AXIMM_90_RUSER_WIDTH,M_AXIMM_89_RUSER_WIDTH,M_AXIMM_88_RUSER_WIDTH,M_AXIMM_87_RUSER_WIDTH,M_AXIMM_86_RUSER_WIDTH,M_AXIMM_85_RUSER_WIDTH,M_AXIMM_84_RUSER_WIDTH,M_AXIMM_83_RUSER_WIDTH,M_AXIMM_82_RUSER_WIDTH,M_AXIMM_81_RUSER_WIDTH,M_AXIMM_80_RUSER_WIDTH,M_AXIMM_79_RUSER_WIDTH,M_AXIMM_78_RUSER_WIDTH,M_AXIMM_77_RUSER_WIDTH,M_AXIMM_76_RUSER_WIDTH,M_AXIMM_75_RUSER_WIDTH,M_AXIMM_74_RUSER_WIDTH,M_AXIMM_73_RUSER_WIDTH,M_AXIMM_72_RUSER_WIDTH,M_AXIMM_71_RUSER_WIDTH,M_AXIMM_70_RUSER_WIDTH,M_AXIMM_69_RUSER_WIDTH,M_AXIMM_68_RUSER_WIDTH,M_AXIMM_67_RUSER_WIDTH,M_AXIMM_66_RUSER_WIDTH,M_AXIMM_65_RUSER_WIDTH,M_AXIMM_64_RUSER_WIDTH,M_AXIMM_63_RUSER_WIDTH,M_AXIMM_62_RUSER_WIDTH,M_AXIMM_61_RUSER_WIDTH,M_AXIMM_60_RUSER_WIDTH,M_AXIMM_59_RUSER_WIDTH,M_AXIMM_58_RUSER_WIDTH,M_AXIMM_57_RUSER_WIDTH,M_AXIMM_56_RUSER_WIDTH,M_AXIMM_55_RUSER_WIDTH,M_AXIMM_54_RUSER_WIDTH,M_AXIMM_53_RUSER_WIDTH,M_AXIMM_52_RUSER_WIDTH,M_AXIMM_51_RUSER_WIDTH,M_AXIMM_50_RUSER_WIDTH,M_AXIMM_49_RUSER_WIDTH,M_AXIMM_48_RUSER_WIDTH,M_AXIMM_47_RUSER_WIDTH,M_AXIMM_46_RUSER_WIDTH,M_AXIMM_45_RUSER_WIDTH,M_AXIMM_44_RUSER_WIDTH,M_AXIMM_43_RUSER_WIDTH,M_AXIMM_42_RUSER_WIDTH,M_AXIMM_41_RUSER_WIDTH,M_AXIMM_40_RUSER_WIDTH,M_AXIMM_39_RUSER_WIDTH,M_AXIMM_38_RUSER_WIDTH,M_AXIMM_37_RUSER_WIDTH,M_AXIMM_36_RUSER_WIDTH,M_AXIMM_35_RUSER_WIDTH,M_AXIMM_34_RUSER_WIDTH,M_AXIMM_33_RUSER_WIDTH,M_AXIMM_32_RUSER_WIDTH,M_AXIMM_31_RUSER_WIDTH,M_AXIMM_30_RUSER_WIDTH,M_AXIMM_29_RUSER_WIDTH,M_AXIMM_28_RUSER_WIDTH,M_AXIMM_27_RUSER_WIDTH,M_AXIMM_26_RUSER_WIDTH,M_AXIMM_25_RUSER_WIDTH,M_AXIMM_24_RUSER_WIDTH,M_AXIMM_23_RUSER_WIDTH,M_AXIMM_22_RUSER_WIDTH,M_AXIMM_21_RUSER_WIDTH,M_AXIMM_20_RUSER_WIDTH,M_AXIMM_19_RUSER_WIDTH,M_AXIMM_18_RUSER_WIDTH,M_AXIMM_17_RUSER_WIDTH,M_AXIMM_16_RUSER_WIDTH,M_AXIMM_15_RUSER_WIDTH,M_AXIMM_14_RUSER_WIDTH,M_AXIMM_13_RUSER_WIDTH,M_AXIMM_12_RUSER_WIDTH,M_AXIMM_11_RUSER_WIDTH,M_AXIMM_10_RUSER_WIDTH,M_AXIMM_9_RUSER_WIDTH,M_AXIMM_8_RUSER_WIDTH,M_AXIMM_7_RUSER_WIDTH,M_AXIMM_6_RUSER_WIDTH,M_AXIMM_5_RUSER_WIDTH,M_AXIMM_4_RUSER_WIDTH,M_AXIMM_3_RUSER_WIDTH,M_AXIMM_2_RUSER_WIDTH,M_AXIMM_1_RUSER_WIDTH,M_AXIMM_0_RUSER_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_WUSER_ARRAY = {M_AXIMM_127_WUSER_WIDTH,M_AXIMM_126_WUSER_WIDTH,M_AXIMM_125_WUSER_WIDTH,M_AXIMM_124_WUSER_WIDTH,M_AXIMM_123_WUSER_WIDTH,M_AXIMM_122_WUSER_WIDTH,M_AXIMM_121_WUSER_WIDTH,M_AXIMM_120_WUSER_WIDTH,M_AXIMM_119_WUSER_WIDTH,M_AXIMM_118_WUSER_WIDTH,M_AXIMM_117_WUSER_WIDTH,M_AXIMM_116_WUSER_WIDTH,M_AXIMM_115_WUSER_WIDTH,M_AXIMM_114_WUSER_WIDTH,M_AXIMM_113_WUSER_WIDTH,M_AXIMM_112_WUSER_WIDTH,M_AXIMM_111_WUSER_WIDTH,M_AXIMM_110_WUSER_WIDTH,M_AXIMM_109_WUSER_WIDTH,M_AXIMM_108_WUSER_WIDTH,M_AXIMM_107_WUSER_WIDTH,M_AXIMM_106_WUSER_WIDTH,M_AXIMM_105_WUSER_WIDTH,M_AXIMM_104_WUSER_WIDTH,M_AXIMM_103_WUSER_WIDTH,M_AXIMM_102_WUSER_WIDTH,M_AXIMM_101_WUSER_WIDTH,M_AXIMM_100_WUSER_WIDTH,M_AXIMM_99_WUSER_WIDTH,M_AXIMM_98_WUSER_WIDTH,M_AXIMM_97_WUSER_WIDTH,M_AXIMM_96_WUSER_WIDTH,M_AXIMM_95_WUSER_WIDTH,M_AXIMM_94_WUSER_WIDTH,M_AXIMM_93_WUSER_WIDTH,M_AXIMM_92_WUSER_WIDTH,M_AXIMM_91_WUSER_WIDTH,M_AXIMM_90_WUSER_WIDTH,M_AXIMM_89_WUSER_WIDTH,M_AXIMM_88_WUSER_WIDTH,M_AXIMM_87_WUSER_WIDTH,M_AXIMM_86_WUSER_WIDTH,M_AXIMM_85_WUSER_WIDTH,M_AXIMM_84_WUSER_WIDTH,M_AXIMM_83_WUSER_WIDTH,M_AXIMM_82_WUSER_WIDTH,M_AXIMM_81_WUSER_WIDTH,M_AXIMM_80_WUSER_WIDTH,M_AXIMM_79_WUSER_WIDTH,M_AXIMM_78_WUSER_WIDTH,M_AXIMM_77_WUSER_WIDTH,M_AXIMM_76_WUSER_WIDTH,M_AXIMM_75_WUSER_WIDTH,M_AXIMM_74_WUSER_WIDTH,M_AXIMM_73_WUSER_WIDTH,M_AXIMM_72_WUSER_WIDTH,M_AXIMM_71_WUSER_WIDTH,M_AXIMM_70_WUSER_WIDTH,M_AXIMM_69_WUSER_WIDTH,M_AXIMM_68_WUSER_WIDTH,M_AXIMM_67_WUSER_WIDTH,M_AXIMM_66_WUSER_WIDTH,M_AXIMM_65_WUSER_WIDTH,M_AXIMM_64_WUSER_WIDTH,M_AXIMM_63_WUSER_WIDTH,M_AXIMM_62_WUSER_WIDTH,M_AXIMM_61_WUSER_WIDTH,M_AXIMM_60_WUSER_WIDTH,M_AXIMM_59_WUSER_WIDTH,M_AXIMM_58_WUSER_WIDTH,M_AXIMM_57_WUSER_WIDTH,M_AXIMM_56_WUSER_WIDTH,M_AXIMM_55_WUSER_WIDTH,M_AXIMM_54_WUSER_WIDTH,M_AXIMM_53_WUSER_WIDTH,M_AXIMM_52_WUSER_WIDTH,M_AXIMM_51_WUSER_WIDTH,M_AXIMM_50_WUSER_WIDTH,M_AXIMM_49_WUSER_WIDTH,M_AXIMM_48_WUSER_WIDTH,M_AXIMM_47_WUSER_WIDTH,M_AXIMM_46_WUSER_WIDTH,M_AXIMM_45_WUSER_WIDTH,M_AXIMM_44_WUSER_WIDTH,M_AXIMM_43_WUSER_WIDTH,M_AXIMM_42_WUSER_WIDTH,M_AXIMM_41_WUSER_WIDTH,M_AXIMM_40_WUSER_WIDTH,M_AXIMM_39_WUSER_WIDTH,M_AXIMM_38_WUSER_WIDTH,M_AXIMM_37_WUSER_WIDTH,M_AXIMM_36_WUSER_WIDTH,M_AXIMM_35_WUSER_WIDTH,M_AXIMM_34_WUSER_WIDTH,M_AXIMM_33_WUSER_WIDTH,M_AXIMM_32_WUSER_WIDTH,M_AXIMM_31_WUSER_WIDTH,M_AXIMM_30_WUSER_WIDTH,M_AXIMM_29_WUSER_WIDTH,M_AXIMM_28_WUSER_WIDTH,M_AXIMM_27_WUSER_WIDTH,M_AXIMM_26_WUSER_WIDTH,M_AXIMM_25_WUSER_WIDTH,M_AXIMM_24_WUSER_WIDTH,M_AXIMM_23_WUSER_WIDTH,M_AXIMM_22_WUSER_WIDTH,M_AXIMM_21_WUSER_WIDTH,M_AXIMM_20_WUSER_WIDTH,M_AXIMM_19_WUSER_WIDTH,M_AXIMM_18_WUSER_WIDTH,M_AXIMM_17_WUSER_WIDTH,M_AXIMM_16_WUSER_WIDTH,M_AXIMM_15_WUSER_WIDTH,M_AXIMM_14_WUSER_WIDTH,M_AXIMM_13_WUSER_WIDTH,M_AXIMM_12_WUSER_WIDTH,M_AXIMM_11_WUSER_WIDTH,M_AXIMM_10_WUSER_WIDTH,M_AXIMM_9_WUSER_WIDTH,M_AXIMM_8_WUSER_WIDTH,M_AXIMM_7_WUSER_WIDTH,M_AXIMM_6_WUSER_WIDTH,M_AXIMM_5_WUSER_WIDTH,M_AXIMM_4_WUSER_WIDTH,M_AXIMM_3_WUSER_WIDTH,M_AXIMM_2_WUSER_WIDTH,M_AXIMM_1_WUSER_WIDTH,M_AXIMM_0_WUSER_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_ARID_ARRAY = {M_AXIMM_127_ARID_WIDTH,M_AXIMM_126_ARID_WIDTH,M_AXIMM_125_ARID_WIDTH,M_AXIMM_124_ARID_WIDTH,M_AXIMM_123_ARID_WIDTH,M_AXIMM_122_ARID_WIDTH,M_AXIMM_121_ARID_WIDTH,M_AXIMM_120_ARID_WIDTH,M_AXIMM_119_ARID_WIDTH,M_AXIMM_118_ARID_WIDTH,M_AXIMM_117_ARID_WIDTH,M_AXIMM_116_ARID_WIDTH,M_AXIMM_115_ARID_WIDTH,M_AXIMM_114_ARID_WIDTH,M_AXIMM_113_ARID_WIDTH,M_AXIMM_112_ARID_WIDTH,M_AXIMM_111_ARID_WIDTH,M_AXIMM_110_ARID_WIDTH,M_AXIMM_109_ARID_WIDTH,M_AXIMM_108_ARID_WIDTH,M_AXIMM_107_ARID_WIDTH,M_AXIMM_106_ARID_WIDTH,M_AXIMM_105_ARID_WIDTH,M_AXIMM_104_ARID_WIDTH,M_AXIMM_103_ARID_WIDTH,M_AXIMM_102_ARID_WIDTH,M_AXIMM_101_ARID_WIDTH,M_AXIMM_100_ARID_WIDTH,M_AXIMM_99_ARID_WIDTH,M_AXIMM_98_ARID_WIDTH,M_AXIMM_97_ARID_WIDTH,M_AXIMM_96_ARID_WIDTH,M_AXIMM_95_ARID_WIDTH,M_AXIMM_94_ARID_WIDTH,M_AXIMM_93_ARID_WIDTH,M_AXIMM_92_ARID_WIDTH,M_AXIMM_91_ARID_WIDTH,M_AXIMM_90_ARID_WIDTH,M_AXIMM_89_ARID_WIDTH,M_AXIMM_88_ARID_WIDTH,M_AXIMM_87_ARID_WIDTH,M_AXIMM_86_ARID_WIDTH,M_AXIMM_85_ARID_WIDTH,M_AXIMM_84_ARID_WIDTH,M_AXIMM_83_ARID_WIDTH,M_AXIMM_82_ARID_WIDTH,M_AXIMM_81_ARID_WIDTH,M_AXIMM_80_ARID_WIDTH,M_AXIMM_79_ARID_WIDTH,M_AXIMM_78_ARID_WIDTH,M_AXIMM_77_ARID_WIDTH,M_AXIMM_76_ARID_WIDTH,M_AXIMM_75_ARID_WIDTH,M_AXIMM_74_ARID_WIDTH,M_AXIMM_73_ARID_WIDTH,M_AXIMM_72_ARID_WIDTH,M_AXIMM_71_ARID_WIDTH,M_AXIMM_70_ARID_WIDTH,M_AXIMM_69_ARID_WIDTH,M_AXIMM_68_ARID_WIDTH,M_AXIMM_67_ARID_WIDTH,M_AXIMM_66_ARID_WIDTH,M_AXIMM_65_ARID_WIDTH,M_AXIMM_64_ARID_WIDTH,M_AXIMM_63_ARID_WIDTH,M_AXIMM_62_ARID_WIDTH,M_AXIMM_61_ARID_WIDTH,M_AXIMM_60_ARID_WIDTH,M_AXIMM_59_ARID_WIDTH,M_AXIMM_58_ARID_WIDTH,M_AXIMM_57_ARID_WIDTH,M_AXIMM_56_ARID_WIDTH,M_AXIMM_55_ARID_WIDTH,M_AXIMM_54_ARID_WIDTH,M_AXIMM_53_ARID_WIDTH,M_AXIMM_52_ARID_WIDTH,M_AXIMM_51_ARID_WIDTH,M_AXIMM_50_ARID_WIDTH,M_AXIMM_49_ARID_WIDTH,M_AXIMM_48_ARID_WIDTH,M_AXIMM_47_ARID_WIDTH,M_AXIMM_46_ARID_WIDTH,M_AXIMM_45_ARID_WIDTH,M_AXIMM_44_ARID_WIDTH,M_AXIMM_43_ARID_WIDTH,M_AXIMM_42_ARID_WIDTH,M_AXIMM_41_ARID_WIDTH,M_AXIMM_40_ARID_WIDTH,M_AXIMM_39_ARID_WIDTH,M_AXIMM_38_ARID_WIDTH,M_AXIMM_37_ARID_WIDTH,M_AXIMM_36_ARID_WIDTH,M_AXIMM_35_ARID_WIDTH,M_AXIMM_34_ARID_WIDTH,M_AXIMM_33_ARID_WIDTH,M_AXIMM_32_ARID_WIDTH,M_AXIMM_31_ARID_WIDTH,M_AXIMM_30_ARID_WIDTH,M_AXIMM_29_ARID_WIDTH,M_AXIMM_28_ARID_WIDTH,M_AXIMM_27_ARID_WIDTH,M_AXIMM_26_ARID_WIDTH,M_AXIMM_25_ARID_WIDTH,M_AXIMM_24_ARID_WIDTH,M_AXIMM_23_ARID_WIDTH,M_AXIMM_22_ARID_WIDTH,M_AXIMM_21_ARID_WIDTH,M_AXIMM_20_ARID_WIDTH,M_AXIMM_19_ARID_WIDTH,M_AXIMM_18_ARID_WIDTH,M_AXIMM_17_ARID_WIDTH,M_AXIMM_16_ARID_WIDTH,M_AXIMM_15_ARID_WIDTH,M_AXIMM_14_ARID_WIDTH,M_AXIMM_13_ARID_WIDTH,M_AXIMM_12_ARID_WIDTH,M_AXIMM_11_ARID_WIDTH,M_AXIMM_10_ARID_WIDTH,M_AXIMM_9_ARID_WIDTH,M_AXIMM_8_ARID_WIDTH,M_AXIMM_7_ARID_WIDTH,M_AXIMM_6_ARID_WIDTH,M_AXIMM_5_ARID_WIDTH,M_AXIMM_4_ARID_WIDTH,M_AXIMM_3_ARID_WIDTH,M_AXIMM_2_ARID_WIDTH,M_AXIMM_1_ARID_WIDTH,M_AXIMM_0_ARID_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_AWID_ARRAY = {M_AXIMM_127_AWID_WIDTH,M_AXIMM_126_AWID_WIDTH,M_AXIMM_125_AWID_WIDTH,M_AXIMM_124_AWID_WIDTH,M_AXIMM_123_AWID_WIDTH,M_AXIMM_122_AWID_WIDTH,M_AXIMM_121_AWID_WIDTH,M_AXIMM_120_AWID_WIDTH,M_AXIMM_119_AWID_WIDTH,M_AXIMM_118_AWID_WIDTH,M_AXIMM_117_AWID_WIDTH,M_AXIMM_116_AWID_WIDTH,M_AXIMM_115_AWID_WIDTH,M_AXIMM_114_AWID_WIDTH,M_AXIMM_113_AWID_WIDTH,M_AXIMM_112_AWID_WIDTH,M_AXIMM_111_AWID_WIDTH,M_AXIMM_110_AWID_WIDTH,M_AXIMM_109_AWID_WIDTH,M_AXIMM_108_AWID_WIDTH,M_AXIMM_107_AWID_WIDTH,M_AXIMM_106_AWID_WIDTH,M_AXIMM_105_AWID_WIDTH,M_AXIMM_104_AWID_WIDTH,M_AXIMM_103_AWID_WIDTH,M_AXIMM_102_AWID_WIDTH,M_AXIMM_101_AWID_WIDTH,M_AXIMM_100_AWID_WIDTH,M_AXIMM_99_AWID_WIDTH,M_AXIMM_98_AWID_WIDTH,M_AXIMM_97_AWID_WIDTH,M_AXIMM_96_AWID_WIDTH,M_AXIMM_95_AWID_WIDTH,M_AXIMM_94_AWID_WIDTH,M_AXIMM_93_AWID_WIDTH,M_AXIMM_92_AWID_WIDTH,M_AXIMM_91_AWID_WIDTH,M_AXIMM_90_AWID_WIDTH,M_AXIMM_89_AWID_WIDTH,M_AXIMM_88_AWID_WIDTH,M_AXIMM_87_AWID_WIDTH,M_AXIMM_86_AWID_WIDTH,M_AXIMM_85_AWID_WIDTH,M_AXIMM_84_AWID_WIDTH,M_AXIMM_83_AWID_WIDTH,M_AXIMM_82_AWID_WIDTH,M_AXIMM_81_AWID_WIDTH,M_AXIMM_80_AWID_WIDTH,M_AXIMM_79_AWID_WIDTH,M_AXIMM_78_AWID_WIDTH,M_AXIMM_77_AWID_WIDTH,M_AXIMM_76_AWID_WIDTH,M_AXIMM_75_AWID_WIDTH,M_AXIMM_74_AWID_WIDTH,M_AXIMM_73_AWID_WIDTH,M_AXIMM_72_AWID_WIDTH,M_AXIMM_71_AWID_WIDTH,M_AXIMM_70_AWID_WIDTH,M_AXIMM_69_AWID_WIDTH,M_AXIMM_68_AWID_WIDTH,M_AXIMM_67_AWID_WIDTH,M_AXIMM_66_AWID_WIDTH,M_AXIMM_65_AWID_WIDTH,M_AXIMM_64_AWID_WIDTH,M_AXIMM_63_AWID_WIDTH,M_AXIMM_62_AWID_WIDTH,M_AXIMM_61_AWID_WIDTH,M_AXIMM_60_AWID_WIDTH,M_AXIMM_59_AWID_WIDTH,M_AXIMM_58_AWID_WIDTH,M_AXIMM_57_AWID_WIDTH,M_AXIMM_56_AWID_WIDTH,M_AXIMM_55_AWID_WIDTH,M_AXIMM_54_AWID_WIDTH,M_AXIMM_53_AWID_WIDTH,M_AXIMM_52_AWID_WIDTH,M_AXIMM_51_AWID_WIDTH,M_AXIMM_50_AWID_WIDTH,M_AXIMM_49_AWID_WIDTH,M_AXIMM_48_AWID_WIDTH,M_AXIMM_47_AWID_WIDTH,M_AXIMM_46_AWID_WIDTH,M_AXIMM_45_AWID_WIDTH,M_AXIMM_44_AWID_WIDTH,M_AXIMM_43_AWID_WIDTH,M_AXIMM_42_AWID_WIDTH,M_AXIMM_41_AWID_WIDTH,M_AXIMM_40_AWID_WIDTH,M_AXIMM_39_AWID_WIDTH,M_AXIMM_38_AWID_WIDTH,M_AXIMM_37_AWID_WIDTH,M_AXIMM_36_AWID_WIDTH,M_AXIMM_35_AWID_WIDTH,M_AXIMM_34_AWID_WIDTH,M_AXIMM_33_AWID_WIDTH,M_AXIMM_32_AWID_WIDTH,M_AXIMM_31_AWID_WIDTH,M_AXIMM_30_AWID_WIDTH,M_AXIMM_29_AWID_WIDTH,M_AXIMM_28_AWID_WIDTH,M_AXIMM_27_AWID_WIDTH,M_AXIMM_26_AWID_WIDTH,M_AXIMM_25_AWID_WIDTH,M_AXIMM_24_AWID_WIDTH,M_AXIMM_23_AWID_WIDTH,M_AXIMM_22_AWID_WIDTH,M_AXIMM_21_AWID_WIDTH,M_AXIMM_20_AWID_WIDTH,M_AXIMM_19_AWID_WIDTH,M_AXIMM_18_AWID_WIDTH,M_AXIMM_17_AWID_WIDTH,M_AXIMM_16_AWID_WIDTH,M_AXIMM_15_AWID_WIDTH,M_AXIMM_14_AWID_WIDTH,M_AXIMM_13_AWID_WIDTH,M_AXIMM_12_AWID_WIDTH,M_AXIMM_11_AWID_WIDTH,M_AXIMM_10_AWID_WIDTH,M_AXIMM_9_AWID_WIDTH,M_AXIMM_8_AWID_WIDTH,M_AXIMM_7_AWID_WIDTH,M_AXIMM_6_AWID_WIDTH,M_AXIMM_5_AWID_WIDTH,M_AXIMM_4_AWID_WIDTH,M_AXIMM_3_AWID_WIDTH,M_AXIMM_2_AWID_WIDTH,M_AXIMM_1_AWID_WIDTH,M_AXIMM_0_AWID_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_BID_ARRAY = {M_AXIMM_127_BID_WIDTH,M_AXIMM_126_BID_WIDTH,M_AXIMM_125_BID_WIDTH,M_AXIMM_124_BID_WIDTH,M_AXIMM_123_BID_WIDTH,M_AXIMM_122_BID_WIDTH,M_AXIMM_121_BID_WIDTH,M_AXIMM_120_BID_WIDTH,M_AXIMM_119_BID_WIDTH,M_AXIMM_118_BID_WIDTH,M_AXIMM_117_BID_WIDTH,M_AXIMM_116_BID_WIDTH,M_AXIMM_115_BID_WIDTH,M_AXIMM_114_BID_WIDTH,M_AXIMM_113_BID_WIDTH,M_AXIMM_112_BID_WIDTH,M_AXIMM_111_BID_WIDTH,M_AXIMM_110_BID_WIDTH,M_AXIMM_109_BID_WIDTH,M_AXIMM_108_BID_WIDTH,M_AXIMM_107_BID_WIDTH,M_AXIMM_106_BID_WIDTH,M_AXIMM_105_BID_WIDTH,M_AXIMM_104_BID_WIDTH,M_AXIMM_103_BID_WIDTH,M_AXIMM_102_BID_WIDTH,M_AXIMM_101_BID_WIDTH,M_AXIMM_100_BID_WIDTH,M_AXIMM_99_BID_WIDTH,M_AXIMM_98_BID_WIDTH,M_AXIMM_97_BID_WIDTH,M_AXIMM_96_BID_WIDTH,M_AXIMM_95_BID_WIDTH,M_AXIMM_94_BID_WIDTH,M_AXIMM_93_BID_WIDTH,M_AXIMM_92_BID_WIDTH,M_AXIMM_91_BID_WIDTH,M_AXIMM_90_BID_WIDTH,M_AXIMM_89_BID_WIDTH,M_AXIMM_88_BID_WIDTH,M_AXIMM_87_BID_WIDTH,M_AXIMM_86_BID_WIDTH,M_AXIMM_85_BID_WIDTH,M_AXIMM_84_BID_WIDTH,M_AXIMM_83_BID_WIDTH,M_AXIMM_82_BID_WIDTH,M_AXIMM_81_BID_WIDTH,M_AXIMM_80_BID_WIDTH,M_AXIMM_79_BID_WIDTH,M_AXIMM_78_BID_WIDTH,M_AXIMM_77_BID_WIDTH,M_AXIMM_76_BID_WIDTH,M_AXIMM_75_BID_WIDTH,M_AXIMM_74_BID_WIDTH,M_AXIMM_73_BID_WIDTH,M_AXIMM_72_BID_WIDTH,M_AXIMM_71_BID_WIDTH,M_AXIMM_70_BID_WIDTH,M_AXIMM_69_BID_WIDTH,M_AXIMM_68_BID_WIDTH,M_AXIMM_67_BID_WIDTH,M_AXIMM_66_BID_WIDTH,M_AXIMM_65_BID_WIDTH,M_AXIMM_64_BID_WIDTH,M_AXIMM_63_BID_WIDTH,M_AXIMM_62_BID_WIDTH,M_AXIMM_61_BID_WIDTH,M_AXIMM_60_BID_WIDTH,M_AXIMM_59_BID_WIDTH,M_AXIMM_58_BID_WIDTH,M_AXIMM_57_BID_WIDTH,M_AXIMM_56_BID_WIDTH,M_AXIMM_55_BID_WIDTH,M_AXIMM_54_BID_WIDTH,M_AXIMM_53_BID_WIDTH,M_AXIMM_52_BID_WIDTH,M_AXIMM_51_BID_WIDTH,M_AXIMM_50_BID_WIDTH,M_AXIMM_49_BID_WIDTH,M_AXIMM_48_BID_WIDTH,M_AXIMM_47_BID_WIDTH,M_AXIMM_46_BID_WIDTH,M_AXIMM_45_BID_WIDTH,M_AXIMM_44_BID_WIDTH,M_AXIMM_43_BID_WIDTH,M_AXIMM_42_BID_WIDTH,M_AXIMM_41_BID_WIDTH,M_AXIMM_40_BID_WIDTH,M_AXIMM_39_BID_WIDTH,M_AXIMM_38_BID_WIDTH,M_AXIMM_37_BID_WIDTH,M_AXIMM_36_BID_WIDTH,M_AXIMM_35_BID_WIDTH,M_AXIMM_34_BID_WIDTH,M_AXIMM_33_BID_WIDTH,M_AXIMM_32_BID_WIDTH,M_AXIMM_31_BID_WIDTH,M_AXIMM_30_BID_WIDTH,M_AXIMM_29_BID_WIDTH,M_AXIMM_28_BID_WIDTH,M_AXIMM_27_BID_WIDTH,M_AXIMM_26_BID_WIDTH,M_AXIMM_25_BID_WIDTH,M_AXIMM_24_BID_WIDTH,M_AXIMM_23_BID_WIDTH,M_AXIMM_22_BID_WIDTH,M_AXIMM_21_BID_WIDTH,M_AXIMM_20_BID_WIDTH,M_AXIMM_19_BID_WIDTH,M_AXIMM_18_BID_WIDTH,M_AXIMM_17_BID_WIDTH,M_AXIMM_16_BID_WIDTH,M_AXIMM_15_BID_WIDTH,M_AXIMM_14_BID_WIDTH,M_AXIMM_13_BID_WIDTH,M_AXIMM_12_BID_WIDTH,M_AXIMM_11_BID_WIDTH,M_AXIMM_10_BID_WIDTH,M_AXIMM_9_BID_WIDTH,M_AXIMM_8_BID_WIDTH,M_AXIMM_7_BID_WIDTH,M_AXIMM_6_BID_WIDTH,M_AXIMM_5_BID_WIDTH,M_AXIMM_4_BID_WIDTH,M_AXIMM_3_BID_WIDTH,M_AXIMM_2_BID_WIDTH,M_AXIMM_1_BID_WIDTH,M_AXIMM_0_BID_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_RID_ARRAY = {M_AXIMM_127_RID_WIDTH,M_AXIMM_126_RID_WIDTH,M_AXIMM_125_RID_WIDTH,M_AXIMM_124_RID_WIDTH,M_AXIMM_123_RID_WIDTH,M_AXIMM_122_RID_WIDTH,M_AXIMM_121_RID_WIDTH,M_AXIMM_120_RID_WIDTH,M_AXIMM_119_RID_WIDTH,M_AXIMM_118_RID_WIDTH,M_AXIMM_117_RID_WIDTH,M_AXIMM_116_RID_WIDTH,M_AXIMM_115_RID_WIDTH,M_AXIMM_114_RID_WIDTH,M_AXIMM_113_RID_WIDTH,M_AXIMM_112_RID_WIDTH,M_AXIMM_111_RID_WIDTH,M_AXIMM_110_RID_WIDTH,M_AXIMM_109_RID_WIDTH,M_AXIMM_108_RID_WIDTH,M_AXIMM_107_RID_WIDTH,M_AXIMM_106_RID_WIDTH,M_AXIMM_105_RID_WIDTH,M_AXIMM_104_RID_WIDTH,M_AXIMM_103_RID_WIDTH,M_AXIMM_102_RID_WIDTH,M_AXIMM_101_RID_WIDTH,M_AXIMM_100_RID_WIDTH,M_AXIMM_99_RID_WIDTH,M_AXIMM_98_RID_WIDTH,M_AXIMM_97_RID_WIDTH,M_AXIMM_96_RID_WIDTH,M_AXIMM_95_RID_WIDTH,M_AXIMM_94_RID_WIDTH,M_AXIMM_93_RID_WIDTH,M_AXIMM_92_RID_WIDTH,M_AXIMM_91_RID_WIDTH,M_AXIMM_90_RID_WIDTH,M_AXIMM_89_RID_WIDTH,M_AXIMM_88_RID_WIDTH,M_AXIMM_87_RID_WIDTH,M_AXIMM_86_RID_WIDTH,M_AXIMM_85_RID_WIDTH,M_AXIMM_84_RID_WIDTH,M_AXIMM_83_RID_WIDTH,M_AXIMM_82_RID_WIDTH,M_AXIMM_81_RID_WIDTH,M_AXIMM_80_RID_WIDTH,M_AXIMM_79_RID_WIDTH,M_AXIMM_78_RID_WIDTH,M_AXIMM_77_RID_WIDTH,M_AXIMM_76_RID_WIDTH,M_AXIMM_75_RID_WIDTH,M_AXIMM_74_RID_WIDTH,M_AXIMM_73_RID_WIDTH,M_AXIMM_72_RID_WIDTH,M_AXIMM_71_RID_WIDTH,M_AXIMM_70_RID_WIDTH,M_AXIMM_69_RID_WIDTH,M_AXIMM_68_RID_WIDTH,M_AXIMM_67_RID_WIDTH,M_AXIMM_66_RID_WIDTH,M_AXIMM_65_RID_WIDTH,M_AXIMM_64_RID_WIDTH,M_AXIMM_63_RID_WIDTH,M_AXIMM_62_RID_WIDTH,M_AXIMM_61_RID_WIDTH,M_AXIMM_60_RID_WIDTH,M_AXIMM_59_RID_WIDTH,M_AXIMM_58_RID_WIDTH,M_AXIMM_57_RID_WIDTH,M_AXIMM_56_RID_WIDTH,M_AXIMM_55_RID_WIDTH,M_AXIMM_54_RID_WIDTH,M_AXIMM_53_RID_WIDTH,M_AXIMM_52_RID_WIDTH,M_AXIMM_51_RID_WIDTH,M_AXIMM_50_RID_WIDTH,M_AXIMM_49_RID_WIDTH,M_AXIMM_48_RID_WIDTH,M_AXIMM_47_RID_WIDTH,M_AXIMM_46_RID_WIDTH,M_AXIMM_45_RID_WIDTH,M_AXIMM_44_RID_WIDTH,M_AXIMM_43_RID_WIDTH,M_AXIMM_42_RID_WIDTH,M_AXIMM_41_RID_WIDTH,M_AXIMM_40_RID_WIDTH,M_AXIMM_39_RID_WIDTH,M_AXIMM_38_RID_WIDTH,M_AXIMM_37_RID_WIDTH,M_AXIMM_36_RID_WIDTH,M_AXIMM_35_RID_WIDTH,M_AXIMM_34_RID_WIDTH,M_AXIMM_33_RID_WIDTH,M_AXIMM_32_RID_WIDTH,M_AXIMM_31_RID_WIDTH,M_AXIMM_30_RID_WIDTH,M_AXIMM_29_RID_WIDTH,M_AXIMM_28_RID_WIDTH,M_AXIMM_27_RID_WIDTH,M_AXIMM_26_RID_WIDTH,M_AXIMM_25_RID_WIDTH,M_AXIMM_24_RID_WIDTH,M_AXIMM_23_RID_WIDTH,M_AXIMM_22_RID_WIDTH,M_AXIMM_21_RID_WIDTH,M_AXIMM_20_RID_WIDTH,M_AXIMM_19_RID_WIDTH,M_AXIMM_18_RID_WIDTH,M_AXIMM_17_RID_WIDTH,M_AXIMM_16_RID_WIDTH,M_AXIMM_15_RID_WIDTH,M_AXIMM_14_RID_WIDTH,M_AXIMM_13_RID_WIDTH,M_AXIMM_12_RID_WIDTH,M_AXIMM_11_RID_WIDTH,M_AXIMM_10_RID_WIDTH,M_AXIMM_9_RID_WIDTH,M_AXIMM_8_RID_WIDTH,M_AXIMM_7_RID_WIDTH,M_AXIMM_6_RID_WIDTH,M_AXIMM_5_RID_WIDTH,M_AXIMM_4_RID_WIDTH,M_AXIMM_3_RID_WIDTH,M_AXIMM_2_RID_WIDTH,M_AXIMM_1_RID_WIDTH,M_AXIMM_0_RID_WIDTH};
    localparam [C_MAX_AXIMMs-1:0] M_AXIMM_WID_ARRAY = {M_AXIMM_127_WID_WIDTH,M_AXIMM_126_WID_WIDTH,M_AXIMM_125_WID_WIDTH,M_AXIMM_124_WID_WIDTH,M_AXIMM_123_WID_WIDTH,M_AXIMM_122_WID_WIDTH,M_AXIMM_121_WID_WIDTH,M_AXIMM_120_WID_WIDTH,M_AXIMM_119_WID_WIDTH,M_AXIMM_118_WID_WIDTH,M_AXIMM_117_WID_WIDTH,M_AXIMM_116_WID_WIDTH,M_AXIMM_115_WID_WIDTH,M_AXIMM_114_WID_WIDTH,M_AXIMM_113_WID_WIDTH,M_AXIMM_112_WID_WIDTH,M_AXIMM_111_WID_WIDTH,M_AXIMM_110_WID_WIDTH,M_AXIMM_109_WID_WIDTH,M_AXIMM_108_WID_WIDTH,M_AXIMM_107_WID_WIDTH,M_AXIMM_106_WID_WIDTH,M_AXIMM_105_WID_WIDTH,M_AXIMM_104_WID_WIDTH,M_AXIMM_103_WID_WIDTH,M_AXIMM_102_WID_WIDTH,M_AXIMM_101_WID_WIDTH,M_AXIMM_100_WID_WIDTH,M_AXIMM_99_WID_WIDTH,M_AXIMM_98_WID_WIDTH,M_AXIMM_97_WID_WIDTH,M_AXIMM_96_WID_WIDTH,M_AXIMM_95_WID_WIDTH,M_AXIMM_94_WID_WIDTH,M_AXIMM_93_WID_WIDTH,M_AXIMM_92_WID_WIDTH,M_AXIMM_91_WID_WIDTH,M_AXIMM_90_WID_WIDTH,M_AXIMM_89_WID_WIDTH,M_AXIMM_88_WID_WIDTH,M_AXIMM_87_WID_WIDTH,M_AXIMM_86_WID_WIDTH,M_AXIMM_85_WID_WIDTH,M_AXIMM_84_WID_WIDTH,M_AXIMM_83_WID_WIDTH,M_AXIMM_82_WID_WIDTH,M_AXIMM_81_WID_WIDTH,M_AXIMM_80_WID_WIDTH,M_AXIMM_79_WID_WIDTH,M_AXIMM_78_WID_WIDTH,M_AXIMM_77_WID_WIDTH,M_AXIMM_76_WID_WIDTH,M_AXIMM_75_WID_WIDTH,M_AXIMM_74_WID_WIDTH,M_AXIMM_73_WID_WIDTH,M_AXIMM_72_WID_WIDTH,M_AXIMM_71_WID_WIDTH,M_AXIMM_70_WID_WIDTH,M_AXIMM_69_WID_WIDTH,M_AXIMM_68_WID_WIDTH,M_AXIMM_67_WID_WIDTH,M_AXIMM_66_WID_WIDTH,M_AXIMM_65_WID_WIDTH,M_AXIMM_64_WID_WIDTH,M_AXIMM_63_WID_WIDTH,M_AXIMM_62_WID_WIDTH,M_AXIMM_61_WID_WIDTH,M_AXIMM_60_WID_WIDTH,M_AXIMM_59_WID_WIDTH,M_AXIMM_58_WID_WIDTH,M_AXIMM_57_WID_WIDTH,M_AXIMM_56_WID_WIDTH,M_AXIMM_55_WID_WIDTH,M_AXIMM_54_WID_WIDTH,M_AXIMM_53_WID_WIDTH,M_AXIMM_52_WID_WIDTH,M_AXIMM_51_WID_WIDTH,M_AXIMM_50_WID_WIDTH,M_AXIMM_49_WID_WIDTH,M_AXIMM_48_WID_WIDTH,M_AXIMM_47_WID_WIDTH,M_AXIMM_46_WID_WIDTH,M_AXIMM_45_WID_WIDTH,M_AXIMM_44_WID_WIDTH,M_AXIMM_43_WID_WIDTH,M_AXIMM_42_WID_WIDTH,M_AXIMM_41_WID_WIDTH,M_AXIMM_40_WID_WIDTH,M_AXIMM_39_WID_WIDTH,M_AXIMM_38_WID_WIDTH,M_AXIMM_37_WID_WIDTH,M_AXIMM_36_WID_WIDTH,M_AXIMM_35_WID_WIDTH,M_AXIMM_34_WID_WIDTH,M_AXIMM_33_WID_WIDTH,M_AXIMM_32_WID_WIDTH,M_AXIMM_31_WID_WIDTH,M_AXIMM_30_WID_WIDTH,M_AXIMM_29_WID_WIDTH,M_AXIMM_28_WID_WIDTH,M_AXIMM_27_WID_WIDTH,M_AXIMM_26_WID_WIDTH,M_AXIMM_25_WID_WIDTH,M_AXIMM_24_WID_WIDTH,M_AXIMM_23_WID_WIDTH,M_AXIMM_22_WID_WIDTH,M_AXIMM_21_WID_WIDTH,M_AXIMM_20_WID_WIDTH,M_AXIMM_19_WID_WIDTH,M_AXIMM_18_WID_WIDTH,M_AXIMM_17_WID_WIDTH,M_AXIMM_16_WID_WIDTH,M_AXIMM_15_WID_WIDTH,M_AXIMM_14_WID_WIDTH,M_AXIMM_13_WID_WIDTH,M_AXIMM_12_WID_WIDTH,M_AXIMM_11_WID_WIDTH,M_AXIMM_10_WID_WIDTH,M_AXIMM_9_WID_WIDTH,M_AXIMM_8_WID_WIDTH,M_AXIMM_7_WID_WIDTH,M_AXIMM_6_WID_WIDTH,M_AXIMM_5_WID_WIDTH,M_AXIMM_4_WID_WIDTH,M_AXIMM_3_WID_WIDTH,M_AXIMM_2_WID_WIDTH,M_AXIMM_1_WID_WIDTH,M_AXIMM_0_WID_WIDTH};
    
    wire [M_AXIMM_ADDR_WIDTH-1:0]   ap_AWADDR [C_NUM_AXIMMs-1:0];
    wire [7:0] ap_AWLEN [C_NUM_AXIMMs-1:0];
    wire [2:0] ap_AWSIZE [C_NUM_AXIMMs-1:0];
    wire [1:0] ap_AWBURST [C_NUM_AXIMMs-1:0];
    wire [1:0] ap_AWLOCK [C_NUM_AXIMMs-1:0];
    wire [3:0] ap_AWCACHE [C_NUM_AXIMMs-1:0];
    wire [2:0] ap_AWPROT [C_NUM_AXIMMs-1:0];
    wire [3:0] ap_AWREGION [C_NUM_AXIMMs-1:0];
    wire [3:0] ap_AWQOS [C_NUM_AXIMMs-1:0];
    wire       ap_AWVALID [C_NUM_AXIMMs-1:0];
    wire       ap_AWREADY [C_NUM_AXIMMs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0]   ap_WDATA [C_NUM_AXIMMs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] ap_WSTRB [C_NUM_AXIMMs-1:0];
    wire       ap_WLAST [C_NUM_AXIMMs-1:0];
    wire       ap_WVALID [C_NUM_AXIMMs-1:0];
    wire       ap_WREADY [C_NUM_AXIMMs-1:0];
    wire [1:0] ap_BRESP [C_NUM_AXIMMs-1:0];
    wire       ap_BVALID [C_NUM_AXIMMs-1:0];
    wire       ap_BREADY [C_NUM_AXIMMs-1:0];
    wire [M_AXIMM_ADDR_WIDTH-1:0]   ap_ARADDR [C_NUM_AXIMMs-1:0];
    wire [7:0] ap_ARLEN [C_NUM_AXIMMs-1:0];
    wire [2:0] ap_ARSIZE [C_NUM_AXIMMs-1:0];
    wire [1:0] ap_ARBURST [C_NUM_AXIMMs-1:0];
    wire [1:0] ap_ARLOCK [C_NUM_AXIMMs-1:0];
    wire [3:0] ap_ARCACHE [C_NUM_AXIMMs-1:0];
    wire [2:0] ap_ARPROT [C_NUM_AXIMMs-1:0];
    wire [3:0] ap_ARREGION [C_NUM_AXIMMs-1:0];
    wire [3:0] ap_ARQOS [C_NUM_AXIMMs-1:0];
    wire       ap_ARVALID [C_NUM_AXIMMs-1:0];
    wire       ap_ARREADY [C_NUM_AXIMMs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0]   ap_RDATA [C_NUM_AXIMMs-1:0];
    wire [1:0] ap_RRESP [C_NUM_AXIMMs-1:0];
    wire       ap_RLAST [C_NUM_AXIMMs-1:0];
    wire       ap_RVALID [C_NUM_AXIMMs-1:0];
    wire       ap_RREADY [C_NUM_AXIMMs-1:0];
    wire [M_AXIMM_ADDR_WIDTH-1:0]   dm_AWADDR [C_NUM_AXIMMs-1:0];
    wire [7:0] dm_AWLEN [C_NUM_AXIMMs-1:0];
    wire [2:0] dm_AWSIZE [C_NUM_AXIMMs-1:0];
    wire [1:0] dm_AWBURST [C_NUM_AXIMMs-1:0];
    wire [1:0] dm_AWLOCK [C_NUM_AXIMMs-1:0];
    wire [3:0] dm_AWCACHE [C_NUM_AXIMMs-1:0];
    wire [2:0] dm_AWPROT [C_NUM_AXIMMs-1:0];
    wire [3:0] dm_AWREGION [C_NUM_AXIMMs-1:0];
    wire [3:0] dm_AWQOS [C_NUM_AXIMMs-1:0];
    wire       dm_AWVALID [C_NUM_AXIMMs-1:0];
    wire       dm_AWREADY [C_NUM_AXIMMs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0]   dm_WDATA [C_NUM_AXIMMs-1:0];
    wire [C_MAX_BIT_WIDTH/8-1:0] dm_WSTRB [C_NUM_AXIMMs-1:0];
    wire       dm_WLAST [C_NUM_AXIMMs-1:0];
    wire       dm_WVALID [C_NUM_AXIMMs-1:0];
    wire       dm_WREADY [C_NUM_AXIMMs-1:0];
    wire [1:0] dm_BRESP [C_NUM_AXIMMs-1:0];
    wire       dm_BVALID [C_NUM_AXIMMs-1:0];
    wire       dm_BREADY [C_NUM_AXIMMs-1:0];
    wire [M_AXIMM_ADDR_WIDTH-1:0]   dm_ARADDR [C_NUM_AXIMMs-1:0];
    wire [7:0] dm_ARLEN [C_NUM_AXIMMs-1:0];
    wire [2:0] dm_ARSIZE [C_NUM_AXIMMs-1:0];
    wire [1:0] dm_ARBURST [C_NUM_AXIMMs-1:0];
    wire [1:0] dm_ARLOCK [C_NUM_AXIMMs-1:0];
    wire [3:0] dm_ARCACHE [C_NUM_AXIMMs-1:0];
    wire [2:0] dm_ARPROT [C_NUM_AXIMMs-1:0];
    wire [3:0] dm_ARREGION [C_NUM_AXIMMs-1:0];
    wire [3:0] dm_ARQOS [C_NUM_AXIMMs-1:0];
    wire       dm_ARVALID [C_NUM_AXIMMs-1:0];
    wire       dm_ARREADY [C_NUM_AXIMMs-1:0];
    wire [C_MAX_BIT_WIDTH-1:0]   dm_RDATA [C_NUM_AXIMMs-1:0];
    wire [1:0] dm_RRESP [C_NUM_AXIMMs-1:0];
    wire       dm_RLAST [C_NUM_AXIMMs-1:0];
    wire       dm_RVALID [C_NUM_AXIMMs-1:0];
    wire       dm_RREADY [C_NUM_AXIMMs-1:0];
    
    //assign inputs to buses, and buses to outputs
    generate
        if(C_NUM_AXIMMs > 0) begin
            assign ap_AWADDR[0][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_0_AWADDR;
            assign ap_AWLEN[0] = AP_AXIMM_0_AWLEN;
            assign ap_AWSIZE[0] = AP_AXIMM_0_AWSIZE;
            assign ap_AWBURST[0] = AP_AXIMM_0_AWBURST;
            assign ap_AWLOCK[0] = AP_AXIMM_0_AWLOCK;
            assign ap_AWCACHE[0] = AP_AXIMM_0_AWCACHE;
            assign ap_AWPROT[0] = AP_AXIMM_0_AWPROT;
            assign ap_AWREGION[0] = AP_AXIMM_0_AWREGION;
            assign ap_AWQOS[0] = AP_AXIMM_0_AWQOS;
            assign ap_AWVALID[0] = AP_AXIMM_0_AWVALID;
            assign AP_AXIMM_0_AWREADY = ap_AWREADY[0];
            assign ap_WDATA[0][M_AXIMM_0_DATA_WIDTH-1:0] = AP_AXIMM_0_WDATA;
            assign ap_WSTRB[0][M_AXIMM_0_DATA_WIDTH/8-1:0] = AP_AXIMM_0_WSTRB;
            assign ap_WLAST[0] = AP_AXIMM_0_WLAST;
            assign ap_WVALID[0] = AP_AXIMM_0_WVALID;
            assign AP_AXIMM_0_WREADY = ap_WREADY[0];
            assign AP_AXIMM_0_BRESP = ap_BRESP[0];
            assign AP_AXIMM_0_BVALID = ap_BVALID[0];
            assign ap_BREADY[0] = AP_AXIMM_0_BREADY;
            assign ap_ARADDR[0][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_0_ARADDR;
            assign ap_ARLEN[0] = AP_AXIMM_0_ARLEN;
            assign ap_ARSIZE[0] = AP_AXIMM_0_ARSIZE;
            assign ap_ARBURST[0] = AP_AXIMM_0_ARBURST;
            assign ap_ARLOCK[0] = AP_AXIMM_0_ARLOCK;
            assign ap_ARCACHE[0] = AP_AXIMM_0_ARCACHE;
            assign ap_ARPROT[0] = AP_AXIMM_0_ARPROT;
            assign ap_ARREGION[0] = AP_AXIMM_0_ARREGION;
            assign ap_ARQOS[0] = AP_AXIMM_0_ARQOS;
            assign ap_ARVALID[0] = AP_AXIMM_0_ARVALID;
            assign AP_AXIMM_0_ARREADY = ap_ARREADY[0];
            assign AP_AXIMM_0_RDATA = ap_RDATA[0][M_AXIMM_0_DATA_WIDTH-1:0];
            assign AP_AXIMM_0_RRESP = ap_RRESP[0];
            assign AP_AXIMM_0_RLAST = ap_RLAST[0];
            assign AP_AXIMM_0_RVALID = ap_RVALID[0];
            assign ap_RREADY[0] = AP_AXIMM_0_RREADY;
            assign M_AXIMM_0_AWADDR = dm_AWADDR[0][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_0_AWLEN = dm_AWLEN[0];
            assign M_AXIMM_0_AWSIZE = dm_AWSIZE[0];
            assign M_AXIMM_0_AWBURST = dm_AWBURST[0];
            assign M_AXIMM_0_AWLOCK = dm_AWLOCK[0];
            assign M_AXIMM_0_AWCACHE = dm_AWCACHE[0];
            assign M_AXIMM_0_AWPROT = dm_AWPROT[0];
            assign M_AXIMM_0_AWREGION = dm_AWREGION[0];
            assign M_AXIMM_0_AWQOS = dm_AWQOS[0];
            assign M_AXIMM_0_AWVALID = dm_AWVALID[0];
            assign dm_AWREADY[0] = M_AXIMM_0_AWREADY;
            assign M_AXIMM_0_WDATA = dm_WDATA[0][M_AXIMM_0_DATA_WIDTH-1:0];
            assign M_AXIMM_0_WSTRB = dm_WSTRB[0][M_AXIMM_0_DATA_WIDTH/8-1:0];
            assign M_AXIMM_0_WLAST = dm_WLAST[0];
            assign M_AXIMM_0_WVALID = dm_WVALID[0];
            assign dm_WREADY[0] = M_AXIMM_0_WREADY;
            assign dm_BRESP[0] = M_AXIMM_0_BRESP;
            assign dm_BVALID[0] = M_AXIMM_0_BVALID;
            assign M_AXIMM_0_BREADY = dm_BREADY[0];
            assign M_AXIMM_0_ARADDR = dm_ARADDR[0][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_0_ARLEN = dm_ARLEN[0];
            assign M_AXIMM_0_ARSIZE = dm_ARSIZE[0];
            assign M_AXIMM_0_ARBURST = dm_ARBURST[0];
            assign M_AXIMM_0_ARLOCK = dm_ARLOCK[0];
            assign M_AXIMM_0_ARCACHE = dm_ARCACHE[0];
            assign M_AXIMM_0_ARPROT = dm_ARPROT[0];
            assign M_AXIMM_0_ARREGION = dm_ARREGION[0];
            assign M_AXIMM_0_ARQOS = dm_ARQOS[0];
            assign M_AXIMM_0_ARVALID = dm_ARVALID[0];
            assign dm_ARREADY[0] = M_AXIMM_0_ARREADY;
            assign dm_RDATA[0][M_AXIMM_0_DATA_WIDTH-1:0] = M_AXIMM_0_RDATA;
            assign dm_RRESP[0] = M_AXIMM_0_RRESP;
            assign dm_RLAST[0] = M_AXIMM_0_RLAST;
            assign dm_RVALID[0] = M_AXIMM_0_RVALID;
            assign M_AXIMM_0_RREADY = dm_RREADY[0];
        end
        if(C_NUM_AXIMMs > 1) begin
            assign ap_AWADDR[1][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_1_AWADDR;
            assign ap_AWLEN[1] = AP_AXIMM_1_AWLEN;
            assign ap_AWSIZE[1] = AP_AXIMM_1_AWSIZE;
            assign ap_AWBURST[1] = AP_AXIMM_1_AWBURST;
            assign ap_AWLOCK[1] = AP_AXIMM_1_AWLOCK;
            assign ap_AWCACHE[1] = AP_AXIMM_1_AWCACHE;
            assign ap_AWPROT[1] = AP_AXIMM_1_AWPROT;
            assign ap_AWREGION[1] = AP_AXIMM_1_AWREGION;
            assign ap_AWQOS[1] = AP_AXIMM_1_AWQOS;
            assign ap_AWVALID[1] = AP_AXIMM_1_AWVALID;
            assign AP_AXIMM_1_AWREADY = ap_AWREADY[1];
            assign ap_WDATA[1][M_AXIMM_1_DATA_WIDTH-1:0] = AP_AXIMM_1_WDATA;
            assign ap_WSTRB[1][M_AXIMM_1_DATA_WIDTH/8-1:0] = AP_AXIMM_1_WSTRB;
            assign ap_WLAST[1] = AP_AXIMM_1_WLAST;
            assign ap_WVALID[1] = AP_AXIMM_1_WVALID;
            assign AP_AXIMM_1_WREADY = ap_WREADY[1];
            assign AP_AXIMM_1_BRESP = ap_BRESP[1];
            assign AP_AXIMM_1_BVALID = ap_BVALID[1];
            assign ap_BREADY[1] = AP_AXIMM_1_BREADY;
            assign ap_ARADDR[1][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_1_ARADDR;
            assign ap_ARLEN[1] = AP_AXIMM_1_ARLEN;
            assign ap_ARSIZE[1] = AP_AXIMM_1_ARSIZE;
            assign ap_ARBURST[1] = AP_AXIMM_1_ARBURST;
            assign ap_ARLOCK[1] = AP_AXIMM_1_ARLOCK;
            assign ap_ARCACHE[1] = AP_AXIMM_1_ARCACHE;
            assign ap_ARPROT[1] = AP_AXIMM_1_ARPROT;
            assign ap_ARREGION[1] = AP_AXIMM_1_ARREGION;
            assign ap_ARQOS[1] = AP_AXIMM_1_ARQOS;
            assign ap_ARVALID[1] = AP_AXIMM_1_ARVALID;
            assign AP_AXIMM_1_ARREADY = ap_ARREADY[1];
            assign AP_AXIMM_1_RDATA = ap_RDATA[1][M_AXIMM_1_DATA_WIDTH-1:0];
            assign AP_AXIMM_1_RRESP = ap_RRESP[1];
            assign AP_AXIMM_1_RLAST = ap_RLAST[1];
            assign AP_AXIMM_1_RVALID = ap_RVALID[1];
            assign ap_RREADY[1] = AP_AXIMM_1_RREADY;
            assign M_AXIMM_1_AWADDR = dm_AWADDR[1][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_1_AWLEN = dm_AWLEN[1];
            assign M_AXIMM_1_AWSIZE = dm_AWSIZE[1];
            assign M_AXIMM_1_AWBURST = dm_AWBURST[1];
            assign M_AXIMM_1_AWLOCK = dm_AWLOCK[1];
            assign M_AXIMM_1_AWCACHE = dm_AWCACHE[1];
            assign M_AXIMM_1_AWPROT = dm_AWPROT[1];
            assign M_AXIMM_1_AWREGION = dm_AWREGION[1];
            assign M_AXIMM_1_AWQOS = dm_AWQOS[1];
            assign M_AXIMM_1_AWVALID = dm_AWVALID[1];
            assign dm_AWREADY[1] = M_AXIMM_1_AWREADY;
            assign M_AXIMM_1_WDATA = dm_WDATA[1][M_AXIMM_1_DATA_WIDTH-1:0];
            assign M_AXIMM_1_WSTRB = dm_WSTRB[1][M_AXIMM_1_DATA_WIDTH/8-1:0];
            assign M_AXIMM_1_WLAST = dm_WLAST[1];
            assign M_AXIMM_1_WVALID = dm_WVALID[1];
            assign dm_WREADY[1] = M_AXIMM_1_WREADY;
            assign dm_BRESP[1] = M_AXIMM_1_BRESP;
            assign dm_BVALID[1] = M_AXIMM_1_BVALID;
            assign M_AXIMM_1_BREADY = dm_BREADY[1];
            assign M_AXIMM_1_ARADDR = dm_ARADDR[1][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_1_ARLEN = dm_ARLEN[1];
            assign M_AXIMM_1_ARSIZE = dm_ARSIZE[1];
            assign M_AXIMM_1_ARBURST = dm_ARBURST[1];
            assign M_AXIMM_1_ARLOCK = dm_ARLOCK[1];
            assign M_AXIMM_1_ARCACHE = dm_ARCACHE[1];
            assign M_AXIMM_1_ARPROT = dm_ARPROT[1];
            assign M_AXIMM_1_ARREGION = dm_ARREGION[1];
            assign M_AXIMM_1_ARQOS = dm_ARQOS[1];
            assign M_AXIMM_1_ARVALID = dm_ARVALID[1];
            assign dm_ARREADY[1] = M_AXIMM_1_ARREADY;
            assign dm_RDATA[1][M_AXIMM_1_DATA_WIDTH-1:0] = M_AXIMM_1_RDATA;
            assign dm_RRESP[1] = M_AXIMM_1_RRESP;
            assign dm_RLAST[1] = M_AXIMM_1_RLAST;
            assign dm_RVALID[1] = M_AXIMM_1_RVALID;
            assign M_AXIMM_1_RREADY = dm_RREADY[1];
        end
        if(C_NUM_AXIMMs > 2) begin
            assign ap_AWADDR[2][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_2_AWADDR;
            assign ap_AWLEN[2] = AP_AXIMM_2_AWLEN;
            assign ap_AWSIZE[2] = AP_AXIMM_2_AWSIZE;
            assign ap_AWBURST[2] = AP_AXIMM_2_AWBURST;
            assign ap_AWLOCK[2] = AP_AXIMM_2_AWLOCK;
            assign ap_AWCACHE[2] = AP_AXIMM_2_AWCACHE;
            assign ap_AWPROT[2] = AP_AXIMM_2_AWPROT;
            assign ap_AWREGION[2] = AP_AXIMM_2_AWREGION;
            assign ap_AWQOS[2] = AP_AXIMM_2_AWQOS;
            assign ap_AWVALID[2] = AP_AXIMM_2_AWVALID;
            assign AP_AXIMM_2_AWREADY = ap_AWREADY[2];
            assign ap_WDATA[2][M_AXIMM_2_DATA_WIDTH-1:0] = AP_AXIMM_2_WDATA;
            assign ap_WSTRB[2][M_AXIMM_2_DATA_WIDTH/8-1:0] = AP_AXIMM_2_WSTRB;
            assign ap_WLAST[2] = AP_AXIMM_2_WLAST;
            assign ap_WVALID[2] = AP_AXIMM_2_WVALID;
            assign AP_AXIMM_2_WREADY = ap_WREADY[2];
            assign AP_AXIMM_2_BRESP = ap_BRESP[2];
            assign AP_AXIMM_2_BVALID = ap_BVALID[2];
            assign ap_BREADY[2] = AP_AXIMM_2_BREADY;
            assign ap_ARADDR[2][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_2_ARADDR;
            assign ap_ARLEN[2] = AP_AXIMM_2_ARLEN;
            assign ap_ARSIZE[2] = AP_AXIMM_2_ARSIZE;
            assign ap_ARBURST[2] = AP_AXIMM_2_ARBURST;
            assign ap_ARLOCK[2] = AP_AXIMM_2_ARLOCK;
            assign ap_ARCACHE[2] = AP_AXIMM_2_ARCACHE;
            assign ap_ARPROT[2] = AP_AXIMM_2_ARPROT;
            assign ap_ARREGION[2] = AP_AXIMM_2_ARREGION;
            assign ap_ARQOS[2] = AP_AXIMM_2_ARQOS;
            assign ap_ARVALID[2] = AP_AXIMM_2_ARVALID;
            assign AP_AXIMM_2_ARREADY = ap_ARREADY[2];
            assign AP_AXIMM_2_RDATA = ap_RDATA[2][M_AXIMM_2_DATA_WIDTH-1:0];
            assign AP_AXIMM_2_RRESP = ap_RRESP[2];
            assign AP_AXIMM_2_RLAST = ap_RLAST[2];
            assign AP_AXIMM_2_RVALID = ap_RVALID[2];
            assign ap_RREADY[2] = AP_AXIMM_2_RREADY;
            assign M_AXIMM_2_AWADDR = dm_AWADDR[2][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_2_AWLEN = dm_AWLEN[2];
            assign M_AXIMM_2_AWSIZE = dm_AWSIZE[2];
            assign M_AXIMM_2_AWBURST = dm_AWBURST[2];
            assign M_AXIMM_2_AWLOCK = dm_AWLOCK[2];
            assign M_AXIMM_2_AWCACHE = dm_AWCACHE[2];
            assign M_AXIMM_2_AWPROT = dm_AWPROT[2];
            assign M_AXIMM_2_AWREGION = dm_AWREGION[2];
            assign M_AXIMM_2_AWQOS = dm_AWQOS[2];
            assign M_AXIMM_2_AWVALID = dm_AWVALID[2];
            assign dm_AWREADY[2] = M_AXIMM_2_AWREADY;
            assign M_AXIMM_2_WDATA = dm_WDATA[2][M_AXIMM_2_DATA_WIDTH-1:0];
            assign M_AXIMM_2_WSTRB = dm_WSTRB[2][M_AXIMM_2_DATA_WIDTH/8-1:0];
            assign M_AXIMM_2_WLAST = dm_WLAST[2];
            assign M_AXIMM_2_WVALID = dm_WVALID[2];
            assign dm_WREADY[2] = M_AXIMM_2_WREADY;
            assign dm_BRESP[2] = M_AXIMM_2_BRESP;
            assign dm_BVALID[2] = M_AXIMM_2_BVALID;
            assign M_AXIMM_2_BREADY = dm_BREADY[2];
            assign M_AXIMM_2_ARADDR = dm_ARADDR[2][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_2_ARLEN = dm_ARLEN[2];
            assign M_AXIMM_2_ARSIZE = dm_ARSIZE[2];
            assign M_AXIMM_2_ARBURST = dm_ARBURST[2];
            assign M_AXIMM_2_ARLOCK = dm_ARLOCK[2];
            assign M_AXIMM_2_ARCACHE = dm_ARCACHE[2];
            assign M_AXIMM_2_ARPROT = dm_ARPROT[2];
            assign M_AXIMM_2_ARREGION = dm_ARREGION[2];
            assign M_AXIMM_2_ARQOS = dm_ARQOS[2];
            assign M_AXIMM_2_ARVALID = dm_ARVALID[2];
            assign dm_ARREADY[2] = M_AXIMM_2_ARREADY;
            assign dm_RDATA[2][M_AXIMM_2_DATA_WIDTH-1:0] = M_AXIMM_2_RDATA;
            assign dm_RRESP[2] = M_AXIMM_2_RRESP;
            assign dm_RLAST[2] = M_AXIMM_2_RLAST;
            assign dm_RVALID[2] = M_AXIMM_2_RVALID;
            assign M_AXIMM_2_RREADY = dm_RREADY[2];
        end
        if(C_NUM_AXIMMs > 3) begin
            assign ap_AWADDR[3][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_3_AWADDR;
            assign ap_AWLEN[3] = AP_AXIMM_3_AWLEN;
            assign ap_AWSIZE[3] = AP_AXIMM_3_AWSIZE;
            assign ap_AWBURST[3] = AP_AXIMM_3_AWBURST;
            assign ap_AWLOCK[3] = AP_AXIMM_3_AWLOCK;
            assign ap_AWCACHE[3] = AP_AXIMM_3_AWCACHE;
            assign ap_AWPROT[3] = AP_AXIMM_3_AWPROT;
            assign ap_AWREGION[3] = AP_AXIMM_3_AWREGION;
            assign ap_AWQOS[3] = AP_AXIMM_3_AWQOS;
            assign ap_AWVALID[3] = AP_AXIMM_3_AWVALID;
            assign AP_AXIMM_3_AWREADY = ap_AWREADY[3];
            assign ap_WDATA[3][M_AXIMM_3_DATA_WIDTH-1:0] = AP_AXIMM_3_WDATA;
            assign ap_WSTRB[3][M_AXIMM_3_DATA_WIDTH/8-1:0] = AP_AXIMM_3_WSTRB;
            assign ap_WLAST[3] = AP_AXIMM_3_WLAST;
            assign ap_WVALID[3] = AP_AXIMM_3_WVALID;
            assign AP_AXIMM_3_WREADY = ap_WREADY[3];
            assign AP_AXIMM_3_BRESP = ap_BRESP[3];
            assign AP_AXIMM_3_BVALID = ap_BVALID[3];
            assign ap_BREADY[3] = AP_AXIMM_3_BREADY;
            assign ap_ARADDR[3][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_3_ARADDR;
            assign ap_ARLEN[3] = AP_AXIMM_3_ARLEN;
            assign ap_ARSIZE[3] = AP_AXIMM_3_ARSIZE;
            assign ap_ARBURST[3] = AP_AXIMM_3_ARBURST;
            assign ap_ARLOCK[3] = AP_AXIMM_3_ARLOCK;
            assign ap_ARCACHE[3] = AP_AXIMM_3_ARCACHE;
            assign ap_ARPROT[3] = AP_AXIMM_3_ARPROT;
            assign ap_ARREGION[3] = AP_AXIMM_3_ARREGION;
            assign ap_ARQOS[3] = AP_AXIMM_3_ARQOS;
            assign ap_ARVALID[3] = AP_AXIMM_3_ARVALID;
            assign AP_AXIMM_3_ARREADY = ap_ARREADY[3];
            assign AP_AXIMM_3_RDATA = ap_RDATA[3][M_AXIMM_3_DATA_WIDTH-1:0];
            assign AP_AXIMM_3_RRESP = ap_RRESP[3];
            assign AP_AXIMM_3_RLAST = ap_RLAST[3];
            assign AP_AXIMM_3_RVALID = ap_RVALID[3];
            assign ap_RREADY[3] = AP_AXIMM_3_RREADY;
            assign M_AXIMM_3_AWADDR = dm_AWADDR[3][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_3_AWLEN = dm_AWLEN[3];
            assign M_AXIMM_3_AWSIZE = dm_AWSIZE[3];
            assign M_AXIMM_3_AWBURST = dm_AWBURST[3];
            assign M_AXIMM_3_AWLOCK = dm_AWLOCK[3];
            assign M_AXIMM_3_AWCACHE = dm_AWCACHE[3];
            assign M_AXIMM_3_AWPROT = dm_AWPROT[3];
            assign M_AXIMM_3_AWREGION = dm_AWREGION[3];
            assign M_AXIMM_3_AWQOS = dm_AWQOS[3];
            assign M_AXIMM_3_AWVALID = dm_AWVALID[3];
            assign dm_AWREADY[3] = M_AXIMM_3_AWREADY;
            assign M_AXIMM_3_WDATA = dm_WDATA[3][M_AXIMM_3_DATA_WIDTH-1:0];
            assign M_AXIMM_3_WSTRB = dm_WSTRB[3][M_AXIMM_3_DATA_WIDTH/8-1:0];
            assign M_AXIMM_3_WLAST = dm_WLAST[3];
            assign M_AXIMM_3_WVALID = dm_WVALID[3];
            assign dm_WREADY[3] = M_AXIMM_3_WREADY;
            assign dm_BRESP[3] = M_AXIMM_3_BRESP;
            assign dm_BVALID[3] = M_AXIMM_3_BVALID;
            assign M_AXIMM_3_BREADY = dm_BREADY[3];
            assign M_AXIMM_3_ARADDR = dm_ARADDR[3][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_3_ARLEN = dm_ARLEN[3];
            assign M_AXIMM_3_ARSIZE = dm_ARSIZE[3];
            assign M_AXIMM_3_ARBURST = dm_ARBURST[3];
            assign M_AXIMM_3_ARLOCK = dm_ARLOCK[3];
            assign M_AXIMM_3_ARCACHE = dm_ARCACHE[3];
            assign M_AXIMM_3_ARPROT = dm_ARPROT[3];
            assign M_AXIMM_3_ARREGION = dm_ARREGION[3];
            assign M_AXIMM_3_ARQOS = dm_ARQOS[3];
            assign M_AXIMM_3_ARVALID = dm_ARVALID[3];
            assign dm_ARREADY[3] = M_AXIMM_3_ARREADY;
            assign dm_RDATA[3][M_AXIMM_3_DATA_WIDTH-1:0] = M_AXIMM_3_RDATA;
            assign dm_RRESP[3] = M_AXIMM_3_RRESP;
            assign dm_RLAST[3] = M_AXIMM_3_RLAST;
            assign dm_RVALID[3] = M_AXIMM_3_RVALID;
            assign M_AXIMM_3_RREADY = dm_RREADY[3];
        end
        if(C_NUM_AXIMMs > 4) begin
            assign ap_AWADDR[4][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_4_AWADDR;
            assign ap_AWLEN[4] = AP_AXIMM_4_AWLEN;
            assign ap_AWSIZE[4] = AP_AXIMM_4_AWSIZE;
            assign ap_AWBURST[4] = AP_AXIMM_4_AWBURST;
            assign ap_AWLOCK[4] = AP_AXIMM_4_AWLOCK;
            assign ap_AWCACHE[4] = AP_AXIMM_4_AWCACHE;
            assign ap_AWPROT[4] = AP_AXIMM_4_AWPROT;
            assign ap_AWREGION[4] = AP_AXIMM_4_AWREGION;
            assign ap_AWQOS[4] = AP_AXIMM_4_AWQOS;
            assign ap_AWVALID[4] = AP_AXIMM_4_AWVALID;
            assign AP_AXIMM_4_AWREADY = ap_AWREADY[4];
            assign ap_WDATA[4][M_AXIMM_4_DATA_WIDTH-1:0] = AP_AXIMM_4_WDATA;
            assign ap_WSTRB[4][M_AXIMM_4_DATA_WIDTH/8-1:0] = AP_AXIMM_4_WSTRB;
            assign ap_WLAST[4] = AP_AXIMM_4_WLAST;
            assign ap_WVALID[4] = AP_AXIMM_4_WVALID;
            assign AP_AXIMM_4_WREADY = ap_WREADY[4];
            assign AP_AXIMM_4_BRESP = ap_BRESP[4];
            assign AP_AXIMM_4_BVALID = ap_BVALID[4];
            assign ap_BREADY[4] = AP_AXIMM_4_BREADY;
            assign ap_ARADDR[4][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_4_ARADDR;
            assign ap_ARLEN[4] = AP_AXIMM_4_ARLEN;
            assign ap_ARSIZE[4] = AP_AXIMM_4_ARSIZE;
            assign ap_ARBURST[4] = AP_AXIMM_4_ARBURST;
            assign ap_ARLOCK[4] = AP_AXIMM_4_ARLOCK;
            assign ap_ARCACHE[4] = AP_AXIMM_4_ARCACHE;
            assign ap_ARPROT[4] = AP_AXIMM_4_ARPROT;
            assign ap_ARREGION[4] = AP_AXIMM_4_ARREGION;
            assign ap_ARQOS[4] = AP_AXIMM_4_ARQOS;
            assign ap_ARVALID[4] = AP_AXIMM_4_ARVALID;
            assign AP_AXIMM_4_ARREADY = ap_ARREADY[4];
            assign AP_AXIMM_4_RDATA = ap_RDATA[4][M_AXIMM_4_DATA_WIDTH-1:0];
            assign AP_AXIMM_4_RRESP = ap_RRESP[4];
            assign AP_AXIMM_4_RLAST = ap_RLAST[4];
            assign AP_AXIMM_4_RVALID = ap_RVALID[4];
            assign ap_RREADY[4] = AP_AXIMM_4_RREADY;
            assign M_AXIMM_4_AWADDR = dm_AWADDR[4][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_4_AWLEN = dm_AWLEN[4];
            assign M_AXIMM_4_AWSIZE = dm_AWSIZE[4];
            assign M_AXIMM_4_AWBURST = dm_AWBURST[4];
            assign M_AXIMM_4_AWLOCK = dm_AWLOCK[4];
            assign M_AXIMM_4_AWCACHE = dm_AWCACHE[4];
            assign M_AXIMM_4_AWPROT = dm_AWPROT[4];
            assign M_AXIMM_4_AWREGION = dm_AWREGION[4];
            assign M_AXIMM_4_AWQOS = dm_AWQOS[4];
            assign M_AXIMM_4_AWVALID = dm_AWVALID[4];
            assign dm_AWREADY[4] = M_AXIMM_4_AWREADY;
            assign M_AXIMM_4_WDATA = dm_WDATA[4][M_AXIMM_4_DATA_WIDTH-1:0];
            assign M_AXIMM_4_WSTRB = dm_WSTRB[4][M_AXIMM_4_DATA_WIDTH/8-1:0];
            assign M_AXIMM_4_WLAST = dm_WLAST[4];
            assign M_AXIMM_4_WVALID = dm_WVALID[4];
            assign dm_WREADY[4] = M_AXIMM_4_WREADY;
            assign dm_BRESP[4] = M_AXIMM_4_BRESP;
            assign dm_BVALID[4] = M_AXIMM_4_BVALID;
            assign M_AXIMM_4_BREADY = dm_BREADY[4];
            assign M_AXIMM_4_ARADDR = dm_ARADDR[4][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_4_ARLEN = dm_ARLEN[4];
            assign M_AXIMM_4_ARSIZE = dm_ARSIZE[4];
            assign M_AXIMM_4_ARBURST = dm_ARBURST[4];
            assign M_AXIMM_4_ARLOCK = dm_ARLOCK[4];
            assign M_AXIMM_4_ARCACHE = dm_ARCACHE[4];
            assign M_AXIMM_4_ARPROT = dm_ARPROT[4];
            assign M_AXIMM_4_ARREGION = dm_ARREGION[4];
            assign M_AXIMM_4_ARQOS = dm_ARQOS[4];
            assign M_AXIMM_4_ARVALID = dm_ARVALID[4];
            assign dm_ARREADY[4] = M_AXIMM_4_ARREADY;
            assign dm_RDATA[4][M_AXIMM_4_DATA_WIDTH-1:0] = M_AXIMM_4_RDATA;
            assign dm_RRESP[4] = M_AXIMM_4_RRESP;
            assign dm_RLAST[4] = M_AXIMM_4_RLAST;
            assign dm_RVALID[4] = M_AXIMM_4_RVALID;
            assign M_AXIMM_4_RREADY = dm_RREADY[4];
        end
        if(C_NUM_AXIMMs > 5) begin
            assign ap_AWADDR[5][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_5_AWADDR;
            assign ap_AWLEN[5] = AP_AXIMM_5_AWLEN;
            assign ap_AWSIZE[5] = AP_AXIMM_5_AWSIZE;
            assign ap_AWBURST[5] = AP_AXIMM_5_AWBURST;
            assign ap_AWLOCK[5] = AP_AXIMM_5_AWLOCK;
            assign ap_AWCACHE[5] = AP_AXIMM_5_AWCACHE;
            assign ap_AWPROT[5] = AP_AXIMM_5_AWPROT;
            assign ap_AWREGION[5] = AP_AXIMM_5_AWREGION;
            assign ap_AWQOS[5] = AP_AXIMM_5_AWQOS;
            assign ap_AWVALID[5] = AP_AXIMM_5_AWVALID;
            assign AP_AXIMM_5_AWREADY = ap_AWREADY[5];
            assign ap_WDATA[5][M_AXIMM_5_DATA_WIDTH-1:0] = AP_AXIMM_5_WDATA;
            assign ap_WSTRB[5][M_AXIMM_5_DATA_WIDTH/8-1:0] = AP_AXIMM_5_WSTRB;
            assign ap_WLAST[5] = AP_AXIMM_5_WLAST;
            assign ap_WVALID[5] = AP_AXIMM_5_WVALID;
            assign AP_AXIMM_5_WREADY = ap_WREADY[5];
            assign AP_AXIMM_5_BRESP = ap_BRESP[5];
            assign AP_AXIMM_5_BVALID = ap_BVALID[5];
            assign ap_BREADY[5] = AP_AXIMM_5_BREADY;
            assign ap_ARADDR[5][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_5_ARADDR;
            assign ap_ARLEN[5] = AP_AXIMM_5_ARLEN;
            assign ap_ARSIZE[5] = AP_AXIMM_5_ARSIZE;
            assign ap_ARBURST[5] = AP_AXIMM_5_ARBURST;
            assign ap_ARLOCK[5] = AP_AXIMM_5_ARLOCK;
            assign ap_ARCACHE[5] = AP_AXIMM_5_ARCACHE;
            assign ap_ARPROT[5] = AP_AXIMM_5_ARPROT;
            assign ap_ARREGION[5] = AP_AXIMM_5_ARREGION;
            assign ap_ARQOS[5] = AP_AXIMM_5_ARQOS;
            assign ap_ARVALID[5] = AP_AXIMM_5_ARVALID;
            assign AP_AXIMM_5_ARREADY = ap_ARREADY[5];
            assign AP_AXIMM_5_RDATA = ap_RDATA[5][M_AXIMM_5_DATA_WIDTH-1:0];
            assign AP_AXIMM_5_RRESP = ap_RRESP[5];
            assign AP_AXIMM_5_RLAST = ap_RLAST[5];
            assign AP_AXIMM_5_RVALID = ap_RVALID[5];
            assign ap_RREADY[5] = AP_AXIMM_5_RREADY;
            assign M_AXIMM_5_AWADDR = dm_AWADDR[5][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_5_AWLEN = dm_AWLEN[5];
            assign M_AXIMM_5_AWSIZE = dm_AWSIZE[5];
            assign M_AXIMM_5_AWBURST = dm_AWBURST[5];
            assign M_AXIMM_5_AWLOCK = dm_AWLOCK[5];
            assign M_AXIMM_5_AWCACHE = dm_AWCACHE[5];
            assign M_AXIMM_5_AWPROT = dm_AWPROT[5];
            assign M_AXIMM_5_AWREGION = dm_AWREGION[5];
            assign M_AXIMM_5_AWQOS = dm_AWQOS[5];
            assign M_AXIMM_5_AWVALID = dm_AWVALID[5];
            assign dm_AWREADY[5] = M_AXIMM_5_AWREADY;
            assign M_AXIMM_5_WDATA = dm_WDATA[5][M_AXIMM_5_DATA_WIDTH-1:0];
            assign M_AXIMM_5_WSTRB = dm_WSTRB[5][M_AXIMM_5_DATA_WIDTH/8-1:0];
            assign M_AXIMM_5_WLAST = dm_WLAST[5];
            assign M_AXIMM_5_WVALID = dm_WVALID[5];
            assign dm_WREADY[5] = M_AXIMM_5_WREADY;
            assign dm_BRESP[5] = M_AXIMM_5_BRESP;
            assign dm_BVALID[5] = M_AXIMM_5_BVALID;
            assign M_AXIMM_5_BREADY = dm_BREADY[5];
            assign M_AXIMM_5_ARADDR = dm_ARADDR[5][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_5_ARLEN = dm_ARLEN[5];
            assign M_AXIMM_5_ARSIZE = dm_ARSIZE[5];
            assign M_AXIMM_5_ARBURST = dm_ARBURST[5];
            assign M_AXIMM_5_ARLOCK = dm_ARLOCK[5];
            assign M_AXIMM_5_ARCACHE = dm_ARCACHE[5];
            assign M_AXIMM_5_ARPROT = dm_ARPROT[5];
            assign M_AXIMM_5_ARREGION = dm_ARREGION[5];
            assign M_AXIMM_5_ARQOS = dm_ARQOS[5];
            assign M_AXIMM_5_ARVALID = dm_ARVALID[5];
            assign dm_ARREADY[5] = M_AXIMM_5_ARREADY;
            assign dm_RDATA[5][M_AXIMM_5_DATA_WIDTH-1:0] = M_AXIMM_5_RDATA;
            assign dm_RRESP[5] = M_AXIMM_5_RRESP;
            assign dm_RLAST[5] = M_AXIMM_5_RLAST;
            assign dm_RVALID[5] = M_AXIMM_5_RVALID;
            assign M_AXIMM_5_RREADY = dm_RREADY[5];
        end
        if(C_NUM_AXIMMs > 6) begin
            assign ap_AWADDR[6][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_6_AWADDR;
            assign ap_AWLEN[6] = AP_AXIMM_6_AWLEN;
            assign ap_AWSIZE[6] = AP_AXIMM_6_AWSIZE;
            assign ap_AWBURST[6] = AP_AXIMM_6_AWBURST;
            assign ap_AWLOCK[6] = AP_AXIMM_6_AWLOCK;
            assign ap_AWCACHE[6] = AP_AXIMM_6_AWCACHE;
            assign ap_AWPROT[6] = AP_AXIMM_6_AWPROT;
            assign ap_AWREGION[6] = AP_AXIMM_6_AWREGION;
            assign ap_AWQOS[6] = AP_AXIMM_6_AWQOS;
            assign ap_AWVALID[6] = AP_AXIMM_6_AWVALID;
            assign AP_AXIMM_6_AWREADY = ap_AWREADY[6];
            assign ap_WDATA[6][M_AXIMM_6_DATA_WIDTH-1:0] = AP_AXIMM_6_WDATA;
            assign ap_WSTRB[6][M_AXIMM_6_DATA_WIDTH/8-1:0] = AP_AXIMM_6_WSTRB;
            assign ap_WLAST[6] = AP_AXIMM_6_WLAST;
            assign ap_WVALID[6] = AP_AXIMM_6_WVALID;
            assign AP_AXIMM_6_WREADY = ap_WREADY[6];
            assign AP_AXIMM_6_BRESP = ap_BRESP[6];
            assign AP_AXIMM_6_BVALID = ap_BVALID[6];
            assign ap_BREADY[6] = AP_AXIMM_6_BREADY;
            assign ap_ARADDR[6][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_6_ARADDR;
            assign ap_ARLEN[6] = AP_AXIMM_6_ARLEN;
            assign ap_ARSIZE[6] = AP_AXIMM_6_ARSIZE;
            assign ap_ARBURST[6] = AP_AXIMM_6_ARBURST;
            assign ap_ARLOCK[6] = AP_AXIMM_6_ARLOCK;
            assign ap_ARCACHE[6] = AP_AXIMM_6_ARCACHE;
            assign ap_ARPROT[6] = AP_AXIMM_6_ARPROT;
            assign ap_ARREGION[6] = AP_AXIMM_6_ARREGION;
            assign ap_ARQOS[6] = AP_AXIMM_6_ARQOS;
            assign ap_ARVALID[6] = AP_AXIMM_6_ARVALID;
            assign AP_AXIMM_6_ARREADY = ap_ARREADY[6];
            assign AP_AXIMM_6_RDATA = ap_RDATA[6][M_AXIMM_6_DATA_WIDTH-1:0];
            assign AP_AXIMM_6_RRESP = ap_RRESP[6];
            assign AP_AXIMM_6_RLAST = ap_RLAST[6];
            assign AP_AXIMM_6_RVALID = ap_RVALID[6];
            assign ap_RREADY[6] = AP_AXIMM_6_RREADY;
            assign M_AXIMM_6_AWADDR = dm_AWADDR[6][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_6_AWLEN = dm_AWLEN[6];
            assign M_AXIMM_6_AWSIZE = dm_AWSIZE[6];
            assign M_AXIMM_6_AWBURST = dm_AWBURST[6];
            assign M_AXIMM_6_AWLOCK = dm_AWLOCK[6];
            assign M_AXIMM_6_AWCACHE = dm_AWCACHE[6];
            assign M_AXIMM_6_AWPROT = dm_AWPROT[6];
            assign M_AXIMM_6_AWREGION = dm_AWREGION[6];
            assign M_AXIMM_6_AWQOS = dm_AWQOS[6];
            assign M_AXIMM_6_AWVALID = dm_AWVALID[6];
            assign dm_AWREADY[6] = M_AXIMM_6_AWREADY;
            assign M_AXIMM_6_WDATA = dm_WDATA[6][M_AXIMM_6_DATA_WIDTH-1:0];
            assign M_AXIMM_6_WSTRB = dm_WSTRB[6][M_AXIMM_6_DATA_WIDTH/8-1:0];
            assign M_AXIMM_6_WLAST = dm_WLAST[6];
            assign M_AXIMM_6_WVALID = dm_WVALID[6];
            assign dm_WREADY[6] = M_AXIMM_6_WREADY;
            assign dm_BRESP[6] = M_AXIMM_6_BRESP;
            assign dm_BVALID[6] = M_AXIMM_6_BVALID;
            assign M_AXIMM_6_BREADY = dm_BREADY[6];
            assign M_AXIMM_6_ARADDR = dm_ARADDR[6][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_6_ARLEN = dm_ARLEN[6];
            assign M_AXIMM_6_ARSIZE = dm_ARSIZE[6];
            assign M_AXIMM_6_ARBURST = dm_ARBURST[6];
            assign M_AXIMM_6_ARLOCK = dm_ARLOCK[6];
            assign M_AXIMM_6_ARCACHE = dm_ARCACHE[6];
            assign M_AXIMM_6_ARPROT = dm_ARPROT[6];
            assign M_AXIMM_6_ARREGION = dm_ARREGION[6];
            assign M_AXIMM_6_ARQOS = dm_ARQOS[6];
            assign M_AXIMM_6_ARVALID = dm_ARVALID[6];
            assign dm_ARREADY[6] = M_AXIMM_6_ARREADY;
            assign dm_RDATA[6][M_AXIMM_6_DATA_WIDTH-1:0] = M_AXIMM_6_RDATA;
            assign dm_RRESP[6] = M_AXIMM_6_RRESP;
            assign dm_RLAST[6] = M_AXIMM_6_RLAST;
            assign dm_RVALID[6] = M_AXIMM_6_RVALID;
            assign M_AXIMM_6_RREADY = dm_RREADY[6];
        end
        if(C_NUM_AXIMMs > 7) begin
            assign ap_AWADDR[7][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_7_AWADDR;
            assign ap_AWLEN[7] = AP_AXIMM_7_AWLEN;
            assign ap_AWSIZE[7] = AP_AXIMM_7_AWSIZE;
            assign ap_AWBURST[7] = AP_AXIMM_7_AWBURST;
            assign ap_AWLOCK[7] = AP_AXIMM_7_AWLOCK;
            assign ap_AWCACHE[7] = AP_AXIMM_7_AWCACHE;
            assign ap_AWPROT[7] = AP_AXIMM_7_AWPROT;
            assign ap_AWREGION[7] = AP_AXIMM_7_AWREGION;
            assign ap_AWQOS[7] = AP_AXIMM_7_AWQOS;
            assign ap_AWVALID[7] = AP_AXIMM_7_AWVALID;
            assign AP_AXIMM_7_AWREADY = ap_AWREADY[7];
            assign ap_WDATA[7][M_AXIMM_7_DATA_WIDTH-1:0] = AP_AXIMM_7_WDATA;
            assign ap_WSTRB[7][M_AXIMM_7_DATA_WIDTH/8-1:0] = AP_AXIMM_7_WSTRB;
            assign ap_WLAST[7] = AP_AXIMM_7_WLAST;
            assign ap_WVALID[7] = AP_AXIMM_7_WVALID;
            assign AP_AXIMM_7_WREADY = ap_WREADY[7];
            assign AP_AXIMM_7_BRESP = ap_BRESP[7];
            assign AP_AXIMM_7_BVALID = ap_BVALID[7];
            assign ap_BREADY[7] = AP_AXIMM_7_BREADY;
            assign ap_ARADDR[7][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_7_ARADDR;
            assign ap_ARLEN[7] = AP_AXIMM_7_ARLEN;
            assign ap_ARSIZE[7] = AP_AXIMM_7_ARSIZE;
            assign ap_ARBURST[7] = AP_AXIMM_7_ARBURST;
            assign ap_ARLOCK[7] = AP_AXIMM_7_ARLOCK;
            assign ap_ARCACHE[7] = AP_AXIMM_7_ARCACHE;
            assign ap_ARPROT[7] = AP_AXIMM_7_ARPROT;
            assign ap_ARREGION[7] = AP_AXIMM_7_ARREGION;
            assign ap_ARQOS[7] = AP_AXIMM_7_ARQOS;
            assign ap_ARVALID[7] = AP_AXIMM_7_ARVALID;
            assign AP_AXIMM_7_ARREADY = ap_ARREADY[7];
            assign AP_AXIMM_7_RDATA = ap_RDATA[7][M_AXIMM_7_DATA_WIDTH-1:0];
            assign AP_AXIMM_7_RRESP = ap_RRESP[7];
            assign AP_AXIMM_7_RLAST = ap_RLAST[7];
            assign AP_AXIMM_7_RVALID = ap_RVALID[7];
            assign ap_RREADY[7] = AP_AXIMM_7_RREADY;
            assign M_AXIMM_7_AWADDR = dm_AWADDR[7][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_7_AWLEN = dm_AWLEN[7];
            assign M_AXIMM_7_AWSIZE = dm_AWSIZE[7];
            assign M_AXIMM_7_AWBURST = dm_AWBURST[7];
            assign M_AXIMM_7_AWLOCK = dm_AWLOCK[7];
            assign M_AXIMM_7_AWCACHE = dm_AWCACHE[7];
            assign M_AXIMM_7_AWPROT = dm_AWPROT[7];
            assign M_AXIMM_7_AWREGION = dm_AWREGION[7];
            assign M_AXIMM_7_AWQOS = dm_AWQOS[7];
            assign M_AXIMM_7_AWVALID = dm_AWVALID[7];
            assign dm_AWREADY[7] = M_AXIMM_7_AWREADY;
            assign M_AXIMM_7_WDATA = dm_WDATA[7][M_AXIMM_7_DATA_WIDTH-1:0];
            assign M_AXIMM_7_WSTRB = dm_WSTRB[7][M_AXIMM_7_DATA_WIDTH/8-1:0];
            assign M_AXIMM_7_WLAST = dm_WLAST[7];
            assign M_AXIMM_7_WVALID = dm_WVALID[7];
            assign dm_WREADY[7] = M_AXIMM_7_WREADY;
            assign dm_BRESP[7] = M_AXIMM_7_BRESP;
            assign dm_BVALID[7] = M_AXIMM_7_BVALID;
            assign M_AXIMM_7_BREADY = dm_BREADY[7];
            assign M_AXIMM_7_ARADDR = dm_ARADDR[7][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_7_ARLEN = dm_ARLEN[7];
            assign M_AXIMM_7_ARSIZE = dm_ARSIZE[7];
            assign M_AXIMM_7_ARBURST = dm_ARBURST[7];
            assign M_AXIMM_7_ARLOCK = dm_ARLOCK[7];
            assign M_AXIMM_7_ARCACHE = dm_ARCACHE[7];
            assign M_AXIMM_7_ARPROT = dm_ARPROT[7];
            assign M_AXIMM_7_ARREGION = dm_ARREGION[7];
            assign M_AXIMM_7_ARQOS = dm_ARQOS[7];
            assign M_AXIMM_7_ARVALID = dm_ARVALID[7];
            assign dm_ARREADY[7] = M_AXIMM_7_ARREADY;
            assign dm_RDATA[7][M_AXIMM_7_DATA_WIDTH-1:0] = M_AXIMM_7_RDATA;
            assign dm_RRESP[7] = M_AXIMM_7_RRESP;
            assign dm_RLAST[7] = M_AXIMM_7_RLAST;
            assign dm_RVALID[7] = M_AXIMM_7_RVALID;
            assign M_AXIMM_7_RREADY = dm_RREADY[7];
        end
        if(C_NUM_AXIMMs > 8) begin
            assign ap_AWADDR[8][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_8_AWADDR;
            assign ap_AWLEN[8] = AP_AXIMM_8_AWLEN;
            assign ap_AWSIZE[8] = AP_AXIMM_8_AWSIZE;
            assign ap_AWBURST[8] = AP_AXIMM_8_AWBURST;
            assign ap_AWLOCK[8] = AP_AXIMM_8_AWLOCK;
            assign ap_AWCACHE[8] = AP_AXIMM_8_AWCACHE;
            assign ap_AWPROT[8] = AP_AXIMM_8_AWPROT;
            assign ap_AWREGION[8] = AP_AXIMM_8_AWREGION;
            assign ap_AWQOS[8] = AP_AXIMM_8_AWQOS;
            assign ap_AWVALID[8] = AP_AXIMM_8_AWVALID;
            assign AP_AXIMM_8_AWREADY = ap_AWREADY[8];
            assign ap_WDATA[8][M_AXIMM_8_DATA_WIDTH-1:0] = AP_AXIMM_8_WDATA;
            assign ap_WSTRB[8][M_AXIMM_8_DATA_WIDTH/8-1:0] = AP_AXIMM_8_WSTRB;
            assign ap_WLAST[8] = AP_AXIMM_8_WLAST;
            assign ap_WVALID[8] = AP_AXIMM_8_WVALID;
            assign AP_AXIMM_8_WREADY = ap_WREADY[8];
            assign AP_AXIMM_8_BRESP = ap_BRESP[8];
            assign AP_AXIMM_8_BVALID = ap_BVALID[8];
            assign ap_BREADY[8] = AP_AXIMM_8_BREADY;
            assign ap_ARADDR[8][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_8_ARADDR;
            assign ap_ARLEN[8] = AP_AXIMM_8_ARLEN;
            assign ap_ARSIZE[8] = AP_AXIMM_8_ARSIZE;
            assign ap_ARBURST[8] = AP_AXIMM_8_ARBURST;
            assign ap_ARLOCK[8] = AP_AXIMM_8_ARLOCK;
            assign ap_ARCACHE[8] = AP_AXIMM_8_ARCACHE;
            assign ap_ARPROT[8] = AP_AXIMM_8_ARPROT;
            assign ap_ARREGION[8] = AP_AXIMM_8_ARREGION;
            assign ap_ARQOS[8] = AP_AXIMM_8_ARQOS;
            assign ap_ARVALID[8] = AP_AXIMM_8_ARVALID;
            assign AP_AXIMM_8_ARREADY = ap_ARREADY[8];
            assign AP_AXIMM_8_RDATA = ap_RDATA[8][M_AXIMM_8_DATA_WIDTH-1:0];
            assign AP_AXIMM_8_RRESP = ap_RRESP[8];
            assign AP_AXIMM_8_RLAST = ap_RLAST[8];
            assign AP_AXIMM_8_RVALID = ap_RVALID[8];
            assign ap_RREADY[8] = AP_AXIMM_8_RREADY;
            assign M_AXIMM_8_AWADDR = dm_AWADDR[8][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_8_AWLEN = dm_AWLEN[8];
            assign M_AXIMM_8_AWSIZE = dm_AWSIZE[8];
            assign M_AXIMM_8_AWBURST = dm_AWBURST[8];
            assign M_AXIMM_8_AWLOCK = dm_AWLOCK[8];
            assign M_AXIMM_8_AWCACHE = dm_AWCACHE[8];
            assign M_AXIMM_8_AWPROT = dm_AWPROT[8];
            assign M_AXIMM_8_AWREGION = dm_AWREGION[8];
            assign M_AXIMM_8_AWQOS = dm_AWQOS[8];
            assign M_AXIMM_8_AWVALID = dm_AWVALID[8];
            assign dm_AWREADY[8] = M_AXIMM_8_AWREADY;
            assign M_AXIMM_8_WDATA = dm_WDATA[8][M_AXIMM_8_DATA_WIDTH-1:0];
            assign M_AXIMM_8_WSTRB = dm_WSTRB[8][M_AXIMM_8_DATA_WIDTH/8-1:0];
            assign M_AXIMM_8_WLAST = dm_WLAST[8];
            assign M_AXIMM_8_WVALID = dm_WVALID[8];
            assign dm_WREADY[8] = M_AXIMM_8_WREADY;
            assign dm_BRESP[8] = M_AXIMM_8_BRESP;
            assign dm_BVALID[8] = M_AXIMM_8_BVALID;
            assign M_AXIMM_8_BREADY = dm_BREADY[8];
            assign M_AXIMM_8_ARADDR = dm_ARADDR[8][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_8_ARLEN = dm_ARLEN[8];
            assign M_AXIMM_8_ARSIZE = dm_ARSIZE[8];
            assign M_AXIMM_8_ARBURST = dm_ARBURST[8];
            assign M_AXIMM_8_ARLOCK = dm_ARLOCK[8];
            assign M_AXIMM_8_ARCACHE = dm_ARCACHE[8];
            assign M_AXIMM_8_ARPROT = dm_ARPROT[8];
            assign M_AXIMM_8_ARREGION = dm_ARREGION[8];
            assign M_AXIMM_8_ARQOS = dm_ARQOS[8];
            assign M_AXIMM_8_ARVALID = dm_ARVALID[8];
            assign dm_ARREADY[8] = M_AXIMM_8_ARREADY;
            assign dm_RDATA[8][M_AXIMM_8_DATA_WIDTH-1:0] = M_AXIMM_8_RDATA;
            assign dm_RRESP[8] = M_AXIMM_8_RRESP;
            assign dm_RLAST[8] = M_AXIMM_8_RLAST;
            assign dm_RVALID[8] = M_AXIMM_8_RVALID;
            assign M_AXIMM_8_RREADY = dm_RREADY[8];
        end
        if(C_NUM_AXIMMs > 9) begin
            assign ap_AWADDR[9][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_9_AWADDR;
            assign ap_AWLEN[9] = AP_AXIMM_9_AWLEN;
            assign ap_AWSIZE[9] = AP_AXIMM_9_AWSIZE;
            assign ap_AWBURST[9] = AP_AXIMM_9_AWBURST;
            assign ap_AWLOCK[9] = AP_AXIMM_9_AWLOCK;
            assign ap_AWCACHE[9] = AP_AXIMM_9_AWCACHE;
            assign ap_AWPROT[9] = AP_AXIMM_9_AWPROT;
            assign ap_AWREGION[9] = AP_AXIMM_9_AWREGION;
            assign ap_AWQOS[9] = AP_AXIMM_9_AWQOS;
            assign ap_AWVALID[9] = AP_AXIMM_9_AWVALID;
            assign AP_AXIMM_9_AWREADY = ap_AWREADY[9];
            assign ap_WDATA[9][M_AXIMM_9_DATA_WIDTH-1:0] = AP_AXIMM_9_WDATA;
            assign ap_WSTRB[9][M_AXIMM_9_DATA_WIDTH/8-1:0] = AP_AXIMM_9_WSTRB;
            assign ap_WLAST[9] = AP_AXIMM_9_WLAST;
            assign ap_WVALID[9] = AP_AXIMM_9_WVALID;
            assign AP_AXIMM_9_WREADY = ap_WREADY[9];
            assign AP_AXIMM_9_BRESP = ap_BRESP[9];
            assign AP_AXIMM_9_BVALID = ap_BVALID[9];
            assign ap_BREADY[9] = AP_AXIMM_9_BREADY;
            assign ap_ARADDR[9][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_9_ARADDR;
            assign ap_ARLEN[9] = AP_AXIMM_9_ARLEN;
            assign ap_ARSIZE[9] = AP_AXIMM_9_ARSIZE;
            assign ap_ARBURST[9] = AP_AXIMM_9_ARBURST;
            assign ap_ARLOCK[9] = AP_AXIMM_9_ARLOCK;
            assign ap_ARCACHE[9] = AP_AXIMM_9_ARCACHE;
            assign ap_ARPROT[9] = AP_AXIMM_9_ARPROT;
            assign ap_ARREGION[9] = AP_AXIMM_9_ARREGION;
            assign ap_ARQOS[9] = AP_AXIMM_9_ARQOS;
            assign ap_ARVALID[9] = AP_AXIMM_9_ARVALID;
            assign AP_AXIMM_9_ARREADY = ap_ARREADY[9];
            assign AP_AXIMM_9_RDATA = ap_RDATA[9][M_AXIMM_9_DATA_WIDTH-1:0];
            assign AP_AXIMM_9_RRESP = ap_RRESP[9];
            assign AP_AXIMM_9_RLAST = ap_RLAST[9];
            assign AP_AXIMM_9_RVALID = ap_RVALID[9];
            assign ap_RREADY[9] = AP_AXIMM_9_RREADY;
            assign M_AXIMM_9_AWADDR = dm_AWADDR[9][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_9_AWLEN = dm_AWLEN[9];
            assign M_AXIMM_9_AWSIZE = dm_AWSIZE[9];
            assign M_AXIMM_9_AWBURST = dm_AWBURST[9];
            assign M_AXIMM_9_AWLOCK = dm_AWLOCK[9];
            assign M_AXIMM_9_AWCACHE = dm_AWCACHE[9];
            assign M_AXIMM_9_AWPROT = dm_AWPROT[9];
            assign M_AXIMM_9_AWREGION = dm_AWREGION[9];
            assign M_AXIMM_9_AWQOS = dm_AWQOS[9];
            assign M_AXIMM_9_AWVALID = dm_AWVALID[9];
            assign dm_AWREADY[9] = M_AXIMM_9_AWREADY;
            assign M_AXIMM_9_WDATA = dm_WDATA[9][M_AXIMM_9_DATA_WIDTH-1:0];
            assign M_AXIMM_9_WSTRB = dm_WSTRB[9][M_AXIMM_9_DATA_WIDTH/8-1:0];
            assign M_AXIMM_9_WLAST = dm_WLAST[9];
            assign M_AXIMM_9_WVALID = dm_WVALID[9];
            assign dm_WREADY[9] = M_AXIMM_9_WREADY;
            assign dm_BRESP[9] = M_AXIMM_9_BRESP;
            assign dm_BVALID[9] = M_AXIMM_9_BVALID;
            assign M_AXIMM_9_BREADY = dm_BREADY[9];
            assign M_AXIMM_9_ARADDR = dm_ARADDR[9][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_9_ARLEN = dm_ARLEN[9];
            assign M_AXIMM_9_ARSIZE = dm_ARSIZE[9];
            assign M_AXIMM_9_ARBURST = dm_ARBURST[9];
            assign M_AXIMM_9_ARLOCK = dm_ARLOCK[9];
            assign M_AXIMM_9_ARCACHE = dm_ARCACHE[9];
            assign M_AXIMM_9_ARPROT = dm_ARPROT[9];
            assign M_AXIMM_9_ARREGION = dm_ARREGION[9];
            assign M_AXIMM_9_ARQOS = dm_ARQOS[9];
            assign M_AXIMM_9_ARVALID = dm_ARVALID[9];
            assign dm_ARREADY[9] = M_AXIMM_9_ARREADY;
            assign dm_RDATA[9][M_AXIMM_9_DATA_WIDTH-1:0] = M_AXIMM_9_RDATA;
            assign dm_RRESP[9] = M_AXIMM_9_RRESP;
            assign dm_RLAST[9] = M_AXIMM_9_RLAST;
            assign dm_RVALID[9] = M_AXIMM_9_RVALID;
            assign M_AXIMM_9_RREADY = dm_RREADY[9];
        end
        if(C_NUM_AXIMMs > 10) begin
            assign ap_AWADDR[10][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_10_AWADDR;
            assign ap_AWLEN[10] = AP_AXIMM_10_AWLEN;
            assign ap_AWSIZE[10] = AP_AXIMM_10_AWSIZE;
            assign ap_AWBURST[10] = AP_AXIMM_10_AWBURST;
            assign ap_AWLOCK[10] = AP_AXIMM_10_AWLOCK;
            assign ap_AWCACHE[10] = AP_AXIMM_10_AWCACHE;
            assign ap_AWPROT[10] = AP_AXIMM_10_AWPROT;
            assign ap_AWREGION[10] = AP_AXIMM_10_AWREGION;
            assign ap_AWQOS[10] = AP_AXIMM_10_AWQOS;
            assign ap_AWVALID[10] = AP_AXIMM_10_AWVALID;
            assign AP_AXIMM_10_AWREADY = ap_AWREADY[10];
            assign ap_WDATA[10][M_AXIMM_10_DATA_WIDTH-1:0] = AP_AXIMM_10_WDATA;
            assign ap_WSTRB[10][M_AXIMM_10_DATA_WIDTH/8-1:0] = AP_AXIMM_10_WSTRB;
            assign ap_WLAST[10] = AP_AXIMM_10_WLAST;
            assign ap_WVALID[10] = AP_AXIMM_10_WVALID;
            assign AP_AXIMM_10_WREADY = ap_WREADY[10];
            assign AP_AXIMM_10_BRESP = ap_BRESP[10];
            assign AP_AXIMM_10_BVALID = ap_BVALID[10];
            assign ap_BREADY[10] = AP_AXIMM_10_BREADY;
            assign ap_ARADDR[10][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_10_ARADDR;
            assign ap_ARLEN[10] = AP_AXIMM_10_ARLEN;
            assign ap_ARSIZE[10] = AP_AXIMM_10_ARSIZE;
            assign ap_ARBURST[10] = AP_AXIMM_10_ARBURST;
            assign ap_ARLOCK[10] = AP_AXIMM_10_ARLOCK;
            assign ap_ARCACHE[10] = AP_AXIMM_10_ARCACHE;
            assign ap_ARPROT[10] = AP_AXIMM_10_ARPROT;
            assign ap_ARREGION[10] = AP_AXIMM_10_ARREGION;
            assign ap_ARQOS[10] = AP_AXIMM_10_ARQOS;
            assign ap_ARVALID[10] = AP_AXIMM_10_ARVALID;
            assign AP_AXIMM_10_ARREADY = ap_ARREADY[10];
            assign AP_AXIMM_10_RDATA = ap_RDATA[10][M_AXIMM_10_DATA_WIDTH-1:0];
            assign AP_AXIMM_10_RRESP = ap_RRESP[10];
            assign AP_AXIMM_10_RLAST = ap_RLAST[10];
            assign AP_AXIMM_10_RVALID = ap_RVALID[10];
            assign ap_RREADY[10] = AP_AXIMM_10_RREADY;
            assign M_AXIMM_10_AWADDR = dm_AWADDR[10][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_10_AWLEN = dm_AWLEN[10];
            assign M_AXIMM_10_AWSIZE = dm_AWSIZE[10];
            assign M_AXIMM_10_AWBURST = dm_AWBURST[10];
            assign M_AXIMM_10_AWLOCK = dm_AWLOCK[10];
            assign M_AXIMM_10_AWCACHE = dm_AWCACHE[10];
            assign M_AXIMM_10_AWPROT = dm_AWPROT[10];
            assign M_AXIMM_10_AWREGION = dm_AWREGION[10];
            assign M_AXIMM_10_AWQOS = dm_AWQOS[10];
            assign M_AXIMM_10_AWVALID = dm_AWVALID[10];
            assign dm_AWREADY[10] = M_AXIMM_10_AWREADY;
            assign M_AXIMM_10_WDATA = dm_WDATA[10][M_AXIMM_10_DATA_WIDTH-1:0];
            assign M_AXIMM_10_WSTRB = dm_WSTRB[10][M_AXIMM_10_DATA_WIDTH/8-1:0];
            assign M_AXIMM_10_WLAST = dm_WLAST[10];
            assign M_AXIMM_10_WVALID = dm_WVALID[10];
            assign dm_WREADY[10] = M_AXIMM_10_WREADY;
            assign dm_BRESP[10] = M_AXIMM_10_BRESP;
            assign dm_BVALID[10] = M_AXIMM_10_BVALID;
            assign M_AXIMM_10_BREADY = dm_BREADY[10];
            assign M_AXIMM_10_ARADDR = dm_ARADDR[10][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_10_ARLEN = dm_ARLEN[10];
            assign M_AXIMM_10_ARSIZE = dm_ARSIZE[10];
            assign M_AXIMM_10_ARBURST = dm_ARBURST[10];
            assign M_AXIMM_10_ARLOCK = dm_ARLOCK[10];
            assign M_AXIMM_10_ARCACHE = dm_ARCACHE[10];
            assign M_AXIMM_10_ARPROT = dm_ARPROT[10];
            assign M_AXIMM_10_ARREGION = dm_ARREGION[10];
            assign M_AXIMM_10_ARQOS = dm_ARQOS[10];
            assign M_AXIMM_10_ARVALID = dm_ARVALID[10];
            assign dm_ARREADY[10] = M_AXIMM_10_ARREADY;
            assign dm_RDATA[10][M_AXIMM_10_DATA_WIDTH-1:0] = M_AXIMM_10_RDATA;
            assign dm_RRESP[10] = M_AXIMM_10_RRESP;
            assign dm_RLAST[10] = M_AXIMM_10_RLAST;
            assign dm_RVALID[10] = M_AXIMM_10_RVALID;
            assign M_AXIMM_10_RREADY = dm_RREADY[10];
        end
        if(C_NUM_AXIMMs > 11) begin
            assign ap_AWADDR[11][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_11_AWADDR;
            assign ap_AWLEN[11] = AP_AXIMM_11_AWLEN;
            assign ap_AWSIZE[11] = AP_AXIMM_11_AWSIZE;
            assign ap_AWBURST[11] = AP_AXIMM_11_AWBURST;
            assign ap_AWLOCK[11] = AP_AXIMM_11_AWLOCK;
            assign ap_AWCACHE[11] = AP_AXIMM_11_AWCACHE;
            assign ap_AWPROT[11] = AP_AXIMM_11_AWPROT;
            assign ap_AWREGION[11] = AP_AXIMM_11_AWREGION;
            assign ap_AWQOS[11] = AP_AXIMM_11_AWQOS;
            assign ap_AWVALID[11] = AP_AXIMM_11_AWVALID;
            assign AP_AXIMM_11_AWREADY = ap_AWREADY[11];
            assign ap_WDATA[11][M_AXIMM_11_DATA_WIDTH-1:0] = AP_AXIMM_11_WDATA;
            assign ap_WSTRB[11][M_AXIMM_11_DATA_WIDTH/8-1:0] = AP_AXIMM_11_WSTRB;
            assign ap_WLAST[11] = AP_AXIMM_11_WLAST;
            assign ap_WVALID[11] = AP_AXIMM_11_WVALID;
            assign AP_AXIMM_11_WREADY = ap_WREADY[11];
            assign AP_AXIMM_11_BRESP = ap_BRESP[11];
            assign AP_AXIMM_11_BVALID = ap_BVALID[11];
            assign ap_BREADY[11] = AP_AXIMM_11_BREADY;
            assign ap_ARADDR[11][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_11_ARADDR;
            assign ap_ARLEN[11] = AP_AXIMM_11_ARLEN;
            assign ap_ARSIZE[11] = AP_AXIMM_11_ARSIZE;
            assign ap_ARBURST[11] = AP_AXIMM_11_ARBURST;
            assign ap_ARLOCK[11] = AP_AXIMM_11_ARLOCK;
            assign ap_ARCACHE[11] = AP_AXIMM_11_ARCACHE;
            assign ap_ARPROT[11] = AP_AXIMM_11_ARPROT;
            assign ap_ARREGION[11] = AP_AXIMM_11_ARREGION;
            assign ap_ARQOS[11] = AP_AXIMM_11_ARQOS;
            assign ap_ARVALID[11] = AP_AXIMM_11_ARVALID;
            assign AP_AXIMM_11_ARREADY = ap_ARREADY[11];
            assign AP_AXIMM_11_RDATA = ap_RDATA[11][M_AXIMM_11_DATA_WIDTH-1:0];
            assign AP_AXIMM_11_RRESP = ap_RRESP[11];
            assign AP_AXIMM_11_RLAST = ap_RLAST[11];
            assign AP_AXIMM_11_RVALID = ap_RVALID[11];
            assign ap_RREADY[11] = AP_AXIMM_11_RREADY;
            assign M_AXIMM_11_AWADDR = dm_AWADDR[11][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_11_AWLEN = dm_AWLEN[11];
            assign M_AXIMM_11_AWSIZE = dm_AWSIZE[11];
            assign M_AXIMM_11_AWBURST = dm_AWBURST[11];
            assign M_AXIMM_11_AWLOCK = dm_AWLOCK[11];
            assign M_AXIMM_11_AWCACHE = dm_AWCACHE[11];
            assign M_AXIMM_11_AWPROT = dm_AWPROT[11];
            assign M_AXIMM_11_AWREGION = dm_AWREGION[11];
            assign M_AXIMM_11_AWQOS = dm_AWQOS[11];
            assign M_AXIMM_11_AWVALID = dm_AWVALID[11];
            assign dm_AWREADY[11] = M_AXIMM_11_AWREADY;
            assign M_AXIMM_11_WDATA = dm_WDATA[11][M_AXIMM_11_DATA_WIDTH-1:0];
            assign M_AXIMM_11_WSTRB = dm_WSTRB[11][M_AXIMM_11_DATA_WIDTH/8-1:0];
            assign M_AXIMM_11_WLAST = dm_WLAST[11];
            assign M_AXIMM_11_WVALID = dm_WVALID[11];
            assign dm_WREADY[11] = M_AXIMM_11_WREADY;
            assign dm_BRESP[11] = M_AXIMM_11_BRESP;
            assign dm_BVALID[11] = M_AXIMM_11_BVALID;
            assign M_AXIMM_11_BREADY = dm_BREADY[11];
            assign M_AXIMM_11_ARADDR = dm_ARADDR[11][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_11_ARLEN = dm_ARLEN[11];
            assign M_AXIMM_11_ARSIZE = dm_ARSIZE[11];
            assign M_AXIMM_11_ARBURST = dm_ARBURST[11];
            assign M_AXIMM_11_ARLOCK = dm_ARLOCK[11];
            assign M_AXIMM_11_ARCACHE = dm_ARCACHE[11];
            assign M_AXIMM_11_ARPROT = dm_ARPROT[11];
            assign M_AXIMM_11_ARREGION = dm_ARREGION[11];
            assign M_AXIMM_11_ARQOS = dm_ARQOS[11];
            assign M_AXIMM_11_ARVALID = dm_ARVALID[11];
            assign dm_ARREADY[11] = M_AXIMM_11_ARREADY;
            assign dm_RDATA[11][M_AXIMM_11_DATA_WIDTH-1:0] = M_AXIMM_11_RDATA;
            assign dm_RRESP[11] = M_AXIMM_11_RRESP;
            assign dm_RLAST[11] = M_AXIMM_11_RLAST;
            assign dm_RVALID[11] = M_AXIMM_11_RVALID;
            assign M_AXIMM_11_RREADY = dm_RREADY[11];
        end
        if(C_NUM_AXIMMs > 12) begin
            assign ap_AWADDR[12][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_12_AWADDR;
            assign ap_AWLEN[12] = AP_AXIMM_12_AWLEN;
            assign ap_AWSIZE[12] = AP_AXIMM_12_AWSIZE;
            assign ap_AWBURST[12] = AP_AXIMM_12_AWBURST;
            assign ap_AWLOCK[12] = AP_AXIMM_12_AWLOCK;
            assign ap_AWCACHE[12] = AP_AXIMM_12_AWCACHE;
            assign ap_AWPROT[12] = AP_AXIMM_12_AWPROT;
            assign ap_AWREGION[12] = AP_AXIMM_12_AWREGION;
            assign ap_AWQOS[12] = AP_AXIMM_12_AWQOS;
            assign ap_AWVALID[12] = AP_AXIMM_12_AWVALID;
            assign AP_AXIMM_12_AWREADY = ap_AWREADY[12];
            assign ap_WDATA[12][M_AXIMM_12_DATA_WIDTH-1:0] = AP_AXIMM_12_WDATA;
            assign ap_WSTRB[12][M_AXIMM_12_DATA_WIDTH/8-1:0] = AP_AXIMM_12_WSTRB;
            assign ap_WLAST[12] = AP_AXIMM_12_WLAST;
            assign ap_WVALID[12] = AP_AXIMM_12_WVALID;
            assign AP_AXIMM_12_WREADY = ap_WREADY[12];
            assign AP_AXIMM_12_BRESP = ap_BRESP[12];
            assign AP_AXIMM_12_BVALID = ap_BVALID[12];
            assign ap_BREADY[12] = AP_AXIMM_12_BREADY;
            assign ap_ARADDR[12][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_12_ARADDR;
            assign ap_ARLEN[12] = AP_AXIMM_12_ARLEN;
            assign ap_ARSIZE[12] = AP_AXIMM_12_ARSIZE;
            assign ap_ARBURST[12] = AP_AXIMM_12_ARBURST;
            assign ap_ARLOCK[12] = AP_AXIMM_12_ARLOCK;
            assign ap_ARCACHE[12] = AP_AXIMM_12_ARCACHE;
            assign ap_ARPROT[12] = AP_AXIMM_12_ARPROT;
            assign ap_ARREGION[12] = AP_AXIMM_12_ARREGION;
            assign ap_ARQOS[12] = AP_AXIMM_12_ARQOS;
            assign ap_ARVALID[12] = AP_AXIMM_12_ARVALID;
            assign AP_AXIMM_12_ARREADY = ap_ARREADY[12];
            assign AP_AXIMM_12_RDATA = ap_RDATA[12][M_AXIMM_12_DATA_WIDTH-1:0];
            assign AP_AXIMM_12_RRESP = ap_RRESP[12];
            assign AP_AXIMM_12_RLAST = ap_RLAST[12];
            assign AP_AXIMM_12_RVALID = ap_RVALID[12];
            assign ap_RREADY[12] = AP_AXIMM_12_RREADY;
            assign M_AXIMM_12_AWADDR = dm_AWADDR[12][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_12_AWLEN = dm_AWLEN[12];
            assign M_AXIMM_12_AWSIZE = dm_AWSIZE[12];
            assign M_AXIMM_12_AWBURST = dm_AWBURST[12];
            assign M_AXIMM_12_AWLOCK = dm_AWLOCK[12];
            assign M_AXIMM_12_AWCACHE = dm_AWCACHE[12];
            assign M_AXIMM_12_AWPROT = dm_AWPROT[12];
            assign M_AXIMM_12_AWREGION = dm_AWREGION[12];
            assign M_AXIMM_12_AWQOS = dm_AWQOS[12];
            assign M_AXIMM_12_AWVALID = dm_AWVALID[12];
            assign dm_AWREADY[12] = M_AXIMM_12_AWREADY;
            assign M_AXIMM_12_WDATA = dm_WDATA[12][M_AXIMM_12_DATA_WIDTH-1:0];
            assign M_AXIMM_12_WSTRB = dm_WSTRB[12][M_AXIMM_12_DATA_WIDTH/8-1:0];
            assign M_AXIMM_12_WLAST = dm_WLAST[12];
            assign M_AXIMM_12_WVALID = dm_WVALID[12];
            assign dm_WREADY[12] = M_AXIMM_12_WREADY;
            assign dm_BRESP[12] = M_AXIMM_12_BRESP;
            assign dm_BVALID[12] = M_AXIMM_12_BVALID;
            assign M_AXIMM_12_BREADY = dm_BREADY[12];
            assign M_AXIMM_12_ARADDR = dm_ARADDR[12][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_12_ARLEN = dm_ARLEN[12];
            assign M_AXIMM_12_ARSIZE = dm_ARSIZE[12];
            assign M_AXIMM_12_ARBURST = dm_ARBURST[12];
            assign M_AXIMM_12_ARLOCK = dm_ARLOCK[12];
            assign M_AXIMM_12_ARCACHE = dm_ARCACHE[12];
            assign M_AXIMM_12_ARPROT = dm_ARPROT[12];
            assign M_AXIMM_12_ARREGION = dm_ARREGION[12];
            assign M_AXIMM_12_ARQOS = dm_ARQOS[12];
            assign M_AXIMM_12_ARVALID = dm_ARVALID[12];
            assign dm_ARREADY[12] = M_AXIMM_12_ARREADY;
            assign dm_RDATA[12][M_AXIMM_12_DATA_WIDTH-1:0] = M_AXIMM_12_RDATA;
            assign dm_RRESP[12] = M_AXIMM_12_RRESP;
            assign dm_RLAST[12] = M_AXIMM_12_RLAST;
            assign dm_RVALID[12] = M_AXIMM_12_RVALID;
            assign M_AXIMM_12_RREADY = dm_RREADY[12];
        end
        if(C_NUM_AXIMMs > 13) begin
            assign ap_AWADDR[13][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_13_AWADDR;
            assign ap_AWLEN[13] = AP_AXIMM_13_AWLEN;
            assign ap_AWSIZE[13] = AP_AXIMM_13_AWSIZE;
            assign ap_AWBURST[13] = AP_AXIMM_13_AWBURST;
            assign ap_AWLOCK[13] = AP_AXIMM_13_AWLOCK;
            assign ap_AWCACHE[13] = AP_AXIMM_13_AWCACHE;
            assign ap_AWPROT[13] = AP_AXIMM_13_AWPROT;
            assign ap_AWREGION[13] = AP_AXIMM_13_AWREGION;
            assign ap_AWQOS[13] = AP_AXIMM_13_AWQOS;
            assign ap_AWVALID[13] = AP_AXIMM_13_AWVALID;
            assign AP_AXIMM_13_AWREADY = ap_AWREADY[13];
            assign ap_WDATA[13][M_AXIMM_13_DATA_WIDTH-1:0] = AP_AXIMM_13_WDATA;
            assign ap_WSTRB[13][M_AXIMM_13_DATA_WIDTH/8-1:0] = AP_AXIMM_13_WSTRB;
            assign ap_WLAST[13] = AP_AXIMM_13_WLAST;
            assign ap_WVALID[13] = AP_AXIMM_13_WVALID;
            assign AP_AXIMM_13_WREADY = ap_WREADY[13];
            assign AP_AXIMM_13_BRESP = ap_BRESP[13];
            assign AP_AXIMM_13_BVALID = ap_BVALID[13];
            assign ap_BREADY[13] = AP_AXIMM_13_BREADY;
            assign ap_ARADDR[13][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_13_ARADDR;
            assign ap_ARLEN[13] = AP_AXIMM_13_ARLEN;
            assign ap_ARSIZE[13] = AP_AXIMM_13_ARSIZE;
            assign ap_ARBURST[13] = AP_AXIMM_13_ARBURST;
            assign ap_ARLOCK[13] = AP_AXIMM_13_ARLOCK;
            assign ap_ARCACHE[13] = AP_AXIMM_13_ARCACHE;
            assign ap_ARPROT[13] = AP_AXIMM_13_ARPROT;
            assign ap_ARREGION[13] = AP_AXIMM_13_ARREGION;
            assign ap_ARQOS[13] = AP_AXIMM_13_ARQOS;
            assign ap_ARVALID[13] = AP_AXIMM_13_ARVALID;
            assign AP_AXIMM_13_ARREADY = ap_ARREADY[13];
            assign AP_AXIMM_13_RDATA = ap_RDATA[13][M_AXIMM_13_DATA_WIDTH-1:0];
            assign AP_AXIMM_13_RRESP = ap_RRESP[13];
            assign AP_AXIMM_13_RLAST = ap_RLAST[13];
            assign AP_AXIMM_13_RVALID = ap_RVALID[13];
            assign ap_RREADY[13] = AP_AXIMM_13_RREADY;
            assign M_AXIMM_13_AWADDR = dm_AWADDR[13][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_13_AWLEN = dm_AWLEN[13];
            assign M_AXIMM_13_AWSIZE = dm_AWSIZE[13];
            assign M_AXIMM_13_AWBURST = dm_AWBURST[13];
            assign M_AXIMM_13_AWLOCK = dm_AWLOCK[13];
            assign M_AXIMM_13_AWCACHE = dm_AWCACHE[13];
            assign M_AXIMM_13_AWPROT = dm_AWPROT[13];
            assign M_AXIMM_13_AWREGION = dm_AWREGION[13];
            assign M_AXIMM_13_AWQOS = dm_AWQOS[13];
            assign M_AXIMM_13_AWVALID = dm_AWVALID[13];
            assign dm_AWREADY[13] = M_AXIMM_13_AWREADY;
            assign M_AXIMM_13_WDATA = dm_WDATA[13][M_AXIMM_13_DATA_WIDTH-1:0];
            assign M_AXIMM_13_WSTRB = dm_WSTRB[13][M_AXIMM_13_DATA_WIDTH/8-1:0];
            assign M_AXIMM_13_WLAST = dm_WLAST[13];
            assign M_AXIMM_13_WVALID = dm_WVALID[13];
            assign dm_WREADY[13] = M_AXIMM_13_WREADY;
            assign dm_BRESP[13] = M_AXIMM_13_BRESP;
            assign dm_BVALID[13] = M_AXIMM_13_BVALID;
            assign M_AXIMM_13_BREADY = dm_BREADY[13];
            assign M_AXIMM_13_ARADDR = dm_ARADDR[13][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_13_ARLEN = dm_ARLEN[13];
            assign M_AXIMM_13_ARSIZE = dm_ARSIZE[13];
            assign M_AXIMM_13_ARBURST = dm_ARBURST[13];
            assign M_AXIMM_13_ARLOCK = dm_ARLOCK[13];
            assign M_AXIMM_13_ARCACHE = dm_ARCACHE[13];
            assign M_AXIMM_13_ARPROT = dm_ARPROT[13];
            assign M_AXIMM_13_ARREGION = dm_ARREGION[13];
            assign M_AXIMM_13_ARQOS = dm_ARQOS[13];
            assign M_AXIMM_13_ARVALID = dm_ARVALID[13];
            assign dm_ARREADY[13] = M_AXIMM_13_ARREADY;
            assign dm_RDATA[13][M_AXIMM_13_DATA_WIDTH-1:0] = M_AXIMM_13_RDATA;
            assign dm_RRESP[13] = M_AXIMM_13_RRESP;
            assign dm_RLAST[13] = M_AXIMM_13_RLAST;
            assign dm_RVALID[13] = M_AXIMM_13_RVALID;
            assign M_AXIMM_13_RREADY = dm_RREADY[13];
        end
        if(C_NUM_AXIMMs > 14) begin
            assign ap_AWADDR[14][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_14_AWADDR;
            assign ap_AWLEN[14] = AP_AXIMM_14_AWLEN;
            assign ap_AWSIZE[14] = AP_AXIMM_14_AWSIZE;
            assign ap_AWBURST[14] = AP_AXIMM_14_AWBURST;
            assign ap_AWLOCK[14] = AP_AXIMM_14_AWLOCK;
            assign ap_AWCACHE[14] = AP_AXIMM_14_AWCACHE;
            assign ap_AWPROT[14] = AP_AXIMM_14_AWPROT;
            assign ap_AWREGION[14] = AP_AXIMM_14_AWREGION;
            assign ap_AWQOS[14] = AP_AXIMM_14_AWQOS;
            assign ap_AWVALID[14] = AP_AXIMM_14_AWVALID;
            assign AP_AXIMM_14_AWREADY = ap_AWREADY[14];
            assign ap_WDATA[14][M_AXIMM_14_DATA_WIDTH-1:0] = AP_AXIMM_14_WDATA;
            assign ap_WSTRB[14][M_AXIMM_14_DATA_WIDTH/8-1:0] = AP_AXIMM_14_WSTRB;
            assign ap_WLAST[14] = AP_AXIMM_14_WLAST;
            assign ap_WVALID[14] = AP_AXIMM_14_WVALID;
            assign AP_AXIMM_14_WREADY = ap_WREADY[14];
            assign AP_AXIMM_14_BRESP = ap_BRESP[14];
            assign AP_AXIMM_14_BVALID = ap_BVALID[14];
            assign ap_BREADY[14] = AP_AXIMM_14_BREADY;
            assign ap_ARADDR[14][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_14_ARADDR;
            assign ap_ARLEN[14] = AP_AXIMM_14_ARLEN;
            assign ap_ARSIZE[14] = AP_AXIMM_14_ARSIZE;
            assign ap_ARBURST[14] = AP_AXIMM_14_ARBURST;
            assign ap_ARLOCK[14] = AP_AXIMM_14_ARLOCK;
            assign ap_ARCACHE[14] = AP_AXIMM_14_ARCACHE;
            assign ap_ARPROT[14] = AP_AXIMM_14_ARPROT;
            assign ap_ARREGION[14] = AP_AXIMM_14_ARREGION;
            assign ap_ARQOS[14] = AP_AXIMM_14_ARQOS;
            assign ap_ARVALID[14] = AP_AXIMM_14_ARVALID;
            assign AP_AXIMM_14_ARREADY = ap_ARREADY[14];
            assign AP_AXIMM_14_RDATA = ap_RDATA[14][M_AXIMM_14_DATA_WIDTH-1:0];
            assign AP_AXIMM_14_RRESP = ap_RRESP[14];
            assign AP_AXIMM_14_RLAST = ap_RLAST[14];
            assign AP_AXIMM_14_RVALID = ap_RVALID[14];
            assign ap_RREADY[14] = AP_AXIMM_14_RREADY;
            assign M_AXIMM_14_AWADDR = dm_AWADDR[14][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_14_AWLEN = dm_AWLEN[14];
            assign M_AXIMM_14_AWSIZE = dm_AWSIZE[14];
            assign M_AXIMM_14_AWBURST = dm_AWBURST[14];
            assign M_AXIMM_14_AWLOCK = dm_AWLOCK[14];
            assign M_AXIMM_14_AWCACHE = dm_AWCACHE[14];
            assign M_AXIMM_14_AWPROT = dm_AWPROT[14];
            assign M_AXIMM_14_AWREGION = dm_AWREGION[14];
            assign M_AXIMM_14_AWQOS = dm_AWQOS[14];
            assign M_AXIMM_14_AWVALID = dm_AWVALID[14];
            assign dm_AWREADY[14] = M_AXIMM_14_AWREADY;
            assign M_AXIMM_14_WDATA = dm_WDATA[14][M_AXIMM_14_DATA_WIDTH-1:0];
            assign M_AXIMM_14_WSTRB = dm_WSTRB[14][M_AXIMM_14_DATA_WIDTH/8-1:0];
            assign M_AXIMM_14_WLAST = dm_WLAST[14];
            assign M_AXIMM_14_WVALID = dm_WVALID[14];
            assign dm_WREADY[14] = M_AXIMM_14_WREADY;
            assign dm_BRESP[14] = M_AXIMM_14_BRESP;
            assign dm_BVALID[14] = M_AXIMM_14_BVALID;
            assign M_AXIMM_14_BREADY = dm_BREADY[14];
            assign M_AXIMM_14_ARADDR = dm_ARADDR[14][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_14_ARLEN = dm_ARLEN[14];
            assign M_AXIMM_14_ARSIZE = dm_ARSIZE[14];
            assign M_AXIMM_14_ARBURST = dm_ARBURST[14];
            assign M_AXIMM_14_ARLOCK = dm_ARLOCK[14];
            assign M_AXIMM_14_ARCACHE = dm_ARCACHE[14];
            assign M_AXIMM_14_ARPROT = dm_ARPROT[14];
            assign M_AXIMM_14_ARREGION = dm_ARREGION[14];
            assign M_AXIMM_14_ARQOS = dm_ARQOS[14];
            assign M_AXIMM_14_ARVALID = dm_ARVALID[14];
            assign dm_ARREADY[14] = M_AXIMM_14_ARREADY;
            assign dm_RDATA[14][M_AXIMM_14_DATA_WIDTH-1:0] = M_AXIMM_14_RDATA;
            assign dm_RRESP[14] = M_AXIMM_14_RRESP;
            assign dm_RLAST[14] = M_AXIMM_14_RLAST;
            assign dm_RVALID[14] = M_AXIMM_14_RVALID;
            assign M_AXIMM_14_RREADY = dm_RREADY[14];
        end
        if(C_NUM_AXIMMs > 15) begin
            assign ap_AWADDR[15][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_15_AWADDR;
            assign ap_AWLEN[15] = AP_AXIMM_15_AWLEN;
            assign ap_AWSIZE[15] = AP_AXIMM_15_AWSIZE;
            assign ap_AWBURST[15] = AP_AXIMM_15_AWBURST;
            assign ap_AWLOCK[15] = AP_AXIMM_15_AWLOCK;
            assign ap_AWCACHE[15] = AP_AXIMM_15_AWCACHE;
            assign ap_AWPROT[15] = AP_AXIMM_15_AWPROT;
            assign ap_AWREGION[15] = AP_AXIMM_15_AWREGION;
            assign ap_AWQOS[15] = AP_AXIMM_15_AWQOS;
            assign ap_AWVALID[15] = AP_AXIMM_15_AWVALID;
            assign AP_AXIMM_15_AWREADY = ap_AWREADY[15];
            assign ap_WDATA[15][M_AXIMM_15_DATA_WIDTH-1:0] = AP_AXIMM_15_WDATA;
            assign ap_WSTRB[15][M_AXIMM_15_DATA_WIDTH/8-1:0] = AP_AXIMM_15_WSTRB;
            assign ap_WLAST[15] = AP_AXIMM_15_WLAST;
            assign ap_WVALID[15] = AP_AXIMM_15_WVALID;
            assign AP_AXIMM_15_WREADY = ap_WREADY[15];
            assign AP_AXIMM_15_BRESP = ap_BRESP[15];
            assign AP_AXIMM_15_BVALID = ap_BVALID[15];
            assign ap_BREADY[15] = AP_AXIMM_15_BREADY;
            assign ap_ARADDR[15][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_15_ARADDR;
            assign ap_ARLEN[15] = AP_AXIMM_15_ARLEN;
            assign ap_ARSIZE[15] = AP_AXIMM_15_ARSIZE;
            assign ap_ARBURST[15] = AP_AXIMM_15_ARBURST;
            assign ap_ARLOCK[15] = AP_AXIMM_15_ARLOCK;
            assign ap_ARCACHE[15] = AP_AXIMM_15_ARCACHE;
            assign ap_ARPROT[15] = AP_AXIMM_15_ARPROT;
            assign ap_ARREGION[15] = AP_AXIMM_15_ARREGION;
            assign ap_ARQOS[15] = AP_AXIMM_15_ARQOS;
            assign ap_ARVALID[15] = AP_AXIMM_15_ARVALID;
            assign AP_AXIMM_15_ARREADY = ap_ARREADY[15];
            assign AP_AXIMM_15_RDATA = ap_RDATA[15][M_AXIMM_15_DATA_WIDTH-1:0];
            assign AP_AXIMM_15_RRESP = ap_RRESP[15];
            assign AP_AXIMM_15_RLAST = ap_RLAST[15];
            assign AP_AXIMM_15_RVALID = ap_RVALID[15];
            assign ap_RREADY[15] = AP_AXIMM_15_RREADY;
            assign M_AXIMM_15_AWADDR = dm_AWADDR[15][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_15_AWLEN = dm_AWLEN[15];
            assign M_AXIMM_15_AWSIZE = dm_AWSIZE[15];
            assign M_AXIMM_15_AWBURST = dm_AWBURST[15];
            assign M_AXIMM_15_AWLOCK = dm_AWLOCK[15];
            assign M_AXIMM_15_AWCACHE = dm_AWCACHE[15];
            assign M_AXIMM_15_AWPROT = dm_AWPROT[15];
            assign M_AXIMM_15_AWREGION = dm_AWREGION[15];
            assign M_AXIMM_15_AWQOS = dm_AWQOS[15];
            assign M_AXIMM_15_AWVALID = dm_AWVALID[15];
            assign dm_AWREADY[15] = M_AXIMM_15_AWREADY;
            assign M_AXIMM_15_WDATA = dm_WDATA[15][M_AXIMM_15_DATA_WIDTH-1:0];
            assign M_AXIMM_15_WSTRB = dm_WSTRB[15][M_AXIMM_15_DATA_WIDTH/8-1:0];
            assign M_AXIMM_15_WLAST = dm_WLAST[15];
            assign M_AXIMM_15_WVALID = dm_WVALID[15];
            assign dm_WREADY[15] = M_AXIMM_15_WREADY;
            assign dm_BRESP[15] = M_AXIMM_15_BRESP;
            assign dm_BVALID[15] = M_AXIMM_15_BVALID;
            assign M_AXIMM_15_BREADY = dm_BREADY[15];
            assign M_AXIMM_15_ARADDR = dm_ARADDR[15][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_15_ARLEN = dm_ARLEN[15];
            assign M_AXIMM_15_ARSIZE = dm_ARSIZE[15];
            assign M_AXIMM_15_ARBURST = dm_ARBURST[15];
            assign M_AXIMM_15_ARLOCK = dm_ARLOCK[15];
            assign M_AXIMM_15_ARCACHE = dm_ARCACHE[15];
            assign M_AXIMM_15_ARPROT = dm_ARPROT[15];
            assign M_AXIMM_15_ARREGION = dm_ARREGION[15];
            assign M_AXIMM_15_ARQOS = dm_ARQOS[15];
            assign M_AXIMM_15_ARVALID = dm_ARVALID[15];
            assign dm_ARREADY[15] = M_AXIMM_15_ARREADY;
            assign dm_RDATA[15][M_AXIMM_15_DATA_WIDTH-1:0] = M_AXIMM_15_RDATA;
            assign dm_RRESP[15] = M_AXIMM_15_RRESP;
            assign dm_RLAST[15] = M_AXIMM_15_RLAST;
            assign dm_RVALID[15] = M_AXIMM_15_RVALID;
            assign M_AXIMM_15_RREADY = dm_RREADY[15];
        end
        if(C_NUM_AXIMMs > 16) begin
            assign ap_AWADDR[16][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_16_AWADDR;
            assign ap_AWLEN[16] = AP_AXIMM_16_AWLEN;
            assign ap_AWSIZE[16] = AP_AXIMM_16_AWSIZE;
            assign ap_AWBURST[16] = AP_AXIMM_16_AWBURST;
            assign ap_AWLOCK[16] = AP_AXIMM_16_AWLOCK;
            assign ap_AWCACHE[16] = AP_AXIMM_16_AWCACHE;
            assign ap_AWPROT[16] = AP_AXIMM_16_AWPROT;
            assign ap_AWREGION[16] = AP_AXIMM_16_AWREGION;
            assign ap_AWQOS[16] = AP_AXIMM_16_AWQOS;
            assign ap_AWVALID[16] = AP_AXIMM_16_AWVALID;
            assign AP_AXIMM_16_AWREADY = ap_AWREADY[16];
            assign ap_WDATA[16][M_AXIMM_16_DATA_WIDTH-1:0] = AP_AXIMM_16_WDATA;
            assign ap_WSTRB[16][M_AXIMM_16_DATA_WIDTH/8-1:0] = AP_AXIMM_16_WSTRB;
            assign ap_WLAST[16] = AP_AXIMM_16_WLAST;
            assign ap_WVALID[16] = AP_AXIMM_16_WVALID;
            assign AP_AXIMM_16_WREADY = ap_WREADY[16];
            assign AP_AXIMM_16_BRESP = ap_BRESP[16];
            assign AP_AXIMM_16_BVALID = ap_BVALID[16];
            assign ap_BREADY[16] = AP_AXIMM_16_BREADY;
            assign ap_ARADDR[16][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_16_ARADDR;
            assign ap_ARLEN[16] = AP_AXIMM_16_ARLEN;
            assign ap_ARSIZE[16] = AP_AXIMM_16_ARSIZE;
            assign ap_ARBURST[16] = AP_AXIMM_16_ARBURST;
            assign ap_ARLOCK[16] = AP_AXIMM_16_ARLOCK;
            assign ap_ARCACHE[16] = AP_AXIMM_16_ARCACHE;
            assign ap_ARPROT[16] = AP_AXIMM_16_ARPROT;
            assign ap_ARREGION[16] = AP_AXIMM_16_ARREGION;
            assign ap_ARQOS[16] = AP_AXIMM_16_ARQOS;
            assign ap_ARVALID[16] = AP_AXIMM_16_ARVALID;
            assign AP_AXIMM_16_ARREADY = ap_ARREADY[16];
            assign AP_AXIMM_16_RDATA = ap_RDATA[16][M_AXIMM_16_DATA_WIDTH-1:0];
            assign AP_AXIMM_16_RRESP = ap_RRESP[16];
            assign AP_AXIMM_16_RLAST = ap_RLAST[16];
            assign AP_AXIMM_16_RVALID = ap_RVALID[16];
            assign ap_RREADY[16] = AP_AXIMM_16_RREADY;
            assign M_AXIMM_16_AWADDR = dm_AWADDR[16][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_16_AWLEN = dm_AWLEN[16];
            assign M_AXIMM_16_AWSIZE = dm_AWSIZE[16];
            assign M_AXIMM_16_AWBURST = dm_AWBURST[16];
            assign M_AXIMM_16_AWLOCK = dm_AWLOCK[16];
            assign M_AXIMM_16_AWCACHE = dm_AWCACHE[16];
            assign M_AXIMM_16_AWPROT = dm_AWPROT[16];
            assign M_AXIMM_16_AWREGION = dm_AWREGION[16];
            assign M_AXIMM_16_AWQOS = dm_AWQOS[16];
            assign M_AXIMM_16_AWVALID = dm_AWVALID[16];
            assign dm_AWREADY[16] = M_AXIMM_16_AWREADY;
            assign M_AXIMM_16_WDATA = dm_WDATA[16][M_AXIMM_16_DATA_WIDTH-1:0];
            assign M_AXIMM_16_WSTRB = dm_WSTRB[16][M_AXIMM_16_DATA_WIDTH/8-1:0];
            assign M_AXIMM_16_WLAST = dm_WLAST[16];
            assign M_AXIMM_16_WVALID = dm_WVALID[16];
            assign dm_WREADY[16] = M_AXIMM_16_WREADY;
            assign dm_BRESP[16] = M_AXIMM_16_BRESP;
            assign dm_BVALID[16] = M_AXIMM_16_BVALID;
            assign M_AXIMM_16_BREADY = dm_BREADY[16];
            assign M_AXIMM_16_ARADDR = dm_ARADDR[16][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_16_ARLEN = dm_ARLEN[16];
            assign M_AXIMM_16_ARSIZE = dm_ARSIZE[16];
            assign M_AXIMM_16_ARBURST = dm_ARBURST[16];
            assign M_AXIMM_16_ARLOCK = dm_ARLOCK[16];
            assign M_AXIMM_16_ARCACHE = dm_ARCACHE[16];
            assign M_AXIMM_16_ARPROT = dm_ARPROT[16];
            assign M_AXIMM_16_ARREGION = dm_ARREGION[16];
            assign M_AXIMM_16_ARQOS = dm_ARQOS[16];
            assign M_AXIMM_16_ARVALID = dm_ARVALID[16];
            assign dm_ARREADY[16] = M_AXIMM_16_ARREADY;
            assign dm_RDATA[16][M_AXIMM_16_DATA_WIDTH-1:0] = M_AXIMM_16_RDATA;
            assign dm_RRESP[16] = M_AXIMM_16_RRESP;
            assign dm_RLAST[16] = M_AXIMM_16_RLAST;
            assign dm_RVALID[16] = M_AXIMM_16_RVALID;
            assign M_AXIMM_16_RREADY = dm_RREADY[16];
        end
        if(C_NUM_AXIMMs > 17) begin
            assign ap_AWADDR[17][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_17_AWADDR;
            assign ap_AWLEN[17] = AP_AXIMM_17_AWLEN;
            assign ap_AWSIZE[17] = AP_AXIMM_17_AWSIZE;
            assign ap_AWBURST[17] = AP_AXIMM_17_AWBURST;
            assign ap_AWLOCK[17] = AP_AXIMM_17_AWLOCK;
            assign ap_AWCACHE[17] = AP_AXIMM_17_AWCACHE;
            assign ap_AWPROT[17] = AP_AXIMM_17_AWPROT;
            assign ap_AWREGION[17] = AP_AXIMM_17_AWREGION;
            assign ap_AWQOS[17] = AP_AXIMM_17_AWQOS;
            assign ap_AWVALID[17] = AP_AXIMM_17_AWVALID;
            assign AP_AXIMM_17_AWREADY = ap_AWREADY[17];
            assign ap_WDATA[17][M_AXIMM_17_DATA_WIDTH-1:0] = AP_AXIMM_17_WDATA;
            assign ap_WSTRB[17][M_AXIMM_17_DATA_WIDTH/8-1:0] = AP_AXIMM_17_WSTRB;
            assign ap_WLAST[17] = AP_AXIMM_17_WLAST;
            assign ap_WVALID[17] = AP_AXIMM_17_WVALID;
            assign AP_AXIMM_17_WREADY = ap_WREADY[17];
            assign AP_AXIMM_17_BRESP = ap_BRESP[17];
            assign AP_AXIMM_17_BVALID = ap_BVALID[17];
            assign ap_BREADY[17] = AP_AXIMM_17_BREADY;
            assign ap_ARADDR[17][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_17_ARADDR;
            assign ap_ARLEN[17] = AP_AXIMM_17_ARLEN;
            assign ap_ARSIZE[17] = AP_AXIMM_17_ARSIZE;
            assign ap_ARBURST[17] = AP_AXIMM_17_ARBURST;
            assign ap_ARLOCK[17] = AP_AXIMM_17_ARLOCK;
            assign ap_ARCACHE[17] = AP_AXIMM_17_ARCACHE;
            assign ap_ARPROT[17] = AP_AXIMM_17_ARPROT;
            assign ap_ARREGION[17] = AP_AXIMM_17_ARREGION;
            assign ap_ARQOS[17] = AP_AXIMM_17_ARQOS;
            assign ap_ARVALID[17] = AP_AXIMM_17_ARVALID;
            assign AP_AXIMM_17_ARREADY = ap_ARREADY[17];
            assign AP_AXIMM_17_RDATA = ap_RDATA[17][M_AXIMM_17_DATA_WIDTH-1:0];
            assign AP_AXIMM_17_RRESP = ap_RRESP[17];
            assign AP_AXIMM_17_RLAST = ap_RLAST[17];
            assign AP_AXIMM_17_RVALID = ap_RVALID[17];
            assign ap_RREADY[17] = AP_AXIMM_17_RREADY;
            assign M_AXIMM_17_AWADDR = dm_AWADDR[17][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_17_AWLEN = dm_AWLEN[17];
            assign M_AXIMM_17_AWSIZE = dm_AWSIZE[17];
            assign M_AXIMM_17_AWBURST = dm_AWBURST[17];
            assign M_AXIMM_17_AWLOCK = dm_AWLOCK[17];
            assign M_AXIMM_17_AWCACHE = dm_AWCACHE[17];
            assign M_AXIMM_17_AWPROT = dm_AWPROT[17];
            assign M_AXIMM_17_AWREGION = dm_AWREGION[17];
            assign M_AXIMM_17_AWQOS = dm_AWQOS[17];
            assign M_AXIMM_17_AWVALID = dm_AWVALID[17];
            assign dm_AWREADY[17] = M_AXIMM_17_AWREADY;
            assign M_AXIMM_17_WDATA = dm_WDATA[17][M_AXIMM_17_DATA_WIDTH-1:0];
            assign M_AXIMM_17_WSTRB = dm_WSTRB[17][M_AXIMM_17_DATA_WIDTH/8-1:0];
            assign M_AXIMM_17_WLAST = dm_WLAST[17];
            assign M_AXIMM_17_WVALID = dm_WVALID[17];
            assign dm_WREADY[17] = M_AXIMM_17_WREADY;
            assign dm_BRESP[17] = M_AXIMM_17_BRESP;
            assign dm_BVALID[17] = M_AXIMM_17_BVALID;
            assign M_AXIMM_17_BREADY = dm_BREADY[17];
            assign M_AXIMM_17_ARADDR = dm_ARADDR[17][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_17_ARLEN = dm_ARLEN[17];
            assign M_AXIMM_17_ARSIZE = dm_ARSIZE[17];
            assign M_AXIMM_17_ARBURST = dm_ARBURST[17];
            assign M_AXIMM_17_ARLOCK = dm_ARLOCK[17];
            assign M_AXIMM_17_ARCACHE = dm_ARCACHE[17];
            assign M_AXIMM_17_ARPROT = dm_ARPROT[17];
            assign M_AXIMM_17_ARREGION = dm_ARREGION[17];
            assign M_AXIMM_17_ARQOS = dm_ARQOS[17];
            assign M_AXIMM_17_ARVALID = dm_ARVALID[17];
            assign dm_ARREADY[17] = M_AXIMM_17_ARREADY;
            assign dm_RDATA[17][M_AXIMM_17_DATA_WIDTH-1:0] = M_AXIMM_17_RDATA;
            assign dm_RRESP[17] = M_AXIMM_17_RRESP;
            assign dm_RLAST[17] = M_AXIMM_17_RLAST;
            assign dm_RVALID[17] = M_AXIMM_17_RVALID;
            assign M_AXIMM_17_RREADY = dm_RREADY[17];
        end
        if(C_NUM_AXIMMs > 18) begin
            assign ap_AWADDR[18][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_18_AWADDR;
            assign ap_AWLEN[18] = AP_AXIMM_18_AWLEN;
            assign ap_AWSIZE[18] = AP_AXIMM_18_AWSIZE;
            assign ap_AWBURST[18] = AP_AXIMM_18_AWBURST;
            assign ap_AWLOCK[18] = AP_AXIMM_18_AWLOCK;
            assign ap_AWCACHE[18] = AP_AXIMM_18_AWCACHE;
            assign ap_AWPROT[18] = AP_AXIMM_18_AWPROT;
            assign ap_AWREGION[18] = AP_AXIMM_18_AWREGION;
            assign ap_AWQOS[18] = AP_AXIMM_18_AWQOS;
            assign ap_AWVALID[18] = AP_AXIMM_18_AWVALID;
            assign AP_AXIMM_18_AWREADY = ap_AWREADY[18];
            assign ap_WDATA[18][M_AXIMM_18_DATA_WIDTH-1:0] = AP_AXIMM_18_WDATA;
            assign ap_WSTRB[18][M_AXIMM_18_DATA_WIDTH/8-1:0] = AP_AXIMM_18_WSTRB;
            assign ap_WLAST[18] = AP_AXIMM_18_WLAST;
            assign ap_WVALID[18] = AP_AXIMM_18_WVALID;
            assign AP_AXIMM_18_WREADY = ap_WREADY[18];
            assign AP_AXIMM_18_BRESP = ap_BRESP[18];
            assign AP_AXIMM_18_BVALID = ap_BVALID[18];
            assign ap_BREADY[18] = AP_AXIMM_18_BREADY;
            assign ap_ARADDR[18][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_18_ARADDR;
            assign ap_ARLEN[18] = AP_AXIMM_18_ARLEN;
            assign ap_ARSIZE[18] = AP_AXIMM_18_ARSIZE;
            assign ap_ARBURST[18] = AP_AXIMM_18_ARBURST;
            assign ap_ARLOCK[18] = AP_AXIMM_18_ARLOCK;
            assign ap_ARCACHE[18] = AP_AXIMM_18_ARCACHE;
            assign ap_ARPROT[18] = AP_AXIMM_18_ARPROT;
            assign ap_ARREGION[18] = AP_AXIMM_18_ARREGION;
            assign ap_ARQOS[18] = AP_AXIMM_18_ARQOS;
            assign ap_ARVALID[18] = AP_AXIMM_18_ARVALID;
            assign AP_AXIMM_18_ARREADY = ap_ARREADY[18];
            assign AP_AXIMM_18_RDATA = ap_RDATA[18][M_AXIMM_18_DATA_WIDTH-1:0];
            assign AP_AXIMM_18_RRESP = ap_RRESP[18];
            assign AP_AXIMM_18_RLAST = ap_RLAST[18];
            assign AP_AXIMM_18_RVALID = ap_RVALID[18];
            assign ap_RREADY[18] = AP_AXIMM_18_RREADY;
            assign M_AXIMM_18_AWADDR = dm_AWADDR[18][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_18_AWLEN = dm_AWLEN[18];
            assign M_AXIMM_18_AWSIZE = dm_AWSIZE[18];
            assign M_AXIMM_18_AWBURST = dm_AWBURST[18];
            assign M_AXIMM_18_AWLOCK = dm_AWLOCK[18];
            assign M_AXIMM_18_AWCACHE = dm_AWCACHE[18];
            assign M_AXIMM_18_AWPROT = dm_AWPROT[18];
            assign M_AXIMM_18_AWREGION = dm_AWREGION[18];
            assign M_AXIMM_18_AWQOS = dm_AWQOS[18];
            assign M_AXIMM_18_AWVALID = dm_AWVALID[18];
            assign dm_AWREADY[18] = M_AXIMM_18_AWREADY;
            assign M_AXIMM_18_WDATA = dm_WDATA[18][M_AXIMM_18_DATA_WIDTH-1:0];
            assign M_AXIMM_18_WSTRB = dm_WSTRB[18][M_AXIMM_18_DATA_WIDTH/8-1:0];
            assign M_AXIMM_18_WLAST = dm_WLAST[18];
            assign M_AXIMM_18_WVALID = dm_WVALID[18];
            assign dm_WREADY[18] = M_AXIMM_18_WREADY;
            assign dm_BRESP[18] = M_AXIMM_18_BRESP;
            assign dm_BVALID[18] = M_AXIMM_18_BVALID;
            assign M_AXIMM_18_BREADY = dm_BREADY[18];
            assign M_AXIMM_18_ARADDR = dm_ARADDR[18][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_18_ARLEN = dm_ARLEN[18];
            assign M_AXIMM_18_ARSIZE = dm_ARSIZE[18];
            assign M_AXIMM_18_ARBURST = dm_ARBURST[18];
            assign M_AXIMM_18_ARLOCK = dm_ARLOCK[18];
            assign M_AXIMM_18_ARCACHE = dm_ARCACHE[18];
            assign M_AXIMM_18_ARPROT = dm_ARPROT[18];
            assign M_AXIMM_18_ARREGION = dm_ARREGION[18];
            assign M_AXIMM_18_ARQOS = dm_ARQOS[18];
            assign M_AXIMM_18_ARVALID = dm_ARVALID[18];
            assign dm_ARREADY[18] = M_AXIMM_18_ARREADY;
            assign dm_RDATA[18][M_AXIMM_18_DATA_WIDTH-1:0] = M_AXIMM_18_RDATA;
            assign dm_RRESP[18] = M_AXIMM_18_RRESP;
            assign dm_RLAST[18] = M_AXIMM_18_RLAST;
            assign dm_RVALID[18] = M_AXIMM_18_RVALID;
            assign M_AXIMM_18_RREADY = dm_RREADY[18];
        end
        if(C_NUM_AXIMMs > 19) begin
            assign ap_AWADDR[19][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_19_AWADDR;
            assign ap_AWLEN[19] = AP_AXIMM_19_AWLEN;
            assign ap_AWSIZE[19] = AP_AXIMM_19_AWSIZE;
            assign ap_AWBURST[19] = AP_AXIMM_19_AWBURST;
            assign ap_AWLOCK[19] = AP_AXIMM_19_AWLOCK;
            assign ap_AWCACHE[19] = AP_AXIMM_19_AWCACHE;
            assign ap_AWPROT[19] = AP_AXIMM_19_AWPROT;
            assign ap_AWREGION[19] = AP_AXIMM_19_AWREGION;
            assign ap_AWQOS[19] = AP_AXIMM_19_AWQOS;
            assign ap_AWVALID[19] = AP_AXIMM_19_AWVALID;
            assign AP_AXIMM_19_AWREADY = ap_AWREADY[19];
            assign ap_WDATA[19][M_AXIMM_19_DATA_WIDTH-1:0] = AP_AXIMM_19_WDATA;
            assign ap_WSTRB[19][M_AXIMM_19_DATA_WIDTH/8-1:0] = AP_AXIMM_19_WSTRB;
            assign ap_WLAST[19] = AP_AXIMM_19_WLAST;
            assign ap_WVALID[19] = AP_AXIMM_19_WVALID;
            assign AP_AXIMM_19_WREADY = ap_WREADY[19];
            assign AP_AXIMM_19_BRESP = ap_BRESP[19];
            assign AP_AXIMM_19_BVALID = ap_BVALID[19];
            assign ap_BREADY[19] = AP_AXIMM_19_BREADY;
            assign ap_ARADDR[19][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_19_ARADDR;
            assign ap_ARLEN[19] = AP_AXIMM_19_ARLEN;
            assign ap_ARSIZE[19] = AP_AXIMM_19_ARSIZE;
            assign ap_ARBURST[19] = AP_AXIMM_19_ARBURST;
            assign ap_ARLOCK[19] = AP_AXIMM_19_ARLOCK;
            assign ap_ARCACHE[19] = AP_AXIMM_19_ARCACHE;
            assign ap_ARPROT[19] = AP_AXIMM_19_ARPROT;
            assign ap_ARREGION[19] = AP_AXIMM_19_ARREGION;
            assign ap_ARQOS[19] = AP_AXIMM_19_ARQOS;
            assign ap_ARVALID[19] = AP_AXIMM_19_ARVALID;
            assign AP_AXIMM_19_ARREADY = ap_ARREADY[19];
            assign AP_AXIMM_19_RDATA = ap_RDATA[19][M_AXIMM_19_DATA_WIDTH-1:0];
            assign AP_AXIMM_19_RRESP = ap_RRESP[19];
            assign AP_AXIMM_19_RLAST = ap_RLAST[19];
            assign AP_AXIMM_19_RVALID = ap_RVALID[19];
            assign ap_RREADY[19] = AP_AXIMM_19_RREADY;
            assign M_AXIMM_19_AWADDR = dm_AWADDR[19][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_19_AWLEN = dm_AWLEN[19];
            assign M_AXIMM_19_AWSIZE = dm_AWSIZE[19];
            assign M_AXIMM_19_AWBURST = dm_AWBURST[19];
            assign M_AXIMM_19_AWLOCK = dm_AWLOCK[19];
            assign M_AXIMM_19_AWCACHE = dm_AWCACHE[19];
            assign M_AXIMM_19_AWPROT = dm_AWPROT[19];
            assign M_AXIMM_19_AWREGION = dm_AWREGION[19];
            assign M_AXIMM_19_AWQOS = dm_AWQOS[19];
            assign M_AXIMM_19_AWVALID = dm_AWVALID[19];
            assign dm_AWREADY[19] = M_AXIMM_19_AWREADY;
            assign M_AXIMM_19_WDATA = dm_WDATA[19][M_AXIMM_19_DATA_WIDTH-1:0];
            assign M_AXIMM_19_WSTRB = dm_WSTRB[19][M_AXIMM_19_DATA_WIDTH/8-1:0];
            assign M_AXIMM_19_WLAST = dm_WLAST[19];
            assign M_AXIMM_19_WVALID = dm_WVALID[19];
            assign dm_WREADY[19] = M_AXIMM_19_WREADY;
            assign dm_BRESP[19] = M_AXIMM_19_BRESP;
            assign dm_BVALID[19] = M_AXIMM_19_BVALID;
            assign M_AXIMM_19_BREADY = dm_BREADY[19];
            assign M_AXIMM_19_ARADDR = dm_ARADDR[19][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_19_ARLEN = dm_ARLEN[19];
            assign M_AXIMM_19_ARSIZE = dm_ARSIZE[19];
            assign M_AXIMM_19_ARBURST = dm_ARBURST[19];
            assign M_AXIMM_19_ARLOCK = dm_ARLOCK[19];
            assign M_AXIMM_19_ARCACHE = dm_ARCACHE[19];
            assign M_AXIMM_19_ARPROT = dm_ARPROT[19];
            assign M_AXIMM_19_ARREGION = dm_ARREGION[19];
            assign M_AXIMM_19_ARQOS = dm_ARQOS[19];
            assign M_AXIMM_19_ARVALID = dm_ARVALID[19];
            assign dm_ARREADY[19] = M_AXIMM_19_ARREADY;
            assign dm_RDATA[19][M_AXIMM_19_DATA_WIDTH-1:0] = M_AXIMM_19_RDATA;
            assign dm_RRESP[19] = M_AXIMM_19_RRESP;
            assign dm_RLAST[19] = M_AXIMM_19_RLAST;
            assign dm_RVALID[19] = M_AXIMM_19_RVALID;
            assign M_AXIMM_19_RREADY = dm_RREADY[19];
        end
        if(C_NUM_AXIMMs > 20) begin
            assign ap_AWADDR[20][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_20_AWADDR;
            assign ap_AWLEN[20] = AP_AXIMM_20_AWLEN;
            assign ap_AWSIZE[20] = AP_AXIMM_20_AWSIZE;
            assign ap_AWBURST[20] = AP_AXIMM_20_AWBURST;
            assign ap_AWLOCK[20] = AP_AXIMM_20_AWLOCK;
            assign ap_AWCACHE[20] = AP_AXIMM_20_AWCACHE;
            assign ap_AWPROT[20] = AP_AXIMM_20_AWPROT;
            assign ap_AWREGION[20] = AP_AXIMM_20_AWREGION;
            assign ap_AWQOS[20] = AP_AXIMM_20_AWQOS;
            assign ap_AWVALID[20] = AP_AXIMM_20_AWVALID;
            assign AP_AXIMM_20_AWREADY = ap_AWREADY[20];
            assign ap_WDATA[20][M_AXIMM_20_DATA_WIDTH-1:0] = AP_AXIMM_20_WDATA;
            assign ap_WSTRB[20][M_AXIMM_20_DATA_WIDTH/8-1:0] = AP_AXIMM_20_WSTRB;
            assign ap_WLAST[20] = AP_AXIMM_20_WLAST;
            assign ap_WVALID[20] = AP_AXIMM_20_WVALID;
            assign AP_AXIMM_20_WREADY = ap_WREADY[20];
            assign AP_AXIMM_20_BRESP = ap_BRESP[20];
            assign AP_AXIMM_20_BVALID = ap_BVALID[20];
            assign ap_BREADY[20] = AP_AXIMM_20_BREADY;
            assign ap_ARADDR[20][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_20_ARADDR;
            assign ap_ARLEN[20] = AP_AXIMM_20_ARLEN;
            assign ap_ARSIZE[20] = AP_AXIMM_20_ARSIZE;
            assign ap_ARBURST[20] = AP_AXIMM_20_ARBURST;
            assign ap_ARLOCK[20] = AP_AXIMM_20_ARLOCK;
            assign ap_ARCACHE[20] = AP_AXIMM_20_ARCACHE;
            assign ap_ARPROT[20] = AP_AXIMM_20_ARPROT;
            assign ap_ARREGION[20] = AP_AXIMM_20_ARREGION;
            assign ap_ARQOS[20] = AP_AXIMM_20_ARQOS;
            assign ap_ARVALID[20] = AP_AXIMM_20_ARVALID;
            assign AP_AXIMM_20_ARREADY = ap_ARREADY[20];
            assign AP_AXIMM_20_RDATA = ap_RDATA[20][M_AXIMM_20_DATA_WIDTH-1:0];
            assign AP_AXIMM_20_RRESP = ap_RRESP[20];
            assign AP_AXIMM_20_RLAST = ap_RLAST[20];
            assign AP_AXIMM_20_RVALID = ap_RVALID[20];
            assign ap_RREADY[20] = AP_AXIMM_20_RREADY;
            assign M_AXIMM_20_AWADDR = dm_AWADDR[20][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_20_AWLEN = dm_AWLEN[20];
            assign M_AXIMM_20_AWSIZE = dm_AWSIZE[20];
            assign M_AXIMM_20_AWBURST = dm_AWBURST[20];
            assign M_AXIMM_20_AWLOCK = dm_AWLOCK[20];
            assign M_AXIMM_20_AWCACHE = dm_AWCACHE[20];
            assign M_AXIMM_20_AWPROT = dm_AWPROT[20];
            assign M_AXIMM_20_AWREGION = dm_AWREGION[20];
            assign M_AXIMM_20_AWQOS = dm_AWQOS[20];
            assign M_AXIMM_20_AWVALID = dm_AWVALID[20];
            assign dm_AWREADY[20] = M_AXIMM_20_AWREADY;
            assign M_AXIMM_20_WDATA = dm_WDATA[20][M_AXIMM_20_DATA_WIDTH-1:0];
            assign M_AXIMM_20_WSTRB = dm_WSTRB[20][M_AXIMM_20_DATA_WIDTH/8-1:0];
            assign M_AXIMM_20_WLAST = dm_WLAST[20];
            assign M_AXIMM_20_WVALID = dm_WVALID[20];
            assign dm_WREADY[20] = M_AXIMM_20_WREADY;
            assign dm_BRESP[20] = M_AXIMM_20_BRESP;
            assign dm_BVALID[20] = M_AXIMM_20_BVALID;
            assign M_AXIMM_20_BREADY = dm_BREADY[20];
            assign M_AXIMM_20_ARADDR = dm_ARADDR[20][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_20_ARLEN = dm_ARLEN[20];
            assign M_AXIMM_20_ARSIZE = dm_ARSIZE[20];
            assign M_AXIMM_20_ARBURST = dm_ARBURST[20];
            assign M_AXIMM_20_ARLOCK = dm_ARLOCK[20];
            assign M_AXIMM_20_ARCACHE = dm_ARCACHE[20];
            assign M_AXIMM_20_ARPROT = dm_ARPROT[20];
            assign M_AXIMM_20_ARREGION = dm_ARREGION[20];
            assign M_AXIMM_20_ARQOS = dm_ARQOS[20];
            assign M_AXIMM_20_ARVALID = dm_ARVALID[20];
            assign dm_ARREADY[20] = M_AXIMM_20_ARREADY;
            assign dm_RDATA[20][M_AXIMM_20_DATA_WIDTH-1:0] = M_AXIMM_20_RDATA;
            assign dm_RRESP[20] = M_AXIMM_20_RRESP;
            assign dm_RLAST[20] = M_AXIMM_20_RLAST;
            assign dm_RVALID[20] = M_AXIMM_20_RVALID;
            assign M_AXIMM_20_RREADY = dm_RREADY[20];
        end
        if(C_NUM_AXIMMs > 21) begin
            assign ap_AWADDR[21][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_21_AWADDR;
            assign ap_AWLEN[21] = AP_AXIMM_21_AWLEN;
            assign ap_AWSIZE[21] = AP_AXIMM_21_AWSIZE;
            assign ap_AWBURST[21] = AP_AXIMM_21_AWBURST;
            assign ap_AWLOCK[21] = AP_AXIMM_21_AWLOCK;
            assign ap_AWCACHE[21] = AP_AXIMM_21_AWCACHE;
            assign ap_AWPROT[21] = AP_AXIMM_21_AWPROT;
            assign ap_AWREGION[21] = AP_AXIMM_21_AWREGION;
            assign ap_AWQOS[21] = AP_AXIMM_21_AWQOS;
            assign ap_AWVALID[21] = AP_AXIMM_21_AWVALID;
            assign AP_AXIMM_21_AWREADY = ap_AWREADY[21];
            assign ap_WDATA[21][M_AXIMM_21_DATA_WIDTH-1:0] = AP_AXIMM_21_WDATA;
            assign ap_WSTRB[21][M_AXIMM_21_DATA_WIDTH/8-1:0] = AP_AXIMM_21_WSTRB;
            assign ap_WLAST[21] = AP_AXIMM_21_WLAST;
            assign ap_WVALID[21] = AP_AXIMM_21_WVALID;
            assign AP_AXIMM_21_WREADY = ap_WREADY[21];
            assign AP_AXIMM_21_BRESP = ap_BRESP[21];
            assign AP_AXIMM_21_BVALID = ap_BVALID[21];
            assign ap_BREADY[21] = AP_AXIMM_21_BREADY;
            assign ap_ARADDR[21][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_21_ARADDR;
            assign ap_ARLEN[21] = AP_AXIMM_21_ARLEN;
            assign ap_ARSIZE[21] = AP_AXIMM_21_ARSIZE;
            assign ap_ARBURST[21] = AP_AXIMM_21_ARBURST;
            assign ap_ARLOCK[21] = AP_AXIMM_21_ARLOCK;
            assign ap_ARCACHE[21] = AP_AXIMM_21_ARCACHE;
            assign ap_ARPROT[21] = AP_AXIMM_21_ARPROT;
            assign ap_ARREGION[21] = AP_AXIMM_21_ARREGION;
            assign ap_ARQOS[21] = AP_AXIMM_21_ARQOS;
            assign ap_ARVALID[21] = AP_AXIMM_21_ARVALID;
            assign AP_AXIMM_21_ARREADY = ap_ARREADY[21];
            assign AP_AXIMM_21_RDATA = ap_RDATA[21][M_AXIMM_21_DATA_WIDTH-1:0];
            assign AP_AXIMM_21_RRESP = ap_RRESP[21];
            assign AP_AXIMM_21_RLAST = ap_RLAST[21];
            assign AP_AXIMM_21_RVALID = ap_RVALID[21];
            assign ap_RREADY[21] = AP_AXIMM_21_RREADY;
            assign M_AXIMM_21_AWADDR = dm_AWADDR[21][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_21_AWLEN = dm_AWLEN[21];
            assign M_AXIMM_21_AWSIZE = dm_AWSIZE[21];
            assign M_AXIMM_21_AWBURST = dm_AWBURST[21];
            assign M_AXIMM_21_AWLOCK = dm_AWLOCK[21];
            assign M_AXIMM_21_AWCACHE = dm_AWCACHE[21];
            assign M_AXIMM_21_AWPROT = dm_AWPROT[21];
            assign M_AXIMM_21_AWREGION = dm_AWREGION[21];
            assign M_AXIMM_21_AWQOS = dm_AWQOS[21];
            assign M_AXIMM_21_AWVALID = dm_AWVALID[21];
            assign dm_AWREADY[21] = M_AXIMM_21_AWREADY;
            assign M_AXIMM_21_WDATA = dm_WDATA[21][M_AXIMM_21_DATA_WIDTH-1:0];
            assign M_AXIMM_21_WSTRB = dm_WSTRB[21][M_AXIMM_21_DATA_WIDTH/8-1:0];
            assign M_AXIMM_21_WLAST = dm_WLAST[21];
            assign M_AXIMM_21_WVALID = dm_WVALID[21];
            assign dm_WREADY[21] = M_AXIMM_21_WREADY;
            assign dm_BRESP[21] = M_AXIMM_21_BRESP;
            assign dm_BVALID[21] = M_AXIMM_21_BVALID;
            assign M_AXIMM_21_BREADY = dm_BREADY[21];
            assign M_AXIMM_21_ARADDR = dm_ARADDR[21][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_21_ARLEN = dm_ARLEN[21];
            assign M_AXIMM_21_ARSIZE = dm_ARSIZE[21];
            assign M_AXIMM_21_ARBURST = dm_ARBURST[21];
            assign M_AXIMM_21_ARLOCK = dm_ARLOCK[21];
            assign M_AXIMM_21_ARCACHE = dm_ARCACHE[21];
            assign M_AXIMM_21_ARPROT = dm_ARPROT[21];
            assign M_AXIMM_21_ARREGION = dm_ARREGION[21];
            assign M_AXIMM_21_ARQOS = dm_ARQOS[21];
            assign M_AXIMM_21_ARVALID = dm_ARVALID[21];
            assign dm_ARREADY[21] = M_AXIMM_21_ARREADY;
            assign dm_RDATA[21][M_AXIMM_21_DATA_WIDTH-1:0] = M_AXIMM_21_RDATA;
            assign dm_RRESP[21] = M_AXIMM_21_RRESP;
            assign dm_RLAST[21] = M_AXIMM_21_RLAST;
            assign dm_RVALID[21] = M_AXIMM_21_RVALID;
            assign M_AXIMM_21_RREADY = dm_RREADY[21];
        end
        if(C_NUM_AXIMMs > 22) begin
            assign ap_AWADDR[22][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_22_AWADDR;
            assign ap_AWLEN[22] = AP_AXIMM_22_AWLEN;
            assign ap_AWSIZE[22] = AP_AXIMM_22_AWSIZE;
            assign ap_AWBURST[22] = AP_AXIMM_22_AWBURST;
            assign ap_AWLOCK[22] = AP_AXIMM_22_AWLOCK;
            assign ap_AWCACHE[22] = AP_AXIMM_22_AWCACHE;
            assign ap_AWPROT[22] = AP_AXIMM_22_AWPROT;
            assign ap_AWREGION[22] = AP_AXIMM_22_AWREGION;
            assign ap_AWQOS[22] = AP_AXIMM_22_AWQOS;
            assign ap_AWVALID[22] = AP_AXIMM_22_AWVALID;
            assign AP_AXIMM_22_AWREADY = ap_AWREADY[22];
            assign ap_WDATA[22][M_AXIMM_22_DATA_WIDTH-1:0] = AP_AXIMM_22_WDATA;
            assign ap_WSTRB[22][M_AXIMM_22_DATA_WIDTH/8-1:0] = AP_AXIMM_22_WSTRB;
            assign ap_WLAST[22] = AP_AXIMM_22_WLAST;
            assign ap_WVALID[22] = AP_AXIMM_22_WVALID;
            assign AP_AXIMM_22_WREADY = ap_WREADY[22];
            assign AP_AXIMM_22_BRESP = ap_BRESP[22];
            assign AP_AXIMM_22_BVALID = ap_BVALID[22];
            assign ap_BREADY[22] = AP_AXIMM_22_BREADY;
            assign ap_ARADDR[22][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_22_ARADDR;
            assign ap_ARLEN[22] = AP_AXIMM_22_ARLEN;
            assign ap_ARSIZE[22] = AP_AXIMM_22_ARSIZE;
            assign ap_ARBURST[22] = AP_AXIMM_22_ARBURST;
            assign ap_ARLOCK[22] = AP_AXIMM_22_ARLOCK;
            assign ap_ARCACHE[22] = AP_AXIMM_22_ARCACHE;
            assign ap_ARPROT[22] = AP_AXIMM_22_ARPROT;
            assign ap_ARREGION[22] = AP_AXIMM_22_ARREGION;
            assign ap_ARQOS[22] = AP_AXIMM_22_ARQOS;
            assign ap_ARVALID[22] = AP_AXIMM_22_ARVALID;
            assign AP_AXIMM_22_ARREADY = ap_ARREADY[22];
            assign AP_AXIMM_22_RDATA = ap_RDATA[22][M_AXIMM_22_DATA_WIDTH-1:0];
            assign AP_AXIMM_22_RRESP = ap_RRESP[22];
            assign AP_AXIMM_22_RLAST = ap_RLAST[22];
            assign AP_AXIMM_22_RVALID = ap_RVALID[22];
            assign ap_RREADY[22] = AP_AXIMM_22_RREADY;
            assign M_AXIMM_22_AWADDR = dm_AWADDR[22][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_22_AWLEN = dm_AWLEN[22];
            assign M_AXIMM_22_AWSIZE = dm_AWSIZE[22];
            assign M_AXIMM_22_AWBURST = dm_AWBURST[22];
            assign M_AXIMM_22_AWLOCK = dm_AWLOCK[22];
            assign M_AXIMM_22_AWCACHE = dm_AWCACHE[22];
            assign M_AXIMM_22_AWPROT = dm_AWPROT[22];
            assign M_AXIMM_22_AWREGION = dm_AWREGION[22];
            assign M_AXIMM_22_AWQOS = dm_AWQOS[22];
            assign M_AXIMM_22_AWVALID = dm_AWVALID[22];
            assign dm_AWREADY[22] = M_AXIMM_22_AWREADY;
            assign M_AXIMM_22_WDATA = dm_WDATA[22][M_AXIMM_22_DATA_WIDTH-1:0];
            assign M_AXIMM_22_WSTRB = dm_WSTRB[22][M_AXIMM_22_DATA_WIDTH/8-1:0];
            assign M_AXIMM_22_WLAST = dm_WLAST[22];
            assign M_AXIMM_22_WVALID = dm_WVALID[22];
            assign dm_WREADY[22] = M_AXIMM_22_WREADY;
            assign dm_BRESP[22] = M_AXIMM_22_BRESP;
            assign dm_BVALID[22] = M_AXIMM_22_BVALID;
            assign M_AXIMM_22_BREADY = dm_BREADY[22];
            assign M_AXIMM_22_ARADDR = dm_ARADDR[22][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_22_ARLEN = dm_ARLEN[22];
            assign M_AXIMM_22_ARSIZE = dm_ARSIZE[22];
            assign M_AXIMM_22_ARBURST = dm_ARBURST[22];
            assign M_AXIMM_22_ARLOCK = dm_ARLOCK[22];
            assign M_AXIMM_22_ARCACHE = dm_ARCACHE[22];
            assign M_AXIMM_22_ARPROT = dm_ARPROT[22];
            assign M_AXIMM_22_ARREGION = dm_ARREGION[22];
            assign M_AXIMM_22_ARQOS = dm_ARQOS[22];
            assign M_AXIMM_22_ARVALID = dm_ARVALID[22];
            assign dm_ARREADY[22] = M_AXIMM_22_ARREADY;
            assign dm_RDATA[22][M_AXIMM_22_DATA_WIDTH-1:0] = M_AXIMM_22_RDATA;
            assign dm_RRESP[22] = M_AXIMM_22_RRESP;
            assign dm_RLAST[22] = M_AXIMM_22_RLAST;
            assign dm_RVALID[22] = M_AXIMM_22_RVALID;
            assign M_AXIMM_22_RREADY = dm_RREADY[22];
        end
        if(C_NUM_AXIMMs > 23) begin
            assign ap_AWADDR[23][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_23_AWADDR;
            assign ap_AWLEN[23] = AP_AXIMM_23_AWLEN;
            assign ap_AWSIZE[23] = AP_AXIMM_23_AWSIZE;
            assign ap_AWBURST[23] = AP_AXIMM_23_AWBURST;
            assign ap_AWLOCK[23] = AP_AXIMM_23_AWLOCK;
            assign ap_AWCACHE[23] = AP_AXIMM_23_AWCACHE;
            assign ap_AWPROT[23] = AP_AXIMM_23_AWPROT;
            assign ap_AWREGION[23] = AP_AXIMM_23_AWREGION;
            assign ap_AWQOS[23] = AP_AXIMM_23_AWQOS;
            assign ap_AWVALID[23] = AP_AXIMM_23_AWVALID;
            assign AP_AXIMM_23_AWREADY = ap_AWREADY[23];
            assign ap_WDATA[23][M_AXIMM_23_DATA_WIDTH-1:0] = AP_AXIMM_23_WDATA;
            assign ap_WSTRB[23][M_AXIMM_23_DATA_WIDTH/8-1:0] = AP_AXIMM_23_WSTRB;
            assign ap_WLAST[23] = AP_AXIMM_23_WLAST;
            assign ap_WVALID[23] = AP_AXIMM_23_WVALID;
            assign AP_AXIMM_23_WREADY = ap_WREADY[23];
            assign AP_AXIMM_23_BRESP = ap_BRESP[23];
            assign AP_AXIMM_23_BVALID = ap_BVALID[23];
            assign ap_BREADY[23] = AP_AXIMM_23_BREADY;
            assign ap_ARADDR[23][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_23_ARADDR;
            assign ap_ARLEN[23] = AP_AXIMM_23_ARLEN;
            assign ap_ARSIZE[23] = AP_AXIMM_23_ARSIZE;
            assign ap_ARBURST[23] = AP_AXIMM_23_ARBURST;
            assign ap_ARLOCK[23] = AP_AXIMM_23_ARLOCK;
            assign ap_ARCACHE[23] = AP_AXIMM_23_ARCACHE;
            assign ap_ARPROT[23] = AP_AXIMM_23_ARPROT;
            assign ap_ARREGION[23] = AP_AXIMM_23_ARREGION;
            assign ap_ARQOS[23] = AP_AXIMM_23_ARQOS;
            assign ap_ARVALID[23] = AP_AXIMM_23_ARVALID;
            assign AP_AXIMM_23_ARREADY = ap_ARREADY[23];
            assign AP_AXIMM_23_RDATA = ap_RDATA[23][M_AXIMM_23_DATA_WIDTH-1:0];
            assign AP_AXIMM_23_RRESP = ap_RRESP[23];
            assign AP_AXIMM_23_RLAST = ap_RLAST[23];
            assign AP_AXIMM_23_RVALID = ap_RVALID[23];
            assign ap_RREADY[23] = AP_AXIMM_23_RREADY;
            assign M_AXIMM_23_AWADDR = dm_AWADDR[23][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_23_AWLEN = dm_AWLEN[23];
            assign M_AXIMM_23_AWSIZE = dm_AWSIZE[23];
            assign M_AXIMM_23_AWBURST = dm_AWBURST[23];
            assign M_AXIMM_23_AWLOCK = dm_AWLOCK[23];
            assign M_AXIMM_23_AWCACHE = dm_AWCACHE[23];
            assign M_AXIMM_23_AWPROT = dm_AWPROT[23];
            assign M_AXIMM_23_AWREGION = dm_AWREGION[23];
            assign M_AXIMM_23_AWQOS = dm_AWQOS[23];
            assign M_AXIMM_23_AWVALID = dm_AWVALID[23];
            assign dm_AWREADY[23] = M_AXIMM_23_AWREADY;
            assign M_AXIMM_23_WDATA = dm_WDATA[23][M_AXIMM_23_DATA_WIDTH-1:0];
            assign M_AXIMM_23_WSTRB = dm_WSTRB[23][M_AXIMM_23_DATA_WIDTH/8-1:0];
            assign M_AXIMM_23_WLAST = dm_WLAST[23];
            assign M_AXIMM_23_WVALID = dm_WVALID[23];
            assign dm_WREADY[23] = M_AXIMM_23_WREADY;
            assign dm_BRESP[23] = M_AXIMM_23_BRESP;
            assign dm_BVALID[23] = M_AXIMM_23_BVALID;
            assign M_AXIMM_23_BREADY = dm_BREADY[23];
            assign M_AXIMM_23_ARADDR = dm_ARADDR[23][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_23_ARLEN = dm_ARLEN[23];
            assign M_AXIMM_23_ARSIZE = dm_ARSIZE[23];
            assign M_AXIMM_23_ARBURST = dm_ARBURST[23];
            assign M_AXIMM_23_ARLOCK = dm_ARLOCK[23];
            assign M_AXIMM_23_ARCACHE = dm_ARCACHE[23];
            assign M_AXIMM_23_ARPROT = dm_ARPROT[23];
            assign M_AXIMM_23_ARREGION = dm_ARREGION[23];
            assign M_AXIMM_23_ARQOS = dm_ARQOS[23];
            assign M_AXIMM_23_ARVALID = dm_ARVALID[23];
            assign dm_ARREADY[23] = M_AXIMM_23_ARREADY;
            assign dm_RDATA[23][M_AXIMM_23_DATA_WIDTH-1:0] = M_AXIMM_23_RDATA;
            assign dm_RRESP[23] = M_AXIMM_23_RRESP;
            assign dm_RLAST[23] = M_AXIMM_23_RLAST;
            assign dm_RVALID[23] = M_AXIMM_23_RVALID;
            assign M_AXIMM_23_RREADY = dm_RREADY[23];
        end
        if(C_NUM_AXIMMs > 24) begin
            assign ap_AWADDR[24][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_24_AWADDR;
            assign ap_AWLEN[24] = AP_AXIMM_24_AWLEN;
            assign ap_AWSIZE[24] = AP_AXIMM_24_AWSIZE;
            assign ap_AWBURST[24] = AP_AXIMM_24_AWBURST;
            assign ap_AWLOCK[24] = AP_AXIMM_24_AWLOCK;
            assign ap_AWCACHE[24] = AP_AXIMM_24_AWCACHE;
            assign ap_AWPROT[24] = AP_AXIMM_24_AWPROT;
            assign ap_AWREGION[24] = AP_AXIMM_24_AWREGION;
            assign ap_AWQOS[24] = AP_AXIMM_24_AWQOS;
            assign ap_AWVALID[24] = AP_AXIMM_24_AWVALID;
            assign AP_AXIMM_24_AWREADY = ap_AWREADY[24];
            assign ap_WDATA[24][M_AXIMM_24_DATA_WIDTH-1:0] = AP_AXIMM_24_WDATA;
            assign ap_WSTRB[24][M_AXIMM_24_DATA_WIDTH/8-1:0] = AP_AXIMM_24_WSTRB;
            assign ap_WLAST[24] = AP_AXIMM_24_WLAST;
            assign ap_WVALID[24] = AP_AXIMM_24_WVALID;
            assign AP_AXIMM_24_WREADY = ap_WREADY[24];
            assign AP_AXIMM_24_BRESP = ap_BRESP[24];
            assign AP_AXIMM_24_BVALID = ap_BVALID[24];
            assign ap_BREADY[24] = AP_AXIMM_24_BREADY;
            assign ap_ARADDR[24][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_24_ARADDR;
            assign ap_ARLEN[24] = AP_AXIMM_24_ARLEN;
            assign ap_ARSIZE[24] = AP_AXIMM_24_ARSIZE;
            assign ap_ARBURST[24] = AP_AXIMM_24_ARBURST;
            assign ap_ARLOCK[24] = AP_AXIMM_24_ARLOCK;
            assign ap_ARCACHE[24] = AP_AXIMM_24_ARCACHE;
            assign ap_ARPROT[24] = AP_AXIMM_24_ARPROT;
            assign ap_ARREGION[24] = AP_AXIMM_24_ARREGION;
            assign ap_ARQOS[24] = AP_AXIMM_24_ARQOS;
            assign ap_ARVALID[24] = AP_AXIMM_24_ARVALID;
            assign AP_AXIMM_24_ARREADY = ap_ARREADY[24];
            assign AP_AXIMM_24_RDATA = ap_RDATA[24][M_AXIMM_24_DATA_WIDTH-1:0];
            assign AP_AXIMM_24_RRESP = ap_RRESP[24];
            assign AP_AXIMM_24_RLAST = ap_RLAST[24];
            assign AP_AXIMM_24_RVALID = ap_RVALID[24];
            assign ap_RREADY[24] = AP_AXIMM_24_RREADY;
            assign M_AXIMM_24_AWADDR = dm_AWADDR[24][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_24_AWLEN = dm_AWLEN[24];
            assign M_AXIMM_24_AWSIZE = dm_AWSIZE[24];
            assign M_AXIMM_24_AWBURST = dm_AWBURST[24];
            assign M_AXIMM_24_AWLOCK = dm_AWLOCK[24];
            assign M_AXIMM_24_AWCACHE = dm_AWCACHE[24];
            assign M_AXIMM_24_AWPROT = dm_AWPROT[24];
            assign M_AXIMM_24_AWREGION = dm_AWREGION[24];
            assign M_AXIMM_24_AWQOS = dm_AWQOS[24];
            assign M_AXIMM_24_AWVALID = dm_AWVALID[24];
            assign dm_AWREADY[24] = M_AXIMM_24_AWREADY;
            assign M_AXIMM_24_WDATA = dm_WDATA[24][M_AXIMM_24_DATA_WIDTH-1:0];
            assign M_AXIMM_24_WSTRB = dm_WSTRB[24][M_AXIMM_24_DATA_WIDTH/8-1:0];
            assign M_AXIMM_24_WLAST = dm_WLAST[24];
            assign M_AXIMM_24_WVALID = dm_WVALID[24];
            assign dm_WREADY[24] = M_AXIMM_24_WREADY;
            assign dm_BRESP[24] = M_AXIMM_24_BRESP;
            assign dm_BVALID[24] = M_AXIMM_24_BVALID;
            assign M_AXIMM_24_BREADY = dm_BREADY[24];
            assign M_AXIMM_24_ARADDR = dm_ARADDR[24][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_24_ARLEN = dm_ARLEN[24];
            assign M_AXIMM_24_ARSIZE = dm_ARSIZE[24];
            assign M_AXIMM_24_ARBURST = dm_ARBURST[24];
            assign M_AXIMM_24_ARLOCK = dm_ARLOCK[24];
            assign M_AXIMM_24_ARCACHE = dm_ARCACHE[24];
            assign M_AXIMM_24_ARPROT = dm_ARPROT[24];
            assign M_AXIMM_24_ARREGION = dm_ARREGION[24];
            assign M_AXIMM_24_ARQOS = dm_ARQOS[24];
            assign M_AXIMM_24_ARVALID = dm_ARVALID[24];
            assign dm_ARREADY[24] = M_AXIMM_24_ARREADY;
            assign dm_RDATA[24][M_AXIMM_24_DATA_WIDTH-1:0] = M_AXIMM_24_RDATA;
            assign dm_RRESP[24] = M_AXIMM_24_RRESP;
            assign dm_RLAST[24] = M_AXIMM_24_RLAST;
            assign dm_RVALID[24] = M_AXIMM_24_RVALID;
            assign M_AXIMM_24_RREADY = dm_RREADY[24];
        end
        if(C_NUM_AXIMMs > 25) begin
            assign ap_AWADDR[25][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_25_AWADDR;
            assign ap_AWLEN[25] = AP_AXIMM_25_AWLEN;
            assign ap_AWSIZE[25] = AP_AXIMM_25_AWSIZE;
            assign ap_AWBURST[25] = AP_AXIMM_25_AWBURST;
            assign ap_AWLOCK[25] = AP_AXIMM_25_AWLOCK;
            assign ap_AWCACHE[25] = AP_AXIMM_25_AWCACHE;
            assign ap_AWPROT[25] = AP_AXIMM_25_AWPROT;
            assign ap_AWREGION[25] = AP_AXIMM_25_AWREGION;
            assign ap_AWQOS[25] = AP_AXIMM_25_AWQOS;
            assign ap_AWVALID[25] = AP_AXIMM_25_AWVALID;
            assign AP_AXIMM_25_AWREADY = ap_AWREADY[25];
            assign ap_WDATA[25][M_AXIMM_25_DATA_WIDTH-1:0] = AP_AXIMM_25_WDATA;
            assign ap_WSTRB[25][M_AXIMM_25_DATA_WIDTH/8-1:0] = AP_AXIMM_25_WSTRB;
            assign ap_WLAST[25] = AP_AXIMM_25_WLAST;
            assign ap_WVALID[25] = AP_AXIMM_25_WVALID;
            assign AP_AXIMM_25_WREADY = ap_WREADY[25];
            assign AP_AXIMM_25_BRESP = ap_BRESP[25];
            assign AP_AXIMM_25_BVALID = ap_BVALID[25];
            assign ap_BREADY[25] = AP_AXIMM_25_BREADY;
            assign ap_ARADDR[25][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_25_ARADDR;
            assign ap_ARLEN[25] = AP_AXIMM_25_ARLEN;
            assign ap_ARSIZE[25] = AP_AXIMM_25_ARSIZE;
            assign ap_ARBURST[25] = AP_AXIMM_25_ARBURST;
            assign ap_ARLOCK[25] = AP_AXIMM_25_ARLOCK;
            assign ap_ARCACHE[25] = AP_AXIMM_25_ARCACHE;
            assign ap_ARPROT[25] = AP_AXIMM_25_ARPROT;
            assign ap_ARREGION[25] = AP_AXIMM_25_ARREGION;
            assign ap_ARQOS[25] = AP_AXIMM_25_ARQOS;
            assign ap_ARVALID[25] = AP_AXIMM_25_ARVALID;
            assign AP_AXIMM_25_ARREADY = ap_ARREADY[25];
            assign AP_AXIMM_25_RDATA = ap_RDATA[25][M_AXIMM_25_DATA_WIDTH-1:0];
            assign AP_AXIMM_25_RRESP = ap_RRESP[25];
            assign AP_AXIMM_25_RLAST = ap_RLAST[25];
            assign AP_AXIMM_25_RVALID = ap_RVALID[25];
            assign ap_RREADY[25] = AP_AXIMM_25_RREADY;
            assign M_AXIMM_25_AWADDR = dm_AWADDR[25][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_25_AWLEN = dm_AWLEN[25];
            assign M_AXIMM_25_AWSIZE = dm_AWSIZE[25];
            assign M_AXIMM_25_AWBURST = dm_AWBURST[25];
            assign M_AXIMM_25_AWLOCK = dm_AWLOCK[25];
            assign M_AXIMM_25_AWCACHE = dm_AWCACHE[25];
            assign M_AXIMM_25_AWPROT = dm_AWPROT[25];
            assign M_AXIMM_25_AWREGION = dm_AWREGION[25];
            assign M_AXIMM_25_AWQOS = dm_AWQOS[25];
            assign M_AXIMM_25_AWVALID = dm_AWVALID[25];
            assign dm_AWREADY[25] = M_AXIMM_25_AWREADY;
            assign M_AXIMM_25_WDATA = dm_WDATA[25][M_AXIMM_25_DATA_WIDTH-1:0];
            assign M_AXIMM_25_WSTRB = dm_WSTRB[25][M_AXIMM_25_DATA_WIDTH/8-1:0];
            assign M_AXIMM_25_WLAST = dm_WLAST[25];
            assign M_AXIMM_25_WVALID = dm_WVALID[25];
            assign dm_WREADY[25] = M_AXIMM_25_WREADY;
            assign dm_BRESP[25] = M_AXIMM_25_BRESP;
            assign dm_BVALID[25] = M_AXIMM_25_BVALID;
            assign M_AXIMM_25_BREADY = dm_BREADY[25];
            assign M_AXIMM_25_ARADDR = dm_ARADDR[25][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_25_ARLEN = dm_ARLEN[25];
            assign M_AXIMM_25_ARSIZE = dm_ARSIZE[25];
            assign M_AXIMM_25_ARBURST = dm_ARBURST[25];
            assign M_AXIMM_25_ARLOCK = dm_ARLOCK[25];
            assign M_AXIMM_25_ARCACHE = dm_ARCACHE[25];
            assign M_AXIMM_25_ARPROT = dm_ARPROT[25];
            assign M_AXIMM_25_ARREGION = dm_ARREGION[25];
            assign M_AXIMM_25_ARQOS = dm_ARQOS[25];
            assign M_AXIMM_25_ARVALID = dm_ARVALID[25];
            assign dm_ARREADY[25] = M_AXIMM_25_ARREADY;
            assign dm_RDATA[25][M_AXIMM_25_DATA_WIDTH-1:0] = M_AXIMM_25_RDATA;
            assign dm_RRESP[25] = M_AXIMM_25_RRESP;
            assign dm_RLAST[25] = M_AXIMM_25_RLAST;
            assign dm_RVALID[25] = M_AXIMM_25_RVALID;
            assign M_AXIMM_25_RREADY = dm_RREADY[25];
        end
        if(C_NUM_AXIMMs > 26) begin
            assign ap_AWADDR[26][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_26_AWADDR;
            assign ap_AWLEN[26] = AP_AXIMM_26_AWLEN;
            assign ap_AWSIZE[26] = AP_AXIMM_26_AWSIZE;
            assign ap_AWBURST[26] = AP_AXIMM_26_AWBURST;
            assign ap_AWLOCK[26] = AP_AXIMM_26_AWLOCK;
            assign ap_AWCACHE[26] = AP_AXIMM_26_AWCACHE;
            assign ap_AWPROT[26] = AP_AXIMM_26_AWPROT;
            assign ap_AWREGION[26] = AP_AXIMM_26_AWREGION;
            assign ap_AWQOS[26] = AP_AXIMM_26_AWQOS;
            assign ap_AWVALID[26] = AP_AXIMM_26_AWVALID;
            assign AP_AXIMM_26_AWREADY = ap_AWREADY[26];
            assign ap_WDATA[26][M_AXIMM_26_DATA_WIDTH-1:0] = AP_AXIMM_26_WDATA;
            assign ap_WSTRB[26][M_AXIMM_26_DATA_WIDTH/8-1:0] = AP_AXIMM_26_WSTRB;
            assign ap_WLAST[26] = AP_AXIMM_26_WLAST;
            assign ap_WVALID[26] = AP_AXIMM_26_WVALID;
            assign AP_AXIMM_26_WREADY = ap_WREADY[26];
            assign AP_AXIMM_26_BRESP = ap_BRESP[26];
            assign AP_AXIMM_26_BVALID = ap_BVALID[26];
            assign ap_BREADY[26] = AP_AXIMM_26_BREADY;
            assign ap_ARADDR[26][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_26_ARADDR;
            assign ap_ARLEN[26] = AP_AXIMM_26_ARLEN;
            assign ap_ARSIZE[26] = AP_AXIMM_26_ARSIZE;
            assign ap_ARBURST[26] = AP_AXIMM_26_ARBURST;
            assign ap_ARLOCK[26] = AP_AXIMM_26_ARLOCK;
            assign ap_ARCACHE[26] = AP_AXIMM_26_ARCACHE;
            assign ap_ARPROT[26] = AP_AXIMM_26_ARPROT;
            assign ap_ARREGION[26] = AP_AXIMM_26_ARREGION;
            assign ap_ARQOS[26] = AP_AXIMM_26_ARQOS;
            assign ap_ARVALID[26] = AP_AXIMM_26_ARVALID;
            assign AP_AXIMM_26_ARREADY = ap_ARREADY[26];
            assign AP_AXIMM_26_RDATA = ap_RDATA[26][M_AXIMM_26_DATA_WIDTH-1:0];
            assign AP_AXIMM_26_RRESP = ap_RRESP[26];
            assign AP_AXIMM_26_RLAST = ap_RLAST[26];
            assign AP_AXIMM_26_RVALID = ap_RVALID[26];
            assign ap_RREADY[26] = AP_AXIMM_26_RREADY;
            assign M_AXIMM_26_AWADDR = dm_AWADDR[26][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_26_AWLEN = dm_AWLEN[26];
            assign M_AXIMM_26_AWSIZE = dm_AWSIZE[26];
            assign M_AXIMM_26_AWBURST = dm_AWBURST[26];
            assign M_AXIMM_26_AWLOCK = dm_AWLOCK[26];
            assign M_AXIMM_26_AWCACHE = dm_AWCACHE[26];
            assign M_AXIMM_26_AWPROT = dm_AWPROT[26];
            assign M_AXIMM_26_AWREGION = dm_AWREGION[26];
            assign M_AXIMM_26_AWQOS = dm_AWQOS[26];
            assign M_AXIMM_26_AWVALID = dm_AWVALID[26];
            assign dm_AWREADY[26] = M_AXIMM_26_AWREADY;
            assign M_AXIMM_26_WDATA = dm_WDATA[26][M_AXIMM_26_DATA_WIDTH-1:0];
            assign M_AXIMM_26_WSTRB = dm_WSTRB[26][M_AXIMM_26_DATA_WIDTH/8-1:0];
            assign M_AXIMM_26_WLAST = dm_WLAST[26];
            assign M_AXIMM_26_WVALID = dm_WVALID[26];
            assign dm_WREADY[26] = M_AXIMM_26_WREADY;
            assign dm_BRESP[26] = M_AXIMM_26_BRESP;
            assign dm_BVALID[26] = M_AXIMM_26_BVALID;
            assign M_AXIMM_26_BREADY = dm_BREADY[26];
            assign M_AXIMM_26_ARADDR = dm_ARADDR[26][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_26_ARLEN = dm_ARLEN[26];
            assign M_AXIMM_26_ARSIZE = dm_ARSIZE[26];
            assign M_AXIMM_26_ARBURST = dm_ARBURST[26];
            assign M_AXIMM_26_ARLOCK = dm_ARLOCK[26];
            assign M_AXIMM_26_ARCACHE = dm_ARCACHE[26];
            assign M_AXIMM_26_ARPROT = dm_ARPROT[26];
            assign M_AXIMM_26_ARREGION = dm_ARREGION[26];
            assign M_AXIMM_26_ARQOS = dm_ARQOS[26];
            assign M_AXIMM_26_ARVALID = dm_ARVALID[26];
            assign dm_ARREADY[26] = M_AXIMM_26_ARREADY;
            assign dm_RDATA[26][M_AXIMM_26_DATA_WIDTH-1:0] = M_AXIMM_26_RDATA;
            assign dm_RRESP[26] = M_AXIMM_26_RRESP;
            assign dm_RLAST[26] = M_AXIMM_26_RLAST;
            assign dm_RVALID[26] = M_AXIMM_26_RVALID;
            assign M_AXIMM_26_RREADY = dm_RREADY[26];
        end
        if(C_NUM_AXIMMs > 27) begin
            assign ap_AWADDR[27][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_27_AWADDR;
            assign ap_AWLEN[27] = AP_AXIMM_27_AWLEN;
            assign ap_AWSIZE[27] = AP_AXIMM_27_AWSIZE;
            assign ap_AWBURST[27] = AP_AXIMM_27_AWBURST;
            assign ap_AWLOCK[27] = AP_AXIMM_27_AWLOCK;
            assign ap_AWCACHE[27] = AP_AXIMM_27_AWCACHE;
            assign ap_AWPROT[27] = AP_AXIMM_27_AWPROT;
            assign ap_AWREGION[27] = AP_AXIMM_27_AWREGION;
            assign ap_AWQOS[27] = AP_AXIMM_27_AWQOS;
            assign ap_AWVALID[27] = AP_AXIMM_27_AWVALID;
            assign AP_AXIMM_27_AWREADY = ap_AWREADY[27];
            assign ap_WDATA[27][M_AXIMM_27_DATA_WIDTH-1:0] = AP_AXIMM_27_WDATA;
            assign ap_WSTRB[27][M_AXIMM_27_DATA_WIDTH/8-1:0] = AP_AXIMM_27_WSTRB;
            assign ap_WLAST[27] = AP_AXIMM_27_WLAST;
            assign ap_WVALID[27] = AP_AXIMM_27_WVALID;
            assign AP_AXIMM_27_WREADY = ap_WREADY[27];
            assign AP_AXIMM_27_BRESP = ap_BRESP[27];
            assign AP_AXIMM_27_BVALID = ap_BVALID[27];
            assign ap_BREADY[27] = AP_AXIMM_27_BREADY;
            assign ap_ARADDR[27][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_27_ARADDR;
            assign ap_ARLEN[27] = AP_AXIMM_27_ARLEN;
            assign ap_ARSIZE[27] = AP_AXIMM_27_ARSIZE;
            assign ap_ARBURST[27] = AP_AXIMM_27_ARBURST;
            assign ap_ARLOCK[27] = AP_AXIMM_27_ARLOCK;
            assign ap_ARCACHE[27] = AP_AXIMM_27_ARCACHE;
            assign ap_ARPROT[27] = AP_AXIMM_27_ARPROT;
            assign ap_ARREGION[27] = AP_AXIMM_27_ARREGION;
            assign ap_ARQOS[27] = AP_AXIMM_27_ARQOS;
            assign ap_ARVALID[27] = AP_AXIMM_27_ARVALID;
            assign AP_AXIMM_27_ARREADY = ap_ARREADY[27];
            assign AP_AXIMM_27_RDATA = ap_RDATA[27][M_AXIMM_27_DATA_WIDTH-1:0];
            assign AP_AXIMM_27_RRESP = ap_RRESP[27];
            assign AP_AXIMM_27_RLAST = ap_RLAST[27];
            assign AP_AXIMM_27_RVALID = ap_RVALID[27];
            assign ap_RREADY[27] = AP_AXIMM_27_RREADY;
            assign M_AXIMM_27_AWADDR = dm_AWADDR[27][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_27_AWLEN = dm_AWLEN[27];
            assign M_AXIMM_27_AWSIZE = dm_AWSIZE[27];
            assign M_AXIMM_27_AWBURST = dm_AWBURST[27];
            assign M_AXIMM_27_AWLOCK = dm_AWLOCK[27];
            assign M_AXIMM_27_AWCACHE = dm_AWCACHE[27];
            assign M_AXIMM_27_AWPROT = dm_AWPROT[27];
            assign M_AXIMM_27_AWREGION = dm_AWREGION[27];
            assign M_AXIMM_27_AWQOS = dm_AWQOS[27];
            assign M_AXIMM_27_AWVALID = dm_AWVALID[27];
            assign dm_AWREADY[27] = M_AXIMM_27_AWREADY;
            assign M_AXIMM_27_WDATA = dm_WDATA[27][M_AXIMM_27_DATA_WIDTH-1:0];
            assign M_AXIMM_27_WSTRB = dm_WSTRB[27][M_AXIMM_27_DATA_WIDTH/8-1:0];
            assign M_AXIMM_27_WLAST = dm_WLAST[27];
            assign M_AXIMM_27_WVALID = dm_WVALID[27];
            assign dm_WREADY[27] = M_AXIMM_27_WREADY;
            assign dm_BRESP[27] = M_AXIMM_27_BRESP;
            assign dm_BVALID[27] = M_AXIMM_27_BVALID;
            assign M_AXIMM_27_BREADY = dm_BREADY[27];
            assign M_AXIMM_27_ARADDR = dm_ARADDR[27][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_27_ARLEN = dm_ARLEN[27];
            assign M_AXIMM_27_ARSIZE = dm_ARSIZE[27];
            assign M_AXIMM_27_ARBURST = dm_ARBURST[27];
            assign M_AXIMM_27_ARLOCK = dm_ARLOCK[27];
            assign M_AXIMM_27_ARCACHE = dm_ARCACHE[27];
            assign M_AXIMM_27_ARPROT = dm_ARPROT[27];
            assign M_AXIMM_27_ARREGION = dm_ARREGION[27];
            assign M_AXIMM_27_ARQOS = dm_ARQOS[27];
            assign M_AXIMM_27_ARVALID = dm_ARVALID[27];
            assign dm_ARREADY[27] = M_AXIMM_27_ARREADY;
            assign dm_RDATA[27][M_AXIMM_27_DATA_WIDTH-1:0] = M_AXIMM_27_RDATA;
            assign dm_RRESP[27] = M_AXIMM_27_RRESP;
            assign dm_RLAST[27] = M_AXIMM_27_RLAST;
            assign dm_RVALID[27] = M_AXIMM_27_RVALID;
            assign M_AXIMM_27_RREADY = dm_RREADY[27];
        end
        if(C_NUM_AXIMMs > 28) begin
            assign ap_AWADDR[28][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_28_AWADDR;
            assign ap_AWLEN[28] = AP_AXIMM_28_AWLEN;
            assign ap_AWSIZE[28] = AP_AXIMM_28_AWSIZE;
            assign ap_AWBURST[28] = AP_AXIMM_28_AWBURST;
            assign ap_AWLOCK[28] = AP_AXIMM_28_AWLOCK;
            assign ap_AWCACHE[28] = AP_AXIMM_28_AWCACHE;
            assign ap_AWPROT[28] = AP_AXIMM_28_AWPROT;
            assign ap_AWREGION[28] = AP_AXIMM_28_AWREGION;
            assign ap_AWQOS[28] = AP_AXIMM_28_AWQOS;
            assign ap_AWVALID[28] = AP_AXIMM_28_AWVALID;
            assign AP_AXIMM_28_AWREADY = ap_AWREADY[28];
            assign ap_WDATA[28][M_AXIMM_28_DATA_WIDTH-1:0] = AP_AXIMM_28_WDATA;
            assign ap_WSTRB[28][M_AXIMM_28_DATA_WIDTH/8-1:0] = AP_AXIMM_28_WSTRB;
            assign ap_WLAST[28] = AP_AXIMM_28_WLAST;
            assign ap_WVALID[28] = AP_AXIMM_28_WVALID;
            assign AP_AXIMM_28_WREADY = ap_WREADY[28];
            assign AP_AXIMM_28_BRESP = ap_BRESP[28];
            assign AP_AXIMM_28_BVALID = ap_BVALID[28];
            assign ap_BREADY[28] = AP_AXIMM_28_BREADY;
            assign ap_ARADDR[28][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_28_ARADDR;
            assign ap_ARLEN[28] = AP_AXIMM_28_ARLEN;
            assign ap_ARSIZE[28] = AP_AXIMM_28_ARSIZE;
            assign ap_ARBURST[28] = AP_AXIMM_28_ARBURST;
            assign ap_ARLOCK[28] = AP_AXIMM_28_ARLOCK;
            assign ap_ARCACHE[28] = AP_AXIMM_28_ARCACHE;
            assign ap_ARPROT[28] = AP_AXIMM_28_ARPROT;
            assign ap_ARREGION[28] = AP_AXIMM_28_ARREGION;
            assign ap_ARQOS[28] = AP_AXIMM_28_ARQOS;
            assign ap_ARVALID[28] = AP_AXIMM_28_ARVALID;
            assign AP_AXIMM_28_ARREADY = ap_ARREADY[28];
            assign AP_AXIMM_28_RDATA = ap_RDATA[28][M_AXIMM_28_DATA_WIDTH-1:0];
            assign AP_AXIMM_28_RRESP = ap_RRESP[28];
            assign AP_AXIMM_28_RLAST = ap_RLAST[28];
            assign AP_AXIMM_28_RVALID = ap_RVALID[28];
            assign ap_RREADY[28] = AP_AXIMM_28_RREADY;
            assign M_AXIMM_28_AWADDR = dm_AWADDR[28][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_28_AWLEN = dm_AWLEN[28];
            assign M_AXIMM_28_AWSIZE = dm_AWSIZE[28];
            assign M_AXIMM_28_AWBURST = dm_AWBURST[28];
            assign M_AXIMM_28_AWLOCK = dm_AWLOCK[28];
            assign M_AXIMM_28_AWCACHE = dm_AWCACHE[28];
            assign M_AXIMM_28_AWPROT = dm_AWPROT[28];
            assign M_AXIMM_28_AWREGION = dm_AWREGION[28];
            assign M_AXIMM_28_AWQOS = dm_AWQOS[28];
            assign M_AXIMM_28_AWVALID = dm_AWVALID[28];
            assign dm_AWREADY[28] = M_AXIMM_28_AWREADY;
            assign M_AXIMM_28_WDATA = dm_WDATA[28][M_AXIMM_28_DATA_WIDTH-1:0];
            assign M_AXIMM_28_WSTRB = dm_WSTRB[28][M_AXIMM_28_DATA_WIDTH/8-1:0];
            assign M_AXIMM_28_WLAST = dm_WLAST[28];
            assign M_AXIMM_28_WVALID = dm_WVALID[28];
            assign dm_WREADY[28] = M_AXIMM_28_WREADY;
            assign dm_BRESP[28] = M_AXIMM_28_BRESP;
            assign dm_BVALID[28] = M_AXIMM_28_BVALID;
            assign M_AXIMM_28_BREADY = dm_BREADY[28];
            assign M_AXIMM_28_ARADDR = dm_ARADDR[28][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_28_ARLEN = dm_ARLEN[28];
            assign M_AXIMM_28_ARSIZE = dm_ARSIZE[28];
            assign M_AXIMM_28_ARBURST = dm_ARBURST[28];
            assign M_AXIMM_28_ARLOCK = dm_ARLOCK[28];
            assign M_AXIMM_28_ARCACHE = dm_ARCACHE[28];
            assign M_AXIMM_28_ARPROT = dm_ARPROT[28];
            assign M_AXIMM_28_ARREGION = dm_ARREGION[28];
            assign M_AXIMM_28_ARQOS = dm_ARQOS[28];
            assign M_AXIMM_28_ARVALID = dm_ARVALID[28];
            assign dm_ARREADY[28] = M_AXIMM_28_ARREADY;
            assign dm_RDATA[28][M_AXIMM_28_DATA_WIDTH-1:0] = M_AXIMM_28_RDATA;
            assign dm_RRESP[28] = M_AXIMM_28_RRESP;
            assign dm_RLAST[28] = M_AXIMM_28_RLAST;
            assign dm_RVALID[28] = M_AXIMM_28_RVALID;
            assign M_AXIMM_28_RREADY = dm_RREADY[28];
        end
        if(C_NUM_AXIMMs > 29) begin
            assign ap_AWADDR[29][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_29_AWADDR;
            assign ap_AWLEN[29] = AP_AXIMM_29_AWLEN;
            assign ap_AWSIZE[29] = AP_AXIMM_29_AWSIZE;
            assign ap_AWBURST[29] = AP_AXIMM_29_AWBURST;
            assign ap_AWLOCK[29] = AP_AXIMM_29_AWLOCK;
            assign ap_AWCACHE[29] = AP_AXIMM_29_AWCACHE;
            assign ap_AWPROT[29] = AP_AXIMM_29_AWPROT;
            assign ap_AWREGION[29] = AP_AXIMM_29_AWREGION;
            assign ap_AWQOS[29] = AP_AXIMM_29_AWQOS;
            assign ap_AWVALID[29] = AP_AXIMM_29_AWVALID;
            assign AP_AXIMM_29_AWREADY = ap_AWREADY[29];
            assign ap_WDATA[29][M_AXIMM_29_DATA_WIDTH-1:0] = AP_AXIMM_29_WDATA;
            assign ap_WSTRB[29][M_AXIMM_29_DATA_WIDTH/8-1:0] = AP_AXIMM_29_WSTRB;
            assign ap_WLAST[29] = AP_AXIMM_29_WLAST;
            assign ap_WVALID[29] = AP_AXIMM_29_WVALID;
            assign AP_AXIMM_29_WREADY = ap_WREADY[29];
            assign AP_AXIMM_29_BRESP = ap_BRESP[29];
            assign AP_AXIMM_29_BVALID = ap_BVALID[29];
            assign ap_BREADY[29] = AP_AXIMM_29_BREADY;
            assign ap_ARADDR[29][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_29_ARADDR;
            assign ap_ARLEN[29] = AP_AXIMM_29_ARLEN;
            assign ap_ARSIZE[29] = AP_AXIMM_29_ARSIZE;
            assign ap_ARBURST[29] = AP_AXIMM_29_ARBURST;
            assign ap_ARLOCK[29] = AP_AXIMM_29_ARLOCK;
            assign ap_ARCACHE[29] = AP_AXIMM_29_ARCACHE;
            assign ap_ARPROT[29] = AP_AXIMM_29_ARPROT;
            assign ap_ARREGION[29] = AP_AXIMM_29_ARREGION;
            assign ap_ARQOS[29] = AP_AXIMM_29_ARQOS;
            assign ap_ARVALID[29] = AP_AXIMM_29_ARVALID;
            assign AP_AXIMM_29_ARREADY = ap_ARREADY[29];
            assign AP_AXIMM_29_RDATA = ap_RDATA[29][M_AXIMM_29_DATA_WIDTH-1:0];
            assign AP_AXIMM_29_RRESP = ap_RRESP[29];
            assign AP_AXIMM_29_RLAST = ap_RLAST[29];
            assign AP_AXIMM_29_RVALID = ap_RVALID[29];
            assign ap_RREADY[29] = AP_AXIMM_29_RREADY;
            assign M_AXIMM_29_AWADDR = dm_AWADDR[29][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_29_AWLEN = dm_AWLEN[29];
            assign M_AXIMM_29_AWSIZE = dm_AWSIZE[29];
            assign M_AXIMM_29_AWBURST = dm_AWBURST[29];
            assign M_AXIMM_29_AWLOCK = dm_AWLOCK[29];
            assign M_AXIMM_29_AWCACHE = dm_AWCACHE[29];
            assign M_AXIMM_29_AWPROT = dm_AWPROT[29];
            assign M_AXIMM_29_AWREGION = dm_AWREGION[29];
            assign M_AXIMM_29_AWQOS = dm_AWQOS[29];
            assign M_AXIMM_29_AWVALID = dm_AWVALID[29];
            assign dm_AWREADY[29] = M_AXIMM_29_AWREADY;
            assign M_AXIMM_29_WDATA = dm_WDATA[29][M_AXIMM_29_DATA_WIDTH-1:0];
            assign M_AXIMM_29_WSTRB = dm_WSTRB[29][M_AXIMM_29_DATA_WIDTH/8-1:0];
            assign M_AXIMM_29_WLAST = dm_WLAST[29];
            assign M_AXIMM_29_WVALID = dm_WVALID[29];
            assign dm_WREADY[29] = M_AXIMM_29_WREADY;
            assign dm_BRESP[29] = M_AXIMM_29_BRESP;
            assign dm_BVALID[29] = M_AXIMM_29_BVALID;
            assign M_AXIMM_29_BREADY = dm_BREADY[29];
            assign M_AXIMM_29_ARADDR = dm_ARADDR[29][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_29_ARLEN = dm_ARLEN[29];
            assign M_AXIMM_29_ARSIZE = dm_ARSIZE[29];
            assign M_AXIMM_29_ARBURST = dm_ARBURST[29];
            assign M_AXIMM_29_ARLOCK = dm_ARLOCK[29];
            assign M_AXIMM_29_ARCACHE = dm_ARCACHE[29];
            assign M_AXIMM_29_ARPROT = dm_ARPROT[29];
            assign M_AXIMM_29_ARREGION = dm_ARREGION[29];
            assign M_AXIMM_29_ARQOS = dm_ARQOS[29];
            assign M_AXIMM_29_ARVALID = dm_ARVALID[29];
            assign dm_ARREADY[29] = M_AXIMM_29_ARREADY;
            assign dm_RDATA[29][M_AXIMM_29_DATA_WIDTH-1:0] = M_AXIMM_29_RDATA;
            assign dm_RRESP[29] = M_AXIMM_29_RRESP;
            assign dm_RLAST[29] = M_AXIMM_29_RLAST;
            assign dm_RVALID[29] = M_AXIMM_29_RVALID;
            assign M_AXIMM_29_RREADY = dm_RREADY[29];
        end
        if(C_NUM_AXIMMs > 30) begin
            assign ap_AWADDR[30][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_30_AWADDR;
            assign ap_AWLEN[30] = AP_AXIMM_30_AWLEN;
            assign ap_AWSIZE[30] = AP_AXIMM_30_AWSIZE;
            assign ap_AWBURST[30] = AP_AXIMM_30_AWBURST;
            assign ap_AWLOCK[30] = AP_AXIMM_30_AWLOCK;
            assign ap_AWCACHE[30] = AP_AXIMM_30_AWCACHE;
            assign ap_AWPROT[30] = AP_AXIMM_30_AWPROT;
            assign ap_AWREGION[30] = AP_AXIMM_30_AWREGION;
            assign ap_AWQOS[30] = AP_AXIMM_30_AWQOS;
            assign ap_AWVALID[30] = AP_AXIMM_30_AWVALID;
            assign AP_AXIMM_30_AWREADY = ap_AWREADY[30];
            assign ap_WDATA[30][M_AXIMM_30_DATA_WIDTH-1:0] = AP_AXIMM_30_WDATA;
            assign ap_WSTRB[30][M_AXIMM_30_DATA_WIDTH/8-1:0] = AP_AXIMM_30_WSTRB;
            assign ap_WLAST[30] = AP_AXIMM_30_WLAST;
            assign ap_WVALID[30] = AP_AXIMM_30_WVALID;
            assign AP_AXIMM_30_WREADY = ap_WREADY[30];
            assign AP_AXIMM_30_BRESP = ap_BRESP[30];
            assign AP_AXIMM_30_BVALID = ap_BVALID[30];
            assign ap_BREADY[30] = AP_AXIMM_30_BREADY;
            assign ap_ARADDR[30][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_30_ARADDR;
            assign ap_ARLEN[30] = AP_AXIMM_30_ARLEN;
            assign ap_ARSIZE[30] = AP_AXIMM_30_ARSIZE;
            assign ap_ARBURST[30] = AP_AXIMM_30_ARBURST;
            assign ap_ARLOCK[30] = AP_AXIMM_30_ARLOCK;
            assign ap_ARCACHE[30] = AP_AXIMM_30_ARCACHE;
            assign ap_ARPROT[30] = AP_AXIMM_30_ARPROT;
            assign ap_ARREGION[30] = AP_AXIMM_30_ARREGION;
            assign ap_ARQOS[30] = AP_AXIMM_30_ARQOS;
            assign ap_ARVALID[30] = AP_AXIMM_30_ARVALID;
            assign AP_AXIMM_30_ARREADY = ap_ARREADY[30];
            assign AP_AXIMM_30_RDATA = ap_RDATA[30][M_AXIMM_30_DATA_WIDTH-1:0];
            assign AP_AXIMM_30_RRESP = ap_RRESP[30];
            assign AP_AXIMM_30_RLAST = ap_RLAST[30];
            assign AP_AXIMM_30_RVALID = ap_RVALID[30];
            assign ap_RREADY[30] = AP_AXIMM_30_RREADY;
            assign M_AXIMM_30_AWADDR = dm_AWADDR[30][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_30_AWLEN = dm_AWLEN[30];
            assign M_AXIMM_30_AWSIZE = dm_AWSIZE[30];
            assign M_AXIMM_30_AWBURST = dm_AWBURST[30];
            assign M_AXIMM_30_AWLOCK = dm_AWLOCK[30];
            assign M_AXIMM_30_AWCACHE = dm_AWCACHE[30];
            assign M_AXIMM_30_AWPROT = dm_AWPROT[30];
            assign M_AXIMM_30_AWREGION = dm_AWREGION[30];
            assign M_AXIMM_30_AWQOS = dm_AWQOS[30];
            assign M_AXIMM_30_AWVALID = dm_AWVALID[30];
            assign dm_AWREADY[30] = M_AXIMM_30_AWREADY;
            assign M_AXIMM_30_WDATA = dm_WDATA[30][M_AXIMM_30_DATA_WIDTH-1:0];
            assign M_AXIMM_30_WSTRB = dm_WSTRB[30][M_AXIMM_30_DATA_WIDTH/8-1:0];
            assign M_AXIMM_30_WLAST = dm_WLAST[30];
            assign M_AXIMM_30_WVALID = dm_WVALID[30];
            assign dm_WREADY[30] = M_AXIMM_30_WREADY;
            assign dm_BRESP[30] = M_AXIMM_30_BRESP;
            assign dm_BVALID[30] = M_AXIMM_30_BVALID;
            assign M_AXIMM_30_BREADY = dm_BREADY[30];
            assign M_AXIMM_30_ARADDR = dm_ARADDR[30][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_30_ARLEN = dm_ARLEN[30];
            assign M_AXIMM_30_ARSIZE = dm_ARSIZE[30];
            assign M_AXIMM_30_ARBURST = dm_ARBURST[30];
            assign M_AXIMM_30_ARLOCK = dm_ARLOCK[30];
            assign M_AXIMM_30_ARCACHE = dm_ARCACHE[30];
            assign M_AXIMM_30_ARPROT = dm_ARPROT[30];
            assign M_AXIMM_30_ARREGION = dm_ARREGION[30];
            assign M_AXIMM_30_ARQOS = dm_ARQOS[30];
            assign M_AXIMM_30_ARVALID = dm_ARVALID[30];
            assign dm_ARREADY[30] = M_AXIMM_30_ARREADY;
            assign dm_RDATA[30][M_AXIMM_30_DATA_WIDTH-1:0] = M_AXIMM_30_RDATA;
            assign dm_RRESP[30] = M_AXIMM_30_RRESP;
            assign dm_RLAST[30] = M_AXIMM_30_RLAST;
            assign dm_RVALID[30] = M_AXIMM_30_RVALID;
            assign M_AXIMM_30_RREADY = dm_RREADY[30];
        end
        if(C_NUM_AXIMMs > 31) begin
            assign ap_AWADDR[31][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_31_AWADDR;
            assign ap_AWLEN[31] = AP_AXIMM_31_AWLEN;
            assign ap_AWSIZE[31] = AP_AXIMM_31_AWSIZE;
            assign ap_AWBURST[31] = AP_AXIMM_31_AWBURST;
            assign ap_AWLOCK[31] = AP_AXIMM_31_AWLOCK;
            assign ap_AWCACHE[31] = AP_AXIMM_31_AWCACHE;
            assign ap_AWPROT[31] = AP_AXIMM_31_AWPROT;
            assign ap_AWREGION[31] = AP_AXIMM_31_AWREGION;
            assign ap_AWQOS[31] = AP_AXIMM_31_AWQOS;
            assign ap_AWVALID[31] = AP_AXIMM_31_AWVALID;
            assign AP_AXIMM_31_AWREADY = ap_AWREADY[31];
            assign ap_WDATA[31][M_AXIMM_31_DATA_WIDTH-1:0] = AP_AXIMM_31_WDATA;
            assign ap_WSTRB[31][M_AXIMM_31_DATA_WIDTH/8-1:0] = AP_AXIMM_31_WSTRB;
            assign ap_WLAST[31] = AP_AXIMM_31_WLAST;
            assign ap_WVALID[31] = AP_AXIMM_31_WVALID;
            assign AP_AXIMM_31_WREADY = ap_WREADY[31];
            assign AP_AXIMM_31_BRESP = ap_BRESP[31];
            assign AP_AXIMM_31_BVALID = ap_BVALID[31];
            assign ap_BREADY[31] = AP_AXIMM_31_BREADY;
            assign ap_ARADDR[31][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_31_ARADDR;
            assign ap_ARLEN[31] = AP_AXIMM_31_ARLEN;
            assign ap_ARSIZE[31] = AP_AXIMM_31_ARSIZE;
            assign ap_ARBURST[31] = AP_AXIMM_31_ARBURST;
            assign ap_ARLOCK[31] = AP_AXIMM_31_ARLOCK;
            assign ap_ARCACHE[31] = AP_AXIMM_31_ARCACHE;
            assign ap_ARPROT[31] = AP_AXIMM_31_ARPROT;
            assign ap_ARREGION[31] = AP_AXIMM_31_ARREGION;
            assign ap_ARQOS[31] = AP_AXIMM_31_ARQOS;
            assign ap_ARVALID[31] = AP_AXIMM_31_ARVALID;
            assign AP_AXIMM_31_ARREADY = ap_ARREADY[31];
            assign AP_AXIMM_31_RDATA = ap_RDATA[31][M_AXIMM_31_DATA_WIDTH-1:0];
            assign AP_AXIMM_31_RRESP = ap_RRESP[31];
            assign AP_AXIMM_31_RLAST = ap_RLAST[31];
            assign AP_AXIMM_31_RVALID = ap_RVALID[31];
            assign ap_RREADY[31] = AP_AXIMM_31_RREADY;
            assign M_AXIMM_31_AWADDR = dm_AWADDR[31][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_31_AWLEN = dm_AWLEN[31];
            assign M_AXIMM_31_AWSIZE = dm_AWSIZE[31];
            assign M_AXIMM_31_AWBURST = dm_AWBURST[31];
            assign M_AXIMM_31_AWLOCK = dm_AWLOCK[31];
            assign M_AXIMM_31_AWCACHE = dm_AWCACHE[31];
            assign M_AXIMM_31_AWPROT = dm_AWPROT[31];
            assign M_AXIMM_31_AWREGION = dm_AWREGION[31];
            assign M_AXIMM_31_AWQOS = dm_AWQOS[31];
            assign M_AXIMM_31_AWVALID = dm_AWVALID[31];
            assign dm_AWREADY[31] = M_AXIMM_31_AWREADY;
            assign M_AXIMM_31_WDATA = dm_WDATA[31][M_AXIMM_31_DATA_WIDTH-1:0];
            assign M_AXIMM_31_WSTRB = dm_WSTRB[31][M_AXIMM_31_DATA_WIDTH/8-1:0];
            assign M_AXIMM_31_WLAST = dm_WLAST[31];
            assign M_AXIMM_31_WVALID = dm_WVALID[31];
            assign dm_WREADY[31] = M_AXIMM_31_WREADY;
            assign dm_BRESP[31] = M_AXIMM_31_BRESP;
            assign dm_BVALID[31] = M_AXIMM_31_BVALID;
            assign M_AXIMM_31_BREADY = dm_BREADY[31];
            assign M_AXIMM_31_ARADDR = dm_ARADDR[31][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_31_ARLEN = dm_ARLEN[31];
            assign M_AXIMM_31_ARSIZE = dm_ARSIZE[31];
            assign M_AXIMM_31_ARBURST = dm_ARBURST[31];
            assign M_AXIMM_31_ARLOCK = dm_ARLOCK[31];
            assign M_AXIMM_31_ARCACHE = dm_ARCACHE[31];
            assign M_AXIMM_31_ARPROT = dm_ARPROT[31];
            assign M_AXIMM_31_ARREGION = dm_ARREGION[31];
            assign M_AXIMM_31_ARQOS = dm_ARQOS[31];
            assign M_AXIMM_31_ARVALID = dm_ARVALID[31];
            assign dm_ARREADY[31] = M_AXIMM_31_ARREADY;
            assign dm_RDATA[31][M_AXIMM_31_DATA_WIDTH-1:0] = M_AXIMM_31_RDATA;
            assign dm_RRESP[31] = M_AXIMM_31_RRESP;
            assign dm_RLAST[31] = M_AXIMM_31_RLAST;
            assign dm_RVALID[31] = M_AXIMM_31_RVALID;
            assign M_AXIMM_31_RREADY = dm_RREADY[31];
        end
        if(C_NUM_AXIMMs > 32) begin
            assign ap_AWADDR[32][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_32_AWADDR;
            assign ap_AWLEN[32] = AP_AXIMM_32_AWLEN;
            assign ap_AWSIZE[32] = AP_AXIMM_32_AWSIZE;
            assign ap_AWBURST[32] = AP_AXIMM_32_AWBURST;
            assign ap_AWLOCK[32] = AP_AXIMM_32_AWLOCK;
            assign ap_AWCACHE[32] = AP_AXIMM_32_AWCACHE;
            assign ap_AWPROT[32] = AP_AXIMM_32_AWPROT;
            assign ap_AWREGION[32] = AP_AXIMM_32_AWREGION;
            assign ap_AWQOS[32] = AP_AXIMM_32_AWQOS;
            assign ap_AWVALID[32] = AP_AXIMM_32_AWVALID;
            assign AP_AXIMM_32_AWREADY = ap_AWREADY[32];
            assign ap_WDATA[32][M_AXIMM_32_DATA_WIDTH-1:0] = AP_AXIMM_32_WDATA;
            assign ap_WSTRB[32][M_AXIMM_32_DATA_WIDTH/8-1:0] = AP_AXIMM_32_WSTRB;
            assign ap_WLAST[32] = AP_AXIMM_32_WLAST;
            assign ap_WVALID[32] = AP_AXIMM_32_WVALID;
            assign AP_AXIMM_32_WREADY = ap_WREADY[32];
            assign AP_AXIMM_32_BRESP = ap_BRESP[32];
            assign AP_AXIMM_32_BVALID = ap_BVALID[32];
            assign ap_BREADY[32] = AP_AXIMM_32_BREADY;
            assign ap_ARADDR[32][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_32_ARADDR;
            assign ap_ARLEN[32] = AP_AXIMM_32_ARLEN;
            assign ap_ARSIZE[32] = AP_AXIMM_32_ARSIZE;
            assign ap_ARBURST[32] = AP_AXIMM_32_ARBURST;
            assign ap_ARLOCK[32] = AP_AXIMM_32_ARLOCK;
            assign ap_ARCACHE[32] = AP_AXIMM_32_ARCACHE;
            assign ap_ARPROT[32] = AP_AXIMM_32_ARPROT;
            assign ap_ARREGION[32] = AP_AXIMM_32_ARREGION;
            assign ap_ARQOS[32] = AP_AXIMM_32_ARQOS;
            assign ap_ARVALID[32] = AP_AXIMM_32_ARVALID;
            assign AP_AXIMM_32_ARREADY = ap_ARREADY[32];
            assign AP_AXIMM_32_RDATA = ap_RDATA[32][M_AXIMM_32_DATA_WIDTH-1:0];
            assign AP_AXIMM_32_RRESP = ap_RRESP[32];
            assign AP_AXIMM_32_RLAST = ap_RLAST[32];
            assign AP_AXIMM_32_RVALID = ap_RVALID[32];
            assign ap_RREADY[32] = AP_AXIMM_32_RREADY;
            assign M_AXIMM_32_AWADDR = dm_AWADDR[32][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_32_AWLEN = dm_AWLEN[32];
            assign M_AXIMM_32_AWSIZE = dm_AWSIZE[32];
            assign M_AXIMM_32_AWBURST = dm_AWBURST[32];
            assign M_AXIMM_32_AWLOCK = dm_AWLOCK[32];
            assign M_AXIMM_32_AWCACHE = dm_AWCACHE[32];
            assign M_AXIMM_32_AWPROT = dm_AWPROT[32];
            assign M_AXIMM_32_AWREGION = dm_AWREGION[32];
            assign M_AXIMM_32_AWQOS = dm_AWQOS[32];
            assign M_AXIMM_32_AWVALID = dm_AWVALID[32];
            assign dm_AWREADY[32] = M_AXIMM_32_AWREADY;
            assign M_AXIMM_32_WDATA = dm_WDATA[32][M_AXIMM_32_DATA_WIDTH-1:0];
            assign M_AXIMM_32_WSTRB = dm_WSTRB[32][M_AXIMM_32_DATA_WIDTH/8-1:0];
            assign M_AXIMM_32_WLAST = dm_WLAST[32];
            assign M_AXIMM_32_WVALID = dm_WVALID[32];
            assign dm_WREADY[32] = M_AXIMM_32_WREADY;
            assign dm_BRESP[32] = M_AXIMM_32_BRESP;
            assign dm_BVALID[32] = M_AXIMM_32_BVALID;
            assign M_AXIMM_32_BREADY = dm_BREADY[32];
            assign M_AXIMM_32_ARADDR = dm_ARADDR[32][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_32_ARLEN = dm_ARLEN[32];
            assign M_AXIMM_32_ARSIZE = dm_ARSIZE[32];
            assign M_AXIMM_32_ARBURST = dm_ARBURST[32];
            assign M_AXIMM_32_ARLOCK = dm_ARLOCK[32];
            assign M_AXIMM_32_ARCACHE = dm_ARCACHE[32];
            assign M_AXIMM_32_ARPROT = dm_ARPROT[32];
            assign M_AXIMM_32_ARREGION = dm_ARREGION[32];
            assign M_AXIMM_32_ARQOS = dm_ARQOS[32];
            assign M_AXIMM_32_ARVALID = dm_ARVALID[32];
            assign dm_ARREADY[32] = M_AXIMM_32_ARREADY;
            assign dm_RDATA[32][M_AXIMM_32_DATA_WIDTH-1:0] = M_AXIMM_32_RDATA;
            assign dm_RRESP[32] = M_AXIMM_32_RRESP;
            assign dm_RLAST[32] = M_AXIMM_32_RLAST;
            assign dm_RVALID[32] = M_AXIMM_32_RVALID;
            assign M_AXIMM_32_RREADY = dm_RREADY[32];
        end
        if(C_NUM_AXIMMs > 33) begin
            assign ap_AWADDR[33][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_33_AWADDR;
            assign ap_AWLEN[33] = AP_AXIMM_33_AWLEN;
            assign ap_AWSIZE[33] = AP_AXIMM_33_AWSIZE;
            assign ap_AWBURST[33] = AP_AXIMM_33_AWBURST;
            assign ap_AWLOCK[33] = AP_AXIMM_33_AWLOCK;
            assign ap_AWCACHE[33] = AP_AXIMM_33_AWCACHE;
            assign ap_AWPROT[33] = AP_AXIMM_33_AWPROT;
            assign ap_AWREGION[33] = AP_AXIMM_33_AWREGION;
            assign ap_AWQOS[33] = AP_AXIMM_33_AWQOS;
            assign ap_AWVALID[33] = AP_AXIMM_33_AWVALID;
            assign AP_AXIMM_33_AWREADY = ap_AWREADY[33];
            assign ap_WDATA[33][M_AXIMM_33_DATA_WIDTH-1:0] = AP_AXIMM_33_WDATA;
            assign ap_WSTRB[33][M_AXIMM_33_DATA_WIDTH/8-1:0] = AP_AXIMM_33_WSTRB;
            assign ap_WLAST[33] = AP_AXIMM_33_WLAST;
            assign ap_WVALID[33] = AP_AXIMM_33_WVALID;
            assign AP_AXIMM_33_WREADY = ap_WREADY[33];
            assign AP_AXIMM_33_BRESP = ap_BRESP[33];
            assign AP_AXIMM_33_BVALID = ap_BVALID[33];
            assign ap_BREADY[33] = AP_AXIMM_33_BREADY;
            assign ap_ARADDR[33][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_33_ARADDR;
            assign ap_ARLEN[33] = AP_AXIMM_33_ARLEN;
            assign ap_ARSIZE[33] = AP_AXIMM_33_ARSIZE;
            assign ap_ARBURST[33] = AP_AXIMM_33_ARBURST;
            assign ap_ARLOCK[33] = AP_AXIMM_33_ARLOCK;
            assign ap_ARCACHE[33] = AP_AXIMM_33_ARCACHE;
            assign ap_ARPROT[33] = AP_AXIMM_33_ARPROT;
            assign ap_ARREGION[33] = AP_AXIMM_33_ARREGION;
            assign ap_ARQOS[33] = AP_AXIMM_33_ARQOS;
            assign ap_ARVALID[33] = AP_AXIMM_33_ARVALID;
            assign AP_AXIMM_33_ARREADY = ap_ARREADY[33];
            assign AP_AXIMM_33_RDATA = ap_RDATA[33][M_AXIMM_33_DATA_WIDTH-1:0];
            assign AP_AXIMM_33_RRESP = ap_RRESP[33];
            assign AP_AXIMM_33_RLAST = ap_RLAST[33];
            assign AP_AXIMM_33_RVALID = ap_RVALID[33];
            assign ap_RREADY[33] = AP_AXIMM_33_RREADY;
            assign M_AXIMM_33_AWADDR = dm_AWADDR[33][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_33_AWLEN = dm_AWLEN[33];
            assign M_AXIMM_33_AWSIZE = dm_AWSIZE[33];
            assign M_AXIMM_33_AWBURST = dm_AWBURST[33];
            assign M_AXIMM_33_AWLOCK = dm_AWLOCK[33];
            assign M_AXIMM_33_AWCACHE = dm_AWCACHE[33];
            assign M_AXIMM_33_AWPROT = dm_AWPROT[33];
            assign M_AXIMM_33_AWREGION = dm_AWREGION[33];
            assign M_AXIMM_33_AWQOS = dm_AWQOS[33];
            assign M_AXIMM_33_AWVALID = dm_AWVALID[33];
            assign dm_AWREADY[33] = M_AXIMM_33_AWREADY;
            assign M_AXIMM_33_WDATA = dm_WDATA[33][M_AXIMM_33_DATA_WIDTH-1:0];
            assign M_AXIMM_33_WSTRB = dm_WSTRB[33][M_AXIMM_33_DATA_WIDTH/8-1:0];
            assign M_AXIMM_33_WLAST = dm_WLAST[33];
            assign M_AXIMM_33_WVALID = dm_WVALID[33];
            assign dm_WREADY[33] = M_AXIMM_33_WREADY;
            assign dm_BRESP[33] = M_AXIMM_33_BRESP;
            assign dm_BVALID[33] = M_AXIMM_33_BVALID;
            assign M_AXIMM_33_BREADY = dm_BREADY[33];
            assign M_AXIMM_33_ARADDR = dm_ARADDR[33][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_33_ARLEN = dm_ARLEN[33];
            assign M_AXIMM_33_ARSIZE = dm_ARSIZE[33];
            assign M_AXIMM_33_ARBURST = dm_ARBURST[33];
            assign M_AXIMM_33_ARLOCK = dm_ARLOCK[33];
            assign M_AXIMM_33_ARCACHE = dm_ARCACHE[33];
            assign M_AXIMM_33_ARPROT = dm_ARPROT[33];
            assign M_AXIMM_33_ARREGION = dm_ARREGION[33];
            assign M_AXIMM_33_ARQOS = dm_ARQOS[33];
            assign M_AXIMM_33_ARVALID = dm_ARVALID[33];
            assign dm_ARREADY[33] = M_AXIMM_33_ARREADY;
            assign dm_RDATA[33][M_AXIMM_33_DATA_WIDTH-1:0] = M_AXIMM_33_RDATA;
            assign dm_RRESP[33] = M_AXIMM_33_RRESP;
            assign dm_RLAST[33] = M_AXIMM_33_RLAST;
            assign dm_RVALID[33] = M_AXIMM_33_RVALID;
            assign M_AXIMM_33_RREADY = dm_RREADY[33];
        end
        if(C_NUM_AXIMMs > 34) begin
            assign ap_AWADDR[34][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_34_AWADDR;
            assign ap_AWLEN[34] = AP_AXIMM_34_AWLEN;
            assign ap_AWSIZE[34] = AP_AXIMM_34_AWSIZE;
            assign ap_AWBURST[34] = AP_AXIMM_34_AWBURST;
            assign ap_AWLOCK[34] = AP_AXIMM_34_AWLOCK;
            assign ap_AWCACHE[34] = AP_AXIMM_34_AWCACHE;
            assign ap_AWPROT[34] = AP_AXIMM_34_AWPROT;
            assign ap_AWREGION[34] = AP_AXIMM_34_AWREGION;
            assign ap_AWQOS[34] = AP_AXIMM_34_AWQOS;
            assign ap_AWVALID[34] = AP_AXIMM_34_AWVALID;
            assign AP_AXIMM_34_AWREADY = ap_AWREADY[34];
            assign ap_WDATA[34][M_AXIMM_34_DATA_WIDTH-1:0] = AP_AXIMM_34_WDATA;
            assign ap_WSTRB[34][M_AXIMM_34_DATA_WIDTH/8-1:0] = AP_AXIMM_34_WSTRB;
            assign ap_WLAST[34] = AP_AXIMM_34_WLAST;
            assign ap_WVALID[34] = AP_AXIMM_34_WVALID;
            assign AP_AXIMM_34_WREADY = ap_WREADY[34];
            assign AP_AXIMM_34_BRESP = ap_BRESP[34];
            assign AP_AXIMM_34_BVALID = ap_BVALID[34];
            assign ap_BREADY[34] = AP_AXIMM_34_BREADY;
            assign ap_ARADDR[34][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_34_ARADDR;
            assign ap_ARLEN[34] = AP_AXIMM_34_ARLEN;
            assign ap_ARSIZE[34] = AP_AXIMM_34_ARSIZE;
            assign ap_ARBURST[34] = AP_AXIMM_34_ARBURST;
            assign ap_ARLOCK[34] = AP_AXIMM_34_ARLOCK;
            assign ap_ARCACHE[34] = AP_AXIMM_34_ARCACHE;
            assign ap_ARPROT[34] = AP_AXIMM_34_ARPROT;
            assign ap_ARREGION[34] = AP_AXIMM_34_ARREGION;
            assign ap_ARQOS[34] = AP_AXIMM_34_ARQOS;
            assign ap_ARVALID[34] = AP_AXIMM_34_ARVALID;
            assign AP_AXIMM_34_ARREADY = ap_ARREADY[34];
            assign AP_AXIMM_34_RDATA = ap_RDATA[34][M_AXIMM_34_DATA_WIDTH-1:0];
            assign AP_AXIMM_34_RRESP = ap_RRESP[34];
            assign AP_AXIMM_34_RLAST = ap_RLAST[34];
            assign AP_AXIMM_34_RVALID = ap_RVALID[34];
            assign ap_RREADY[34] = AP_AXIMM_34_RREADY;
            assign M_AXIMM_34_AWADDR = dm_AWADDR[34][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_34_AWLEN = dm_AWLEN[34];
            assign M_AXIMM_34_AWSIZE = dm_AWSIZE[34];
            assign M_AXIMM_34_AWBURST = dm_AWBURST[34];
            assign M_AXIMM_34_AWLOCK = dm_AWLOCK[34];
            assign M_AXIMM_34_AWCACHE = dm_AWCACHE[34];
            assign M_AXIMM_34_AWPROT = dm_AWPROT[34];
            assign M_AXIMM_34_AWREGION = dm_AWREGION[34];
            assign M_AXIMM_34_AWQOS = dm_AWQOS[34];
            assign M_AXIMM_34_AWVALID = dm_AWVALID[34];
            assign dm_AWREADY[34] = M_AXIMM_34_AWREADY;
            assign M_AXIMM_34_WDATA = dm_WDATA[34][M_AXIMM_34_DATA_WIDTH-1:0];
            assign M_AXIMM_34_WSTRB = dm_WSTRB[34][M_AXIMM_34_DATA_WIDTH/8-1:0];
            assign M_AXIMM_34_WLAST = dm_WLAST[34];
            assign M_AXIMM_34_WVALID = dm_WVALID[34];
            assign dm_WREADY[34] = M_AXIMM_34_WREADY;
            assign dm_BRESP[34] = M_AXIMM_34_BRESP;
            assign dm_BVALID[34] = M_AXIMM_34_BVALID;
            assign M_AXIMM_34_BREADY = dm_BREADY[34];
            assign M_AXIMM_34_ARADDR = dm_ARADDR[34][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_34_ARLEN = dm_ARLEN[34];
            assign M_AXIMM_34_ARSIZE = dm_ARSIZE[34];
            assign M_AXIMM_34_ARBURST = dm_ARBURST[34];
            assign M_AXIMM_34_ARLOCK = dm_ARLOCK[34];
            assign M_AXIMM_34_ARCACHE = dm_ARCACHE[34];
            assign M_AXIMM_34_ARPROT = dm_ARPROT[34];
            assign M_AXIMM_34_ARREGION = dm_ARREGION[34];
            assign M_AXIMM_34_ARQOS = dm_ARQOS[34];
            assign M_AXIMM_34_ARVALID = dm_ARVALID[34];
            assign dm_ARREADY[34] = M_AXIMM_34_ARREADY;
            assign dm_RDATA[34][M_AXIMM_34_DATA_WIDTH-1:0] = M_AXIMM_34_RDATA;
            assign dm_RRESP[34] = M_AXIMM_34_RRESP;
            assign dm_RLAST[34] = M_AXIMM_34_RLAST;
            assign dm_RVALID[34] = M_AXIMM_34_RVALID;
            assign M_AXIMM_34_RREADY = dm_RREADY[34];
        end
        if(C_NUM_AXIMMs > 35) begin
            assign ap_AWADDR[35][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_35_AWADDR;
            assign ap_AWLEN[35] = AP_AXIMM_35_AWLEN;
            assign ap_AWSIZE[35] = AP_AXIMM_35_AWSIZE;
            assign ap_AWBURST[35] = AP_AXIMM_35_AWBURST;
            assign ap_AWLOCK[35] = AP_AXIMM_35_AWLOCK;
            assign ap_AWCACHE[35] = AP_AXIMM_35_AWCACHE;
            assign ap_AWPROT[35] = AP_AXIMM_35_AWPROT;
            assign ap_AWREGION[35] = AP_AXIMM_35_AWREGION;
            assign ap_AWQOS[35] = AP_AXIMM_35_AWQOS;
            assign ap_AWVALID[35] = AP_AXIMM_35_AWVALID;
            assign AP_AXIMM_35_AWREADY = ap_AWREADY[35];
            assign ap_WDATA[35][M_AXIMM_35_DATA_WIDTH-1:0] = AP_AXIMM_35_WDATA;
            assign ap_WSTRB[35][M_AXIMM_35_DATA_WIDTH/8-1:0] = AP_AXIMM_35_WSTRB;
            assign ap_WLAST[35] = AP_AXIMM_35_WLAST;
            assign ap_WVALID[35] = AP_AXIMM_35_WVALID;
            assign AP_AXIMM_35_WREADY = ap_WREADY[35];
            assign AP_AXIMM_35_BRESP = ap_BRESP[35];
            assign AP_AXIMM_35_BVALID = ap_BVALID[35];
            assign ap_BREADY[35] = AP_AXIMM_35_BREADY;
            assign ap_ARADDR[35][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_35_ARADDR;
            assign ap_ARLEN[35] = AP_AXIMM_35_ARLEN;
            assign ap_ARSIZE[35] = AP_AXIMM_35_ARSIZE;
            assign ap_ARBURST[35] = AP_AXIMM_35_ARBURST;
            assign ap_ARLOCK[35] = AP_AXIMM_35_ARLOCK;
            assign ap_ARCACHE[35] = AP_AXIMM_35_ARCACHE;
            assign ap_ARPROT[35] = AP_AXIMM_35_ARPROT;
            assign ap_ARREGION[35] = AP_AXIMM_35_ARREGION;
            assign ap_ARQOS[35] = AP_AXIMM_35_ARQOS;
            assign ap_ARVALID[35] = AP_AXIMM_35_ARVALID;
            assign AP_AXIMM_35_ARREADY = ap_ARREADY[35];
            assign AP_AXIMM_35_RDATA = ap_RDATA[35][M_AXIMM_35_DATA_WIDTH-1:0];
            assign AP_AXIMM_35_RRESP = ap_RRESP[35];
            assign AP_AXIMM_35_RLAST = ap_RLAST[35];
            assign AP_AXIMM_35_RVALID = ap_RVALID[35];
            assign ap_RREADY[35] = AP_AXIMM_35_RREADY;
            assign M_AXIMM_35_AWADDR = dm_AWADDR[35][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_35_AWLEN = dm_AWLEN[35];
            assign M_AXIMM_35_AWSIZE = dm_AWSIZE[35];
            assign M_AXIMM_35_AWBURST = dm_AWBURST[35];
            assign M_AXIMM_35_AWLOCK = dm_AWLOCK[35];
            assign M_AXIMM_35_AWCACHE = dm_AWCACHE[35];
            assign M_AXIMM_35_AWPROT = dm_AWPROT[35];
            assign M_AXIMM_35_AWREGION = dm_AWREGION[35];
            assign M_AXIMM_35_AWQOS = dm_AWQOS[35];
            assign M_AXIMM_35_AWVALID = dm_AWVALID[35];
            assign dm_AWREADY[35] = M_AXIMM_35_AWREADY;
            assign M_AXIMM_35_WDATA = dm_WDATA[35][M_AXIMM_35_DATA_WIDTH-1:0];
            assign M_AXIMM_35_WSTRB = dm_WSTRB[35][M_AXIMM_35_DATA_WIDTH/8-1:0];
            assign M_AXIMM_35_WLAST = dm_WLAST[35];
            assign M_AXIMM_35_WVALID = dm_WVALID[35];
            assign dm_WREADY[35] = M_AXIMM_35_WREADY;
            assign dm_BRESP[35] = M_AXIMM_35_BRESP;
            assign dm_BVALID[35] = M_AXIMM_35_BVALID;
            assign M_AXIMM_35_BREADY = dm_BREADY[35];
            assign M_AXIMM_35_ARADDR = dm_ARADDR[35][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_35_ARLEN = dm_ARLEN[35];
            assign M_AXIMM_35_ARSIZE = dm_ARSIZE[35];
            assign M_AXIMM_35_ARBURST = dm_ARBURST[35];
            assign M_AXIMM_35_ARLOCK = dm_ARLOCK[35];
            assign M_AXIMM_35_ARCACHE = dm_ARCACHE[35];
            assign M_AXIMM_35_ARPROT = dm_ARPROT[35];
            assign M_AXIMM_35_ARREGION = dm_ARREGION[35];
            assign M_AXIMM_35_ARQOS = dm_ARQOS[35];
            assign M_AXIMM_35_ARVALID = dm_ARVALID[35];
            assign dm_ARREADY[35] = M_AXIMM_35_ARREADY;
            assign dm_RDATA[35][M_AXIMM_35_DATA_WIDTH-1:0] = M_AXIMM_35_RDATA;
            assign dm_RRESP[35] = M_AXIMM_35_RRESP;
            assign dm_RLAST[35] = M_AXIMM_35_RLAST;
            assign dm_RVALID[35] = M_AXIMM_35_RVALID;
            assign M_AXIMM_35_RREADY = dm_RREADY[35];
        end
        if(C_NUM_AXIMMs > 36) begin
            assign ap_AWADDR[36][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_36_AWADDR;
            assign ap_AWLEN[36] = AP_AXIMM_36_AWLEN;
            assign ap_AWSIZE[36] = AP_AXIMM_36_AWSIZE;
            assign ap_AWBURST[36] = AP_AXIMM_36_AWBURST;
            assign ap_AWLOCK[36] = AP_AXIMM_36_AWLOCK;
            assign ap_AWCACHE[36] = AP_AXIMM_36_AWCACHE;
            assign ap_AWPROT[36] = AP_AXIMM_36_AWPROT;
            assign ap_AWREGION[36] = AP_AXIMM_36_AWREGION;
            assign ap_AWQOS[36] = AP_AXIMM_36_AWQOS;
            assign ap_AWVALID[36] = AP_AXIMM_36_AWVALID;
            assign AP_AXIMM_36_AWREADY = ap_AWREADY[36];
            assign ap_WDATA[36][M_AXIMM_36_DATA_WIDTH-1:0] = AP_AXIMM_36_WDATA;
            assign ap_WSTRB[36][M_AXIMM_36_DATA_WIDTH/8-1:0] = AP_AXIMM_36_WSTRB;
            assign ap_WLAST[36] = AP_AXIMM_36_WLAST;
            assign ap_WVALID[36] = AP_AXIMM_36_WVALID;
            assign AP_AXIMM_36_WREADY = ap_WREADY[36];
            assign AP_AXIMM_36_BRESP = ap_BRESP[36];
            assign AP_AXIMM_36_BVALID = ap_BVALID[36];
            assign ap_BREADY[36] = AP_AXIMM_36_BREADY;
            assign ap_ARADDR[36][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_36_ARADDR;
            assign ap_ARLEN[36] = AP_AXIMM_36_ARLEN;
            assign ap_ARSIZE[36] = AP_AXIMM_36_ARSIZE;
            assign ap_ARBURST[36] = AP_AXIMM_36_ARBURST;
            assign ap_ARLOCK[36] = AP_AXIMM_36_ARLOCK;
            assign ap_ARCACHE[36] = AP_AXIMM_36_ARCACHE;
            assign ap_ARPROT[36] = AP_AXIMM_36_ARPROT;
            assign ap_ARREGION[36] = AP_AXIMM_36_ARREGION;
            assign ap_ARQOS[36] = AP_AXIMM_36_ARQOS;
            assign ap_ARVALID[36] = AP_AXIMM_36_ARVALID;
            assign AP_AXIMM_36_ARREADY = ap_ARREADY[36];
            assign AP_AXIMM_36_RDATA = ap_RDATA[36][M_AXIMM_36_DATA_WIDTH-1:0];
            assign AP_AXIMM_36_RRESP = ap_RRESP[36];
            assign AP_AXIMM_36_RLAST = ap_RLAST[36];
            assign AP_AXIMM_36_RVALID = ap_RVALID[36];
            assign ap_RREADY[36] = AP_AXIMM_36_RREADY;
            assign M_AXIMM_36_AWADDR = dm_AWADDR[36][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_36_AWLEN = dm_AWLEN[36];
            assign M_AXIMM_36_AWSIZE = dm_AWSIZE[36];
            assign M_AXIMM_36_AWBURST = dm_AWBURST[36];
            assign M_AXIMM_36_AWLOCK = dm_AWLOCK[36];
            assign M_AXIMM_36_AWCACHE = dm_AWCACHE[36];
            assign M_AXIMM_36_AWPROT = dm_AWPROT[36];
            assign M_AXIMM_36_AWREGION = dm_AWREGION[36];
            assign M_AXIMM_36_AWQOS = dm_AWQOS[36];
            assign M_AXIMM_36_AWVALID = dm_AWVALID[36];
            assign dm_AWREADY[36] = M_AXIMM_36_AWREADY;
            assign M_AXIMM_36_WDATA = dm_WDATA[36][M_AXIMM_36_DATA_WIDTH-1:0];
            assign M_AXIMM_36_WSTRB = dm_WSTRB[36][M_AXIMM_36_DATA_WIDTH/8-1:0];
            assign M_AXIMM_36_WLAST = dm_WLAST[36];
            assign M_AXIMM_36_WVALID = dm_WVALID[36];
            assign dm_WREADY[36] = M_AXIMM_36_WREADY;
            assign dm_BRESP[36] = M_AXIMM_36_BRESP;
            assign dm_BVALID[36] = M_AXIMM_36_BVALID;
            assign M_AXIMM_36_BREADY = dm_BREADY[36];
            assign M_AXIMM_36_ARADDR = dm_ARADDR[36][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_36_ARLEN = dm_ARLEN[36];
            assign M_AXIMM_36_ARSIZE = dm_ARSIZE[36];
            assign M_AXIMM_36_ARBURST = dm_ARBURST[36];
            assign M_AXIMM_36_ARLOCK = dm_ARLOCK[36];
            assign M_AXIMM_36_ARCACHE = dm_ARCACHE[36];
            assign M_AXIMM_36_ARPROT = dm_ARPROT[36];
            assign M_AXIMM_36_ARREGION = dm_ARREGION[36];
            assign M_AXIMM_36_ARQOS = dm_ARQOS[36];
            assign M_AXIMM_36_ARVALID = dm_ARVALID[36];
            assign dm_ARREADY[36] = M_AXIMM_36_ARREADY;
            assign dm_RDATA[36][M_AXIMM_36_DATA_WIDTH-1:0] = M_AXIMM_36_RDATA;
            assign dm_RRESP[36] = M_AXIMM_36_RRESP;
            assign dm_RLAST[36] = M_AXIMM_36_RLAST;
            assign dm_RVALID[36] = M_AXIMM_36_RVALID;
            assign M_AXIMM_36_RREADY = dm_RREADY[36];
        end
        if(C_NUM_AXIMMs > 37) begin
            assign ap_AWADDR[37][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_37_AWADDR;
            assign ap_AWLEN[37] = AP_AXIMM_37_AWLEN;
            assign ap_AWSIZE[37] = AP_AXIMM_37_AWSIZE;
            assign ap_AWBURST[37] = AP_AXIMM_37_AWBURST;
            assign ap_AWLOCK[37] = AP_AXIMM_37_AWLOCK;
            assign ap_AWCACHE[37] = AP_AXIMM_37_AWCACHE;
            assign ap_AWPROT[37] = AP_AXIMM_37_AWPROT;
            assign ap_AWREGION[37] = AP_AXIMM_37_AWREGION;
            assign ap_AWQOS[37] = AP_AXIMM_37_AWQOS;
            assign ap_AWVALID[37] = AP_AXIMM_37_AWVALID;
            assign AP_AXIMM_37_AWREADY = ap_AWREADY[37];
            assign ap_WDATA[37][M_AXIMM_37_DATA_WIDTH-1:0] = AP_AXIMM_37_WDATA;
            assign ap_WSTRB[37][M_AXIMM_37_DATA_WIDTH/8-1:0] = AP_AXIMM_37_WSTRB;
            assign ap_WLAST[37] = AP_AXIMM_37_WLAST;
            assign ap_WVALID[37] = AP_AXIMM_37_WVALID;
            assign AP_AXIMM_37_WREADY = ap_WREADY[37];
            assign AP_AXIMM_37_BRESP = ap_BRESP[37];
            assign AP_AXIMM_37_BVALID = ap_BVALID[37];
            assign ap_BREADY[37] = AP_AXIMM_37_BREADY;
            assign ap_ARADDR[37][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_37_ARADDR;
            assign ap_ARLEN[37] = AP_AXIMM_37_ARLEN;
            assign ap_ARSIZE[37] = AP_AXIMM_37_ARSIZE;
            assign ap_ARBURST[37] = AP_AXIMM_37_ARBURST;
            assign ap_ARLOCK[37] = AP_AXIMM_37_ARLOCK;
            assign ap_ARCACHE[37] = AP_AXIMM_37_ARCACHE;
            assign ap_ARPROT[37] = AP_AXIMM_37_ARPROT;
            assign ap_ARREGION[37] = AP_AXIMM_37_ARREGION;
            assign ap_ARQOS[37] = AP_AXIMM_37_ARQOS;
            assign ap_ARVALID[37] = AP_AXIMM_37_ARVALID;
            assign AP_AXIMM_37_ARREADY = ap_ARREADY[37];
            assign AP_AXIMM_37_RDATA = ap_RDATA[37][M_AXIMM_37_DATA_WIDTH-1:0];
            assign AP_AXIMM_37_RRESP = ap_RRESP[37];
            assign AP_AXIMM_37_RLAST = ap_RLAST[37];
            assign AP_AXIMM_37_RVALID = ap_RVALID[37];
            assign ap_RREADY[37] = AP_AXIMM_37_RREADY;
            assign M_AXIMM_37_AWADDR = dm_AWADDR[37][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_37_AWLEN = dm_AWLEN[37];
            assign M_AXIMM_37_AWSIZE = dm_AWSIZE[37];
            assign M_AXIMM_37_AWBURST = dm_AWBURST[37];
            assign M_AXIMM_37_AWLOCK = dm_AWLOCK[37];
            assign M_AXIMM_37_AWCACHE = dm_AWCACHE[37];
            assign M_AXIMM_37_AWPROT = dm_AWPROT[37];
            assign M_AXIMM_37_AWREGION = dm_AWREGION[37];
            assign M_AXIMM_37_AWQOS = dm_AWQOS[37];
            assign M_AXIMM_37_AWVALID = dm_AWVALID[37];
            assign dm_AWREADY[37] = M_AXIMM_37_AWREADY;
            assign M_AXIMM_37_WDATA = dm_WDATA[37][M_AXIMM_37_DATA_WIDTH-1:0];
            assign M_AXIMM_37_WSTRB = dm_WSTRB[37][M_AXIMM_37_DATA_WIDTH/8-1:0];
            assign M_AXIMM_37_WLAST = dm_WLAST[37];
            assign M_AXIMM_37_WVALID = dm_WVALID[37];
            assign dm_WREADY[37] = M_AXIMM_37_WREADY;
            assign dm_BRESP[37] = M_AXIMM_37_BRESP;
            assign dm_BVALID[37] = M_AXIMM_37_BVALID;
            assign M_AXIMM_37_BREADY = dm_BREADY[37];
            assign M_AXIMM_37_ARADDR = dm_ARADDR[37][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_37_ARLEN = dm_ARLEN[37];
            assign M_AXIMM_37_ARSIZE = dm_ARSIZE[37];
            assign M_AXIMM_37_ARBURST = dm_ARBURST[37];
            assign M_AXIMM_37_ARLOCK = dm_ARLOCK[37];
            assign M_AXIMM_37_ARCACHE = dm_ARCACHE[37];
            assign M_AXIMM_37_ARPROT = dm_ARPROT[37];
            assign M_AXIMM_37_ARREGION = dm_ARREGION[37];
            assign M_AXIMM_37_ARQOS = dm_ARQOS[37];
            assign M_AXIMM_37_ARVALID = dm_ARVALID[37];
            assign dm_ARREADY[37] = M_AXIMM_37_ARREADY;
            assign dm_RDATA[37][M_AXIMM_37_DATA_WIDTH-1:0] = M_AXIMM_37_RDATA;
            assign dm_RRESP[37] = M_AXIMM_37_RRESP;
            assign dm_RLAST[37] = M_AXIMM_37_RLAST;
            assign dm_RVALID[37] = M_AXIMM_37_RVALID;
            assign M_AXIMM_37_RREADY = dm_RREADY[37];
        end
        if(C_NUM_AXIMMs > 38) begin
            assign ap_AWADDR[38][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_38_AWADDR;
            assign ap_AWLEN[38] = AP_AXIMM_38_AWLEN;
            assign ap_AWSIZE[38] = AP_AXIMM_38_AWSIZE;
            assign ap_AWBURST[38] = AP_AXIMM_38_AWBURST;
            assign ap_AWLOCK[38] = AP_AXIMM_38_AWLOCK;
            assign ap_AWCACHE[38] = AP_AXIMM_38_AWCACHE;
            assign ap_AWPROT[38] = AP_AXIMM_38_AWPROT;
            assign ap_AWREGION[38] = AP_AXIMM_38_AWREGION;
            assign ap_AWQOS[38] = AP_AXIMM_38_AWQOS;
            assign ap_AWVALID[38] = AP_AXIMM_38_AWVALID;
            assign AP_AXIMM_38_AWREADY = ap_AWREADY[38];
            assign ap_WDATA[38][M_AXIMM_38_DATA_WIDTH-1:0] = AP_AXIMM_38_WDATA;
            assign ap_WSTRB[38][M_AXIMM_38_DATA_WIDTH/8-1:0] = AP_AXIMM_38_WSTRB;
            assign ap_WLAST[38] = AP_AXIMM_38_WLAST;
            assign ap_WVALID[38] = AP_AXIMM_38_WVALID;
            assign AP_AXIMM_38_WREADY = ap_WREADY[38];
            assign AP_AXIMM_38_BRESP = ap_BRESP[38];
            assign AP_AXIMM_38_BVALID = ap_BVALID[38];
            assign ap_BREADY[38] = AP_AXIMM_38_BREADY;
            assign ap_ARADDR[38][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_38_ARADDR;
            assign ap_ARLEN[38] = AP_AXIMM_38_ARLEN;
            assign ap_ARSIZE[38] = AP_AXIMM_38_ARSIZE;
            assign ap_ARBURST[38] = AP_AXIMM_38_ARBURST;
            assign ap_ARLOCK[38] = AP_AXIMM_38_ARLOCK;
            assign ap_ARCACHE[38] = AP_AXIMM_38_ARCACHE;
            assign ap_ARPROT[38] = AP_AXIMM_38_ARPROT;
            assign ap_ARREGION[38] = AP_AXIMM_38_ARREGION;
            assign ap_ARQOS[38] = AP_AXIMM_38_ARQOS;
            assign ap_ARVALID[38] = AP_AXIMM_38_ARVALID;
            assign AP_AXIMM_38_ARREADY = ap_ARREADY[38];
            assign AP_AXIMM_38_RDATA = ap_RDATA[38][M_AXIMM_38_DATA_WIDTH-1:0];
            assign AP_AXIMM_38_RRESP = ap_RRESP[38];
            assign AP_AXIMM_38_RLAST = ap_RLAST[38];
            assign AP_AXIMM_38_RVALID = ap_RVALID[38];
            assign ap_RREADY[38] = AP_AXIMM_38_RREADY;
            assign M_AXIMM_38_AWADDR = dm_AWADDR[38][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_38_AWLEN = dm_AWLEN[38];
            assign M_AXIMM_38_AWSIZE = dm_AWSIZE[38];
            assign M_AXIMM_38_AWBURST = dm_AWBURST[38];
            assign M_AXIMM_38_AWLOCK = dm_AWLOCK[38];
            assign M_AXIMM_38_AWCACHE = dm_AWCACHE[38];
            assign M_AXIMM_38_AWPROT = dm_AWPROT[38];
            assign M_AXIMM_38_AWREGION = dm_AWREGION[38];
            assign M_AXIMM_38_AWQOS = dm_AWQOS[38];
            assign M_AXIMM_38_AWVALID = dm_AWVALID[38];
            assign dm_AWREADY[38] = M_AXIMM_38_AWREADY;
            assign M_AXIMM_38_WDATA = dm_WDATA[38][M_AXIMM_38_DATA_WIDTH-1:0];
            assign M_AXIMM_38_WSTRB = dm_WSTRB[38][M_AXIMM_38_DATA_WIDTH/8-1:0];
            assign M_AXIMM_38_WLAST = dm_WLAST[38];
            assign M_AXIMM_38_WVALID = dm_WVALID[38];
            assign dm_WREADY[38] = M_AXIMM_38_WREADY;
            assign dm_BRESP[38] = M_AXIMM_38_BRESP;
            assign dm_BVALID[38] = M_AXIMM_38_BVALID;
            assign M_AXIMM_38_BREADY = dm_BREADY[38];
            assign M_AXIMM_38_ARADDR = dm_ARADDR[38][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_38_ARLEN = dm_ARLEN[38];
            assign M_AXIMM_38_ARSIZE = dm_ARSIZE[38];
            assign M_AXIMM_38_ARBURST = dm_ARBURST[38];
            assign M_AXIMM_38_ARLOCK = dm_ARLOCK[38];
            assign M_AXIMM_38_ARCACHE = dm_ARCACHE[38];
            assign M_AXIMM_38_ARPROT = dm_ARPROT[38];
            assign M_AXIMM_38_ARREGION = dm_ARREGION[38];
            assign M_AXIMM_38_ARQOS = dm_ARQOS[38];
            assign M_AXIMM_38_ARVALID = dm_ARVALID[38];
            assign dm_ARREADY[38] = M_AXIMM_38_ARREADY;
            assign dm_RDATA[38][M_AXIMM_38_DATA_WIDTH-1:0] = M_AXIMM_38_RDATA;
            assign dm_RRESP[38] = M_AXIMM_38_RRESP;
            assign dm_RLAST[38] = M_AXIMM_38_RLAST;
            assign dm_RVALID[38] = M_AXIMM_38_RVALID;
            assign M_AXIMM_38_RREADY = dm_RREADY[38];
        end
        if(C_NUM_AXIMMs > 39) begin
            assign ap_AWADDR[39][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_39_AWADDR;
            assign ap_AWLEN[39] = AP_AXIMM_39_AWLEN;
            assign ap_AWSIZE[39] = AP_AXIMM_39_AWSIZE;
            assign ap_AWBURST[39] = AP_AXIMM_39_AWBURST;
            assign ap_AWLOCK[39] = AP_AXIMM_39_AWLOCK;
            assign ap_AWCACHE[39] = AP_AXIMM_39_AWCACHE;
            assign ap_AWPROT[39] = AP_AXIMM_39_AWPROT;
            assign ap_AWREGION[39] = AP_AXIMM_39_AWREGION;
            assign ap_AWQOS[39] = AP_AXIMM_39_AWQOS;
            assign ap_AWVALID[39] = AP_AXIMM_39_AWVALID;
            assign AP_AXIMM_39_AWREADY = ap_AWREADY[39];
            assign ap_WDATA[39][M_AXIMM_39_DATA_WIDTH-1:0] = AP_AXIMM_39_WDATA;
            assign ap_WSTRB[39][M_AXIMM_39_DATA_WIDTH/8-1:0] = AP_AXIMM_39_WSTRB;
            assign ap_WLAST[39] = AP_AXIMM_39_WLAST;
            assign ap_WVALID[39] = AP_AXIMM_39_WVALID;
            assign AP_AXIMM_39_WREADY = ap_WREADY[39];
            assign AP_AXIMM_39_BRESP = ap_BRESP[39];
            assign AP_AXIMM_39_BVALID = ap_BVALID[39];
            assign ap_BREADY[39] = AP_AXIMM_39_BREADY;
            assign ap_ARADDR[39][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_39_ARADDR;
            assign ap_ARLEN[39] = AP_AXIMM_39_ARLEN;
            assign ap_ARSIZE[39] = AP_AXIMM_39_ARSIZE;
            assign ap_ARBURST[39] = AP_AXIMM_39_ARBURST;
            assign ap_ARLOCK[39] = AP_AXIMM_39_ARLOCK;
            assign ap_ARCACHE[39] = AP_AXIMM_39_ARCACHE;
            assign ap_ARPROT[39] = AP_AXIMM_39_ARPROT;
            assign ap_ARREGION[39] = AP_AXIMM_39_ARREGION;
            assign ap_ARQOS[39] = AP_AXIMM_39_ARQOS;
            assign ap_ARVALID[39] = AP_AXIMM_39_ARVALID;
            assign AP_AXIMM_39_ARREADY = ap_ARREADY[39];
            assign AP_AXIMM_39_RDATA = ap_RDATA[39][M_AXIMM_39_DATA_WIDTH-1:0];
            assign AP_AXIMM_39_RRESP = ap_RRESP[39];
            assign AP_AXIMM_39_RLAST = ap_RLAST[39];
            assign AP_AXIMM_39_RVALID = ap_RVALID[39];
            assign ap_RREADY[39] = AP_AXIMM_39_RREADY;
            assign M_AXIMM_39_AWADDR = dm_AWADDR[39][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_39_AWLEN = dm_AWLEN[39];
            assign M_AXIMM_39_AWSIZE = dm_AWSIZE[39];
            assign M_AXIMM_39_AWBURST = dm_AWBURST[39];
            assign M_AXIMM_39_AWLOCK = dm_AWLOCK[39];
            assign M_AXIMM_39_AWCACHE = dm_AWCACHE[39];
            assign M_AXIMM_39_AWPROT = dm_AWPROT[39];
            assign M_AXIMM_39_AWREGION = dm_AWREGION[39];
            assign M_AXIMM_39_AWQOS = dm_AWQOS[39];
            assign M_AXIMM_39_AWVALID = dm_AWVALID[39];
            assign dm_AWREADY[39] = M_AXIMM_39_AWREADY;
            assign M_AXIMM_39_WDATA = dm_WDATA[39][M_AXIMM_39_DATA_WIDTH-1:0];
            assign M_AXIMM_39_WSTRB = dm_WSTRB[39][M_AXIMM_39_DATA_WIDTH/8-1:0];
            assign M_AXIMM_39_WLAST = dm_WLAST[39];
            assign M_AXIMM_39_WVALID = dm_WVALID[39];
            assign dm_WREADY[39] = M_AXIMM_39_WREADY;
            assign dm_BRESP[39] = M_AXIMM_39_BRESP;
            assign dm_BVALID[39] = M_AXIMM_39_BVALID;
            assign M_AXIMM_39_BREADY = dm_BREADY[39];
            assign M_AXIMM_39_ARADDR = dm_ARADDR[39][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_39_ARLEN = dm_ARLEN[39];
            assign M_AXIMM_39_ARSIZE = dm_ARSIZE[39];
            assign M_AXIMM_39_ARBURST = dm_ARBURST[39];
            assign M_AXIMM_39_ARLOCK = dm_ARLOCK[39];
            assign M_AXIMM_39_ARCACHE = dm_ARCACHE[39];
            assign M_AXIMM_39_ARPROT = dm_ARPROT[39];
            assign M_AXIMM_39_ARREGION = dm_ARREGION[39];
            assign M_AXIMM_39_ARQOS = dm_ARQOS[39];
            assign M_AXIMM_39_ARVALID = dm_ARVALID[39];
            assign dm_ARREADY[39] = M_AXIMM_39_ARREADY;
            assign dm_RDATA[39][M_AXIMM_39_DATA_WIDTH-1:0] = M_AXIMM_39_RDATA;
            assign dm_RRESP[39] = M_AXIMM_39_RRESP;
            assign dm_RLAST[39] = M_AXIMM_39_RLAST;
            assign dm_RVALID[39] = M_AXIMM_39_RVALID;
            assign M_AXIMM_39_RREADY = dm_RREADY[39];
        end
        if(C_NUM_AXIMMs > 40) begin
            assign ap_AWADDR[40][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_40_AWADDR;
            assign ap_AWLEN[40] = AP_AXIMM_40_AWLEN;
            assign ap_AWSIZE[40] = AP_AXIMM_40_AWSIZE;
            assign ap_AWBURST[40] = AP_AXIMM_40_AWBURST;
            assign ap_AWLOCK[40] = AP_AXIMM_40_AWLOCK;
            assign ap_AWCACHE[40] = AP_AXIMM_40_AWCACHE;
            assign ap_AWPROT[40] = AP_AXIMM_40_AWPROT;
            assign ap_AWREGION[40] = AP_AXIMM_40_AWREGION;
            assign ap_AWQOS[40] = AP_AXIMM_40_AWQOS;
            assign ap_AWVALID[40] = AP_AXIMM_40_AWVALID;
            assign AP_AXIMM_40_AWREADY = ap_AWREADY[40];
            assign ap_WDATA[40][M_AXIMM_40_DATA_WIDTH-1:0] = AP_AXIMM_40_WDATA;
            assign ap_WSTRB[40][M_AXIMM_40_DATA_WIDTH/8-1:0] = AP_AXIMM_40_WSTRB;
            assign ap_WLAST[40] = AP_AXIMM_40_WLAST;
            assign ap_WVALID[40] = AP_AXIMM_40_WVALID;
            assign AP_AXIMM_40_WREADY = ap_WREADY[40];
            assign AP_AXIMM_40_BRESP = ap_BRESP[40];
            assign AP_AXIMM_40_BVALID = ap_BVALID[40];
            assign ap_BREADY[40] = AP_AXIMM_40_BREADY;
            assign ap_ARADDR[40][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_40_ARADDR;
            assign ap_ARLEN[40] = AP_AXIMM_40_ARLEN;
            assign ap_ARSIZE[40] = AP_AXIMM_40_ARSIZE;
            assign ap_ARBURST[40] = AP_AXIMM_40_ARBURST;
            assign ap_ARLOCK[40] = AP_AXIMM_40_ARLOCK;
            assign ap_ARCACHE[40] = AP_AXIMM_40_ARCACHE;
            assign ap_ARPROT[40] = AP_AXIMM_40_ARPROT;
            assign ap_ARREGION[40] = AP_AXIMM_40_ARREGION;
            assign ap_ARQOS[40] = AP_AXIMM_40_ARQOS;
            assign ap_ARVALID[40] = AP_AXIMM_40_ARVALID;
            assign AP_AXIMM_40_ARREADY = ap_ARREADY[40];
            assign AP_AXIMM_40_RDATA = ap_RDATA[40][M_AXIMM_40_DATA_WIDTH-1:0];
            assign AP_AXIMM_40_RRESP = ap_RRESP[40];
            assign AP_AXIMM_40_RLAST = ap_RLAST[40];
            assign AP_AXIMM_40_RVALID = ap_RVALID[40];
            assign ap_RREADY[40] = AP_AXIMM_40_RREADY;
            assign M_AXIMM_40_AWADDR = dm_AWADDR[40][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_40_AWLEN = dm_AWLEN[40];
            assign M_AXIMM_40_AWSIZE = dm_AWSIZE[40];
            assign M_AXIMM_40_AWBURST = dm_AWBURST[40];
            assign M_AXIMM_40_AWLOCK = dm_AWLOCK[40];
            assign M_AXIMM_40_AWCACHE = dm_AWCACHE[40];
            assign M_AXIMM_40_AWPROT = dm_AWPROT[40];
            assign M_AXIMM_40_AWREGION = dm_AWREGION[40];
            assign M_AXIMM_40_AWQOS = dm_AWQOS[40];
            assign M_AXIMM_40_AWVALID = dm_AWVALID[40];
            assign dm_AWREADY[40] = M_AXIMM_40_AWREADY;
            assign M_AXIMM_40_WDATA = dm_WDATA[40][M_AXIMM_40_DATA_WIDTH-1:0];
            assign M_AXIMM_40_WSTRB = dm_WSTRB[40][M_AXIMM_40_DATA_WIDTH/8-1:0];
            assign M_AXIMM_40_WLAST = dm_WLAST[40];
            assign M_AXIMM_40_WVALID = dm_WVALID[40];
            assign dm_WREADY[40] = M_AXIMM_40_WREADY;
            assign dm_BRESP[40] = M_AXIMM_40_BRESP;
            assign dm_BVALID[40] = M_AXIMM_40_BVALID;
            assign M_AXIMM_40_BREADY = dm_BREADY[40];
            assign M_AXIMM_40_ARADDR = dm_ARADDR[40][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_40_ARLEN = dm_ARLEN[40];
            assign M_AXIMM_40_ARSIZE = dm_ARSIZE[40];
            assign M_AXIMM_40_ARBURST = dm_ARBURST[40];
            assign M_AXIMM_40_ARLOCK = dm_ARLOCK[40];
            assign M_AXIMM_40_ARCACHE = dm_ARCACHE[40];
            assign M_AXIMM_40_ARPROT = dm_ARPROT[40];
            assign M_AXIMM_40_ARREGION = dm_ARREGION[40];
            assign M_AXIMM_40_ARQOS = dm_ARQOS[40];
            assign M_AXIMM_40_ARVALID = dm_ARVALID[40];
            assign dm_ARREADY[40] = M_AXIMM_40_ARREADY;
            assign dm_RDATA[40][M_AXIMM_40_DATA_WIDTH-1:0] = M_AXIMM_40_RDATA;
            assign dm_RRESP[40] = M_AXIMM_40_RRESP;
            assign dm_RLAST[40] = M_AXIMM_40_RLAST;
            assign dm_RVALID[40] = M_AXIMM_40_RVALID;
            assign M_AXIMM_40_RREADY = dm_RREADY[40];
        end
        if(C_NUM_AXIMMs > 41) begin
            assign ap_AWADDR[41][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_41_AWADDR;
            assign ap_AWLEN[41] = AP_AXIMM_41_AWLEN;
            assign ap_AWSIZE[41] = AP_AXIMM_41_AWSIZE;
            assign ap_AWBURST[41] = AP_AXIMM_41_AWBURST;
            assign ap_AWLOCK[41] = AP_AXIMM_41_AWLOCK;
            assign ap_AWCACHE[41] = AP_AXIMM_41_AWCACHE;
            assign ap_AWPROT[41] = AP_AXIMM_41_AWPROT;
            assign ap_AWREGION[41] = AP_AXIMM_41_AWREGION;
            assign ap_AWQOS[41] = AP_AXIMM_41_AWQOS;
            assign ap_AWVALID[41] = AP_AXIMM_41_AWVALID;
            assign AP_AXIMM_41_AWREADY = ap_AWREADY[41];
            assign ap_WDATA[41][M_AXIMM_41_DATA_WIDTH-1:0] = AP_AXIMM_41_WDATA;
            assign ap_WSTRB[41][M_AXIMM_41_DATA_WIDTH/8-1:0] = AP_AXIMM_41_WSTRB;
            assign ap_WLAST[41] = AP_AXIMM_41_WLAST;
            assign ap_WVALID[41] = AP_AXIMM_41_WVALID;
            assign AP_AXIMM_41_WREADY = ap_WREADY[41];
            assign AP_AXIMM_41_BRESP = ap_BRESP[41];
            assign AP_AXIMM_41_BVALID = ap_BVALID[41];
            assign ap_BREADY[41] = AP_AXIMM_41_BREADY;
            assign ap_ARADDR[41][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_41_ARADDR;
            assign ap_ARLEN[41] = AP_AXIMM_41_ARLEN;
            assign ap_ARSIZE[41] = AP_AXIMM_41_ARSIZE;
            assign ap_ARBURST[41] = AP_AXIMM_41_ARBURST;
            assign ap_ARLOCK[41] = AP_AXIMM_41_ARLOCK;
            assign ap_ARCACHE[41] = AP_AXIMM_41_ARCACHE;
            assign ap_ARPROT[41] = AP_AXIMM_41_ARPROT;
            assign ap_ARREGION[41] = AP_AXIMM_41_ARREGION;
            assign ap_ARQOS[41] = AP_AXIMM_41_ARQOS;
            assign ap_ARVALID[41] = AP_AXIMM_41_ARVALID;
            assign AP_AXIMM_41_ARREADY = ap_ARREADY[41];
            assign AP_AXIMM_41_RDATA = ap_RDATA[41][M_AXIMM_41_DATA_WIDTH-1:0];
            assign AP_AXIMM_41_RRESP = ap_RRESP[41];
            assign AP_AXIMM_41_RLAST = ap_RLAST[41];
            assign AP_AXIMM_41_RVALID = ap_RVALID[41];
            assign ap_RREADY[41] = AP_AXIMM_41_RREADY;
            assign M_AXIMM_41_AWADDR = dm_AWADDR[41][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_41_AWLEN = dm_AWLEN[41];
            assign M_AXIMM_41_AWSIZE = dm_AWSIZE[41];
            assign M_AXIMM_41_AWBURST = dm_AWBURST[41];
            assign M_AXIMM_41_AWLOCK = dm_AWLOCK[41];
            assign M_AXIMM_41_AWCACHE = dm_AWCACHE[41];
            assign M_AXIMM_41_AWPROT = dm_AWPROT[41];
            assign M_AXIMM_41_AWREGION = dm_AWREGION[41];
            assign M_AXIMM_41_AWQOS = dm_AWQOS[41];
            assign M_AXIMM_41_AWVALID = dm_AWVALID[41];
            assign dm_AWREADY[41] = M_AXIMM_41_AWREADY;
            assign M_AXIMM_41_WDATA = dm_WDATA[41][M_AXIMM_41_DATA_WIDTH-1:0];
            assign M_AXIMM_41_WSTRB = dm_WSTRB[41][M_AXIMM_41_DATA_WIDTH/8-1:0];
            assign M_AXIMM_41_WLAST = dm_WLAST[41];
            assign M_AXIMM_41_WVALID = dm_WVALID[41];
            assign dm_WREADY[41] = M_AXIMM_41_WREADY;
            assign dm_BRESP[41] = M_AXIMM_41_BRESP;
            assign dm_BVALID[41] = M_AXIMM_41_BVALID;
            assign M_AXIMM_41_BREADY = dm_BREADY[41];
            assign M_AXIMM_41_ARADDR = dm_ARADDR[41][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_41_ARLEN = dm_ARLEN[41];
            assign M_AXIMM_41_ARSIZE = dm_ARSIZE[41];
            assign M_AXIMM_41_ARBURST = dm_ARBURST[41];
            assign M_AXIMM_41_ARLOCK = dm_ARLOCK[41];
            assign M_AXIMM_41_ARCACHE = dm_ARCACHE[41];
            assign M_AXIMM_41_ARPROT = dm_ARPROT[41];
            assign M_AXIMM_41_ARREGION = dm_ARREGION[41];
            assign M_AXIMM_41_ARQOS = dm_ARQOS[41];
            assign M_AXIMM_41_ARVALID = dm_ARVALID[41];
            assign dm_ARREADY[41] = M_AXIMM_41_ARREADY;
            assign dm_RDATA[41][M_AXIMM_41_DATA_WIDTH-1:0] = M_AXIMM_41_RDATA;
            assign dm_RRESP[41] = M_AXIMM_41_RRESP;
            assign dm_RLAST[41] = M_AXIMM_41_RLAST;
            assign dm_RVALID[41] = M_AXIMM_41_RVALID;
            assign M_AXIMM_41_RREADY = dm_RREADY[41];
        end
        if(C_NUM_AXIMMs > 42) begin
            assign ap_AWADDR[42][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_42_AWADDR;
            assign ap_AWLEN[42] = AP_AXIMM_42_AWLEN;
            assign ap_AWSIZE[42] = AP_AXIMM_42_AWSIZE;
            assign ap_AWBURST[42] = AP_AXIMM_42_AWBURST;
            assign ap_AWLOCK[42] = AP_AXIMM_42_AWLOCK;
            assign ap_AWCACHE[42] = AP_AXIMM_42_AWCACHE;
            assign ap_AWPROT[42] = AP_AXIMM_42_AWPROT;
            assign ap_AWREGION[42] = AP_AXIMM_42_AWREGION;
            assign ap_AWQOS[42] = AP_AXIMM_42_AWQOS;
            assign ap_AWVALID[42] = AP_AXIMM_42_AWVALID;
            assign AP_AXIMM_42_AWREADY = ap_AWREADY[42];
            assign ap_WDATA[42][M_AXIMM_42_DATA_WIDTH-1:0] = AP_AXIMM_42_WDATA;
            assign ap_WSTRB[42][M_AXIMM_42_DATA_WIDTH/8-1:0] = AP_AXIMM_42_WSTRB;
            assign ap_WLAST[42] = AP_AXIMM_42_WLAST;
            assign ap_WVALID[42] = AP_AXIMM_42_WVALID;
            assign AP_AXIMM_42_WREADY = ap_WREADY[42];
            assign AP_AXIMM_42_BRESP = ap_BRESP[42];
            assign AP_AXIMM_42_BVALID = ap_BVALID[42];
            assign ap_BREADY[42] = AP_AXIMM_42_BREADY;
            assign ap_ARADDR[42][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_42_ARADDR;
            assign ap_ARLEN[42] = AP_AXIMM_42_ARLEN;
            assign ap_ARSIZE[42] = AP_AXIMM_42_ARSIZE;
            assign ap_ARBURST[42] = AP_AXIMM_42_ARBURST;
            assign ap_ARLOCK[42] = AP_AXIMM_42_ARLOCK;
            assign ap_ARCACHE[42] = AP_AXIMM_42_ARCACHE;
            assign ap_ARPROT[42] = AP_AXIMM_42_ARPROT;
            assign ap_ARREGION[42] = AP_AXIMM_42_ARREGION;
            assign ap_ARQOS[42] = AP_AXIMM_42_ARQOS;
            assign ap_ARVALID[42] = AP_AXIMM_42_ARVALID;
            assign AP_AXIMM_42_ARREADY = ap_ARREADY[42];
            assign AP_AXIMM_42_RDATA = ap_RDATA[42][M_AXIMM_42_DATA_WIDTH-1:0];
            assign AP_AXIMM_42_RRESP = ap_RRESP[42];
            assign AP_AXIMM_42_RLAST = ap_RLAST[42];
            assign AP_AXIMM_42_RVALID = ap_RVALID[42];
            assign ap_RREADY[42] = AP_AXIMM_42_RREADY;
            assign M_AXIMM_42_AWADDR = dm_AWADDR[42][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_42_AWLEN = dm_AWLEN[42];
            assign M_AXIMM_42_AWSIZE = dm_AWSIZE[42];
            assign M_AXIMM_42_AWBURST = dm_AWBURST[42];
            assign M_AXIMM_42_AWLOCK = dm_AWLOCK[42];
            assign M_AXIMM_42_AWCACHE = dm_AWCACHE[42];
            assign M_AXIMM_42_AWPROT = dm_AWPROT[42];
            assign M_AXIMM_42_AWREGION = dm_AWREGION[42];
            assign M_AXIMM_42_AWQOS = dm_AWQOS[42];
            assign M_AXIMM_42_AWVALID = dm_AWVALID[42];
            assign dm_AWREADY[42] = M_AXIMM_42_AWREADY;
            assign M_AXIMM_42_WDATA = dm_WDATA[42][M_AXIMM_42_DATA_WIDTH-1:0];
            assign M_AXIMM_42_WSTRB = dm_WSTRB[42][M_AXIMM_42_DATA_WIDTH/8-1:0];
            assign M_AXIMM_42_WLAST = dm_WLAST[42];
            assign M_AXIMM_42_WVALID = dm_WVALID[42];
            assign dm_WREADY[42] = M_AXIMM_42_WREADY;
            assign dm_BRESP[42] = M_AXIMM_42_BRESP;
            assign dm_BVALID[42] = M_AXIMM_42_BVALID;
            assign M_AXIMM_42_BREADY = dm_BREADY[42];
            assign M_AXIMM_42_ARADDR = dm_ARADDR[42][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_42_ARLEN = dm_ARLEN[42];
            assign M_AXIMM_42_ARSIZE = dm_ARSIZE[42];
            assign M_AXIMM_42_ARBURST = dm_ARBURST[42];
            assign M_AXIMM_42_ARLOCK = dm_ARLOCK[42];
            assign M_AXIMM_42_ARCACHE = dm_ARCACHE[42];
            assign M_AXIMM_42_ARPROT = dm_ARPROT[42];
            assign M_AXIMM_42_ARREGION = dm_ARREGION[42];
            assign M_AXIMM_42_ARQOS = dm_ARQOS[42];
            assign M_AXIMM_42_ARVALID = dm_ARVALID[42];
            assign dm_ARREADY[42] = M_AXIMM_42_ARREADY;
            assign dm_RDATA[42][M_AXIMM_42_DATA_WIDTH-1:0] = M_AXIMM_42_RDATA;
            assign dm_RRESP[42] = M_AXIMM_42_RRESP;
            assign dm_RLAST[42] = M_AXIMM_42_RLAST;
            assign dm_RVALID[42] = M_AXIMM_42_RVALID;
            assign M_AXIMM_42_RREADY = dm_RREADY[42];
        end
        if(C_NUM_AXIMMs > 43) begin
            assign ap_AWADDR[43][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_43_AWADDR;
            assign ap_AWLEN[43] = AP_AXIMM_43_AWLEN;
            assign ap_AWSIZE[43] = AP_AXIMM_43_AWSIZE;
            assign ap_AWBURST[43] = AP_AXIMM_43_AWBURST;
            assign ap_AWLOCK[43] = AP_AXIMM_43_AWLOCK;
            assign ap_AWCACHE[43] = AP_AXIMM_43_AWCACHE;
            assign ap_AWPROT[43] = AP_AXIMM_43_AWPROT;
            assign ap_AWREGION[43] = AP_AXIMM_43_AWREGION;
            assign ap_AWQOS[43] = AP_AXIMM_43_AWQOS;
            assign ap_AWVALID[43] = AP_AXIMM_43_AWVALID;
            assign AP_AXIMM_43_AWREADY = ap_AWREADY[43];
            assign ap_WDATA[43][M_AXIMM_43_DATA_WIDTH-1:0] = AP_AXIMM_43_WDATA;
            assign ap_WSTRB[43][M_AXIMM_43_DATA_WIDTH/8-1:0] = AP_AXIMM_43_WSTRB;
            assign ap_WLAST[43] = AP_AXIMM_43_WLAST;
            assign ap_WVALID[43] = AP_AXIMM_43_WVALID;
            assign AP_AXIMM_43_WREADY = ap_WREADY[43];
            assign AP_AXIMM_43_BRESP = ap_BRESP[43];
            assign AP_AXIMM_43_BVALID = ap_BVALID[43];
            assign ap_BREADY[43] = AP_AXIMM_43_BREADY;
            assign ap_ARADDR[43][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_43_ARADDR;
            assign ap_ARLEN[43] = AP_AXIMM_43_ARLEN;
            assign ap_ARSIZE[43] = AP_AXIMM_43_ARSIZE;
            assign ap_ARBURST[43] = AP_AXIMM_43_ARBURST;
            assign ap_ARLOCK[43] = AP_AXIMM_43_ARLOCK;
            assign ap_ARCACHE[43] = AP_AXIMM_43_ARCACHE;
            assign ap_ARPROT[43] = AP_AXIMM_43_ARPROT;
            assign ap_ARREGION[43] = AP_AXIMM_43_ARREGION;
            assign ap_ARQOS[43] = AP_AXIMM_43_ARQOS;
            assign ap_ARVALID[43] = AP_AXIMM_43_ARVALID;
            assign AP_AXIMM_43_ARREADY = ap_ARREADY[43];
            assign AP_AXIMM_43_RDATA = ap_RDATA[43][M_AXIMM_43_DATA_WIDTH-1:0];
            assign AP_AXIMM_43_RRESP = ap_RRESP[43];
            assign AP_AXIMM_43_RLAST = ap_RLAST[43];
            assign AP_AXIMM_43_RVALID = ap_RVALID[43];
            assign ap_RREADY[43] = AP_AXIMM_43_RREADY;
            assign M_AXIMM_43_AWADDR = dm_AWADDR[43][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_43_AWLEN = dm_AWLEN[43];
            assign M_AXIMM_43_AWSIZE = dm_AWSIZE[43];
            assign M_AXIMM_43_AWBURST = dm_AWBURST[43];
            assign M_AXIMM_43_AWLOCK = dm_AWLOCK[43];
            assign M_AXIMM_43_AWCACHE = dm_AWCACHE[43];
            assign M_AXIMM_43_AWPROT = dm_AWPROT[43];
            assign M_AXIMM_43_AWREGION = dm_AWREGION[43];
            assign M_AXIMM_43_AWQOS = dm_AWQOS[43];
            assign M_AXIMM_43_AWVALID = dm_AWVALID[43];
            assign dm_AWREADY[43] = M_AXIMM_43_AWREADY;
            assign M_AXIMM_43_WDATA = dm_WDATA[43][M_AXIMM_43_DATA_WIDTH-1:0];
            assign M_AXIMM_43_WSTRB = dm_WSTRB[43][M_AXIMM_43_DATA_WIDTH/8-1:0];
            assign M_AXIMM_43_WLAST = dm_WLAST[43];
            assign M_AXIMM_43_WVALID = dm_WVALID[43];
            assign dm_WREADY[43] = M_AXIMM_43_WREADY;
            assign dm_BRESP[43] = M_AXIMM_43_BRESP;
            assign dm_BVALID[43] = M_AXIMM_43_BVALID;
            assign M_AXIMM_43_BREADY = dm_BREADY[43];
            assign M_AXIMM_43_ARADDR = dm_ARADDR[43][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_43_ARLEN = dm_ARLEN[43];
            assign M_AXIMM_43_ARSIZE = dm_ARSIZE[43];
            assign M_AXIMM_43_ARBURST = dm_ARBURST[43];
            assign M_AXIMM_43_ARLOCK = dm_ARLOCK[43];
            assign M_AXIMM_43_ARCACHE = dm_ARCACHE[43];
            assign M_AXIMM_43_ARPROT = dm_ARPROT[43];
            assign M_AXIMM_43_ARREGION = dm_ARREGION[43];
            assign M_AXIMM_43_ARQOS = dm_ARQOS[43];
            assign M_AXIMM_43_ARVALID = dm_ARVALID[43];
            assign dm_ARREADY[43] = M_AXIMM_43_ARREADY;
            assign dm_RDATA[43][M_AXIMM_43_DATA_WIDTH-1:0] = M_AXIMM_43_RDATA;
            assign dm_RRESP[43] = M_AXIMM_43_RRESP;
            assign dm_RLAST[43] = M_AXIMM_43_RLAST;
            assign dm_RVALID[43] = M_AXIMM_43_RVALID;
            assign M_AXIMM_43_RREADY = dm_RREADY[43];
        end
        if(C_NUM_AXIMMs > 44) begin
            assign ap_AWADDR[44][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_44_AWADDR;
            assign ap_AWLEN[44] = AP_AXIMM_44_AWLEN;
            assign ap_AWSIZE[44] = AP_AXIMM_44_AWSIZE;
            assign ap_AWBURST[44] = AP_AXIMM_44_AWBURST;
            assign ap_AWLOCK[44] = AP_AXIMM_44_AWLOCK;
            assign ap_AWCACHE[44] = AP_AXIMM_44_AWCACHE;
            assign ap_AWPROT[44] = AP_AXIMM_44_AWPROT;
            assign ap_AWREGION[44] = AP_AXIMM_44_AWREGION;
            assign ap_AWQOS[44] = AP_AXIMM_44_AWQOS;
            assign ap_AWVALID[44] = AP_AXIMM_44_AWVALID;
            assign AP_AXIMM_44_AWREADY = ap_AWREADY[44];
            assign ap_WDATA[44][M_AXIMM_44_DATA_WIDTH-1:0] = AP_AXIMM_44_WDATA;
            assign ap_WSTRB[44][M_AXIMM_44_DATA_WIDTH/8-1:0] = AP_AXIMM_44_WSTRB;
            assign ap_WLAST[44] = AP_AXIMM_44_WLAST;
            assign ap_WVALID[44] = AP_AXIMM_44_WVALID;
            assign AP_AXIMM_44_WREADY = ap_WREADY[44];
            assign AP_AXIMM_44_BRESP = ap_BRESP[44];
            assign AP_AXIMM_44_BVALID = ap_BVALID[44];
            assign ap_BREADY[44] = AP_AXIMM_44_BREADY;
            assign ap_ARADDR[44][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_44_ARADDR;
            assign ap_ARLEN[44] = AP_AXIMM_44_ARLEN;
            assign ap_ARSIZE[44] = AP_AXIMM_44_ARSIZE;
            assign ap_ARBURST[44] = AP_AXIMM_44_ARBURST;
            assign ap_ARLOCK[44] = AP_AXIMM_44_ARLOCK;
            assign ap_ARCACHE[44] = AP_AXIMM_44_ARCACHE;
            assign ap_ARPROT[44] = AP_AXIMM_44_ARPROT;
            assign ap_ARREGION[44] = AP_AXIMM_44_ARREGION;
            assign ap_ARQOS[44] = AP_AXIMM_44_ARQOS;
            assign ap_ARVALID[44] = AP_AXIMM_44_ARVALID;
            assign AP_AXIMM_44_ARREADY = ap_ARREADY[44];
            assign AP_AXIMM_44_RDATA = ap_RDATA[44][M_AXIMM_44_DATA_WIDTH-1:0];
            assign AP_AXIMM_44_RRESP = ap_RRESP[44];
            assign AP_AXIMM_44_RLAST = ap_RLAST[44];
            assign AP_AXIMM_44_RVALID = ap_RVALID[44];
            assign ap_RREADY[44] = AP_AXIMM_44_RREADY;
            assign M_AXIMM_44_AWADDR = dm_AWADDR[44][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_44_AWLEN = dm_AWLEN[44];
            assign M_AXIMM_44_AWSIZE = dm_AWSIZE[44];
            assign M_AXIMM_44_AWBURST = dm_AWBURST[44];
            assign M_AXIMM_44_AWLOCK = dm_AWLOCK[44];
            assign M_AXIMM_44_AWCACHE = dm_AWCACHE[44];
            assign M_AXIMM_44_AWPROT = dm_AWPROT[44];
            assign M_AXIMM_44_AWREGION = dm_AWREGION[44];
            assign M_AXIMM_44_AWQOS = dm_AWQOS[44];
            assign M_AXIMM_44_AWVALID = dm_AWVALID[44];
            assign dm_AWREADY[44] = M_AXIMM_44_AWREADY;
            assign M_AXIMM_44_WDATA = dm_WDATA[44][M_AXIMM_44_DATA_WIDTH-1:0];
            assign M_AXIMM_44_WSTRB = dm_WSTRB[44][M_AXIMM_44_DATA_WIDTH/8-1:0];
            assign M_AXIMM_44_WLAST = dm_WLAST[44];
            assign M_AXIMM_44_WVALID = dm_WVALID[44];
            assign dm_WREADY[44] = M_AXIMM_44_WREADY;
            assign dm_BRESP[44] = M_AXIMM_44_BRESP;
            assign dm_BVALID[44] = M_AXIMM_44_BVALID;
            assign M_AXIMM_44_BREADY = dm_BREADY[44];
            assign M_AXIMM_44_ARADDR = dm_ARADDR[44][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_44_ARLEN = dm_ARLEN[44];
            assign M_AXIMM_44_ARSIZE = dm_ARSIZE[44];
            assign M_AXIMM_44_ARBURST = dm_ARBURST[44];
            assign M_AXIMM_44_ARLOCK = dm_ARLOCK[44];
            assign M_AXIMM_44_ARCACHE = dm_ARCACHE[44];
            assign M_AXIMM_44_ARPROT = dm_ARPROT[44];
            assign M_AXIMM_44_ARREGION = dm_ARREGION[44];
            assign M_AXIMM_44_ARQOS = dm_ARQOS[44];
            assign M_AXIMM_44_ARVALID = dm_ARVALID[44];
            assign dm_ARREADY[44] = M_AXIMM_44_ARREADY;
            assign dm_RDATA[44][M_AXIMM_44_DATA_WIDTH-1:0] = M_AXIMM_44_RDATA;
            assign dm_RRESP[44] = M_AXIMM_44_RRESP;
            assign dm_RLAST[44] = M_AXIMM_44_RLAST;
            assign dm_RVALID[44] = M_AXIMM_44_RVALID;
            assign M_AXIMM_44_RREADY = dm_RREADY[44];
        end
        if(C_NUM_AXIMMs > 45) begin
            assign ap_AWADDR[45][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_45_AWADDR;
            assign ap_AWLEN[45] = AP_AXIMM_45_AWLEN;
            assign ap_AWSIZE[45] = AP_AXIMM_45_AWSIZE;
            assign ap_AWBURST[45] = AP_AXIMM_45_AWBURST;
            assign ap_AWLOCK[45] = AP_AXIMM_45_AWLOCK;
            assign ap_AWCACHE[45] = AP_AXIMM_45_AWCACHE;
            assign ap_AWPROT[45] = AP_AXIMM_45_AWPROT;
            assign ap_AWREGION[45] = AP_AXIMM_45_AWREGION;
            assign ap_AWQOS[45] = AP_AXIMM_45_AWQOS;
            assign ap_AWVALID[45] = AP_AXIMM_45_AWVALID;
            assign AP_AXIMM_45_AWREADY = ap_AWREADY[45];
            assign ap_WDATA[45][M_AXIMM_45_DATA_WIDTH-1:0] = AP_AXIMM_45_WDATA;
            assign ap_WSTRB[45][M_AXIMM_45_DATA_WIDTH/8-1:0] = AP_AXIMM_45_WSTRB;
            assign ap_WLAST[45] = AP_AXIMM_45_WLAST;
            assign ap_WVALID[45] = AP_AXIMM_45_WVALID;
            assign AP_AXIMM_45_WREADY = ap_WREADY[45];
            assign AP_AXIMM_45_BRESP = ap_BRESP[45];
            assign AP_AXIMM_45_BVALID = ap_BVALID[45];
            assign ap_BREADY[45] = AP_AXIMM_45_BREADY;
            assign ap_ARADDR[45][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_45_ARADDR;
            assign ap_ARLEN[45] = AP_AXIMM_45_ARLEN;
            assign ap_ARSIZE[45] = AP_AXIMM_45_ARSIZE;
            assign ap_ARBURST[45] = AP_AXIMM_45_ARBURST;
            assign ap_ARLOCK[45] = AP_AXIMM_45_ARLOCK;
            assign ap_ARCACHE[45] = AP_AXIMM_45_ARCACHE;
            assign ap_ARPROT[45] = AP_AXIMM_45_ARPROT;
            assign ap_ARREGION[45] = AP_AXIMM_45_ARREGION;
            assign ap_ARQOS[45] = AP_AXIMM_45_ARQOS;
            assign ap_ARVALID[45] = AP_AXIMM_45_ARVALID;
            assign AP_AXIMM_45_ARREADY = ap_ARREADY[45];
            assign AP_AXIMM_45_RDATA = ap_RDATA[45][M_AXIMM_45_DATA_WIDTH-1:0];
            assign AP_AXIMM_45_RRESP = ap_RRESP[45];
            assign AP_AXIMM_45_RLAST = ap_RLAST[45];
            assign AP_AXIMM_45_RVALID = ap_RVALID[45];
            assign ap_RREADY[45] = AP_AXIMM_45_RREADY;
            assign M_AXIMM_45_AWADDR = dm_AWADDR[45][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_45_AWLEN = dm_AWLEN[45];
            assign M_AXIMM_45_AWSIZE = dm_AWSIZE[45];
            assign M_AXIMM_45_AWBURST = dm_AWBURST[45];
            assign M_AXIMM_45_AWLOCK = dm_AWLOCK[45];
            assign M_AXIMM_45_AWCACHE = dm_AWCACHE[45];
            assign M_AXIMM_45_AWPROT = dm_AWPROT[45];
            assign M_AXIMM_45_AWREGION = dm_AWREGION[45];
            assign M_AXIMM_45_AWQOS = dm_AWQOS[45];
            assign M_AXIMM_45_AWVALID = dm_AWVALID[45];
            assign dm_AWREADY[45] = M_AXIMM_45_AWREADY;
            assign M_AXIMM_45_WDATA = dm_WDATA[45][M_AXIMM_45_DATA_WIDTH-1:0];
            assign M_AXIMM_45_WSTRB = dm_WSTRB[45][M_AXIMM_45_DATA_WIDTH/8-1:0];
            assign M_AXIMM_45_WLAST = dm_WLAST[45];
            assign M_AXIMM_45_WVALID = dm_WVALID[45];
            assign dm_WREADY[45] = M_AXIMM_45_WREADY;
            assign dm_BRESP[45] = M_AXIMM_45_BRESP;
            assign dm_BVALID[45] = M_AXIMM_45_BVALID;
            assign M_AXIMM_45_BREADY = dm_BREADY[45];
            assign M_AXIMM_45_ARADDR = dm_ARADDR[45][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_45_ARLEN = dm_ARLEN[45];
            assign M_AXIMM_45_ARSIZE = dm_ARSIZE[45];
            assign M_AXIMM_45_ARBURST = dm_ARBURST[45];
            assign M_AXIMM_45_ARLOCK = dm_ARLOCK[45];
            assign M_AXIMM_45_ARCACHE = dm_ARCACHE[45];
            assign M_AXIMM_45_ARPROT = dm_ARPROT[45];
            assign M_AXIMM_45_ARREGION = dm_ARREGION[45];
            assign M_AXIMM_45_ARQOS = dm_ARQOS[45];
            assign M_AXIMM_45_ARVALID = dm_ARVALID[45];
            assign dm_ARREADY[45] = M_AXIMM_45_ARREADY;
            assign dm_RDATA[45][M_AXIMM_45_DATA_WIDTH-1:0] = M_AXIMM_45_RDATA;
            assign dm_RRESP[45] = M_AXIMM_45_RRESP;
            assign dm_RLAST[45] = M_AXIMM_45_RLAST;
            assign dm_RVALID[45] = M_AXIMM_45_RVALID;
            assign M_AXIMM_45_RREADY = dm_RREADY[45];
        end
        if(C_NUM_AXIMMs > 46) begin
            assign ap_AWADDR[46][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_46_AWADDR;
            assign ap_AWLEN[46] = AP_AXIMM_46_AWLEN;
            assign ap_AWSIZE[46] = AP_AXIMM_46_AWSIZE;
            assign ap_AWBURST[46] = AP_AXIMM_46_AWBURST;
            assign ap_AWLOCK[46] = AP_AXIMM_46_AWLOCK;
            assign ap_AWCACHE[46] = AP_AXIMM_46_AWCACHE;
            assign ap_AWPROT[46] = AP_AXIMM_46_AWPROT;
            assign ap_AWREGION[46] = AP_AXIMM_46_AWREGION;
            assign ap_AWQOS[46] = AP_AXIMM_46_AWQOS;
            assign ap_AWVALID[46] = AP_AXIMM_46_AWVALID;
            assign AP_AXIMM_46_AWREADY = ap_AWREADY[46];
            assign ap_WDATA[46][M_AXIMM_46_DATA_WIDTH-1:0] = AP_AXIMM_46_WDATA;
            assign ap_WSTRB[46][M_AXIMM_46_DATA_WIDTH/8-1:0] = AP_AXIMM_46_WSTRB;
            assign ap_WLAST[46] = AP_AXIMM_46_WLAST;
            assign ap_WVALID[46] = AP_AXIMM_46_WVALID;
            assign AP_AXIMM_46_WREADY = ap_WREADY[46];
            assign AP_AXIMM_46_BRESP = ap_BRESP[46];
            assign AP_AXIMM_46_BVALID = ap_BVALID[46];
            assign ap_BREADY[46] = AP_AXIMM_46_BREADY;
            assign ap_ARADDR[46][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_46_ARADDR;
            assign ap_ARLEN[46] = AP_AXIMM_46_ARLEN;
            assign ap_ARSIZE[46] = AP_AXIMM_46_ARSIZE;
            assign ap_ARBURST[46] = AP_AXIMM_46_ARBURST;
            assign ap_ARLOCK[46] = AP_AXIMM_46_ARLOCK;
            assign ap_ARCACHE[46] = AP_AXIMM_46_ARCACHE;
            assign ap_ARPROT[46] = AP_AXIMM_46_ARPROT;
            assign ap_ARREGION[46] = AP_AXIMM_46_ARREGION;
            assign ap_ARQOS[46] = AP_AXIMM_46_ARQOS;
            assign ap_ARVALID[46] = AP_AXIMM_46_ARVALID;
            assign AP_AXIMM_46_ARREADY = ap_ARREADY[46];
            assign AP_AXIMM_46_RDATA = ap_RDATA[46][M_AXIMM_46_DATA_WIDTH-1:0];
            assign AP_AXIMM_46_RRESP = ap_RRESP[46];
            assign AP_AXIMM_46_RLAST = ap_RLAST[46];
            assign AP_AXIMM_46_RVALID = ap_RVALID[46];
            assign ap_RREADY[46] = AP_AXIMM_46_RREADY;
            assign M_AXIMM_46_AWADDR = dm_AWADDR[46][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_46_AWLEN = dm_AWLEN[46];
            assign M_AXIMM_46_AWSIZE = dm_AWSIZE[46];
            assign M_AXIMM_46_AWBURST = dm_AWBURST[46];
            assign M_AXIMM_46_AWLOCK = dm_AWLOCK[46];
            assign M_AXIMM_46_AWCACHE = dm_AWCACHE[46];
            assign M_AXIMM_46_AWPROT = dm_AWPROT[46];
            assign M_AXIMM_46_AWREGION = dm_AWREGION[46];
            assign M_AXIMM_46_AWQOS = dm_AWQOS[46];
            assign M_AXIMM_46_AWVALID = dm_AWVALID[46];
            assign dm_AWREADY[46] = M_AXIMM_46_AWREADY;
            assign M_AXIMM_46_WDATA = dm_WDATA[46][M_AXIMM_46_DATA_WIDTH-1:0];
            assign M_AXIMM_46_WSTRB = dm_WSTRB[46][M_AXIMM_46_DATA_WIDTH/8-1:0];
            assign M_AXIMM_46_WLAST = dm_WLAST[46];
            assign M_AXIMM_46_WVALID = dm_WVALID[46];
            assign dm_WREADY[46] = M_AXIMM_46_WREADY;
            assign dm_BRESP[46] = M_AXIMM_46_BRESP;
            assign dm_BVALID[46] = M_AXIMM_46_BVALID;
            assign M_AXIMM_46_BREADY = dm_BREADY[46];
            assign M_AXIMM_46_ARADDR = dm_ARADDR[46][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_46_ARLEN = dm_ARLEN[46];
            assign M_AXIMM_46_ARSIZE = dm_ARSIZE[46];
            assign M_AXIMM_46_ARBURST = dm_ARBURST[46];
            assign M_AXIMM_46_ARLOCK = dm_ARLOCK[46];
            assign M_AXIMM_46_ARCACHE = dm_ARCACHE[46];
            assign M_AXIMM_46_ARPROT = dm_ARPROT[46];
            assign M_AXIMM_46_ARREGION = dm_ARREGION[46];
            assign M_AXIMM_46_ARQOS = dm_ARQOS[46];
            assign M_AXIMM_46_ARVALID = dm_ARVALID[46];
            assign dm_ARREADY[46] = M_AXIMM_46_ARREADY;
            assign dm_RDATA[46][M_AXIMM_46_DATA_WIDTH-1:0] = M_AXIMM_46_RDATA;
            assign dm_RRESP[46] = M_AXIMM_46_RRESP;
            assign dm_RLAST[46] = M_AXIMM_46_RLAST;
            assign dm_RVALID[46] = M_AXIMM_46_RVALID;
            assign M_AXIMM_46_RREADY = dm_RREADY[46];
        end
        if(C_NUM_AXIMMs > 47) begin
            assign ap_AWADDR[47][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_47_AWADDR;
            assign ap_AWLEN[47] = AP_AXIMM_47_AWLEN;
            assign ap_AWSIZE[47] = AP_AXIMM_47_AWSIZE;
            assign ap_AWBURST[47] = AP_AXIMM_47_AWBURST;
            assign ap_AWLOCK[47] = AP_AXIMM_47_AWLOCK;
            assign ap_AWCACHE[47] = AP_AXIMM_47_AWCACHE;
            assign ap_AWPROT[47] = AP_AXIMM_47_AWPROT;
            assign ap_AWREGION[47] = AP_AXIMM_47_AWREGION;
            assign ap_AWQOS[47] = AP_AXIMM_47_AWQOS;
            assign ap_AWVALID[47] = AP_AXIMM_47_AWVALID;
            assign AP_AXIMM_47_AWREADY = ap_AWREADY[47];
            assign ap_WDATA[47][M_AXIMM_47_DATA_WIDTH-1:0] = AP_AXIMM_47_WDATA;
            assign ap_WSTRB[47][M_AXIMM_47_DATA_WIDTH/8-1:0] = AP_AXIMM_47_WSTRB;
            assign ap_WLAST[47] = AP_AXIMM_47_WLAST;
            assign ap_WVALID[47] = AP_AXIMM_47_WVALID;
            assign AP_AXIMM_47_WREADY = ap_WREADY[47];
            assign AP_AXIMM_47_BRESP = ap_BRESP[47];
            assign AP_AXIMM_47_BVALID = ap_BVALID[47];
            assign ap_BREADY[47] = AP_AXIMM_47_BREADY;
            assign ap_ARADDR[47][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_47_ARADDR;
            assign ap_ARLEN[47] = AP_AXIMM_47_ARLEN;
            assign ap_ARSIZE[47] = AP_AXIMM_47_ARSIZE;
            assign ap_ARBURST[47] = AP_AXIMM_47_ARBURST;
            assign ap_ARLOCK[47] = AP_AXIMM_47_ARLOCK;
            assign ap_ARCACHE[47] = AP_AXIMM_47_ARCACHE;
            assign ap_ARPROT[47] = AP_AXIMM_47_ARPROT;
            assign ap_ARREGION[47] = AP_AXIMM_47_ARREGION;
            assign ap_ARQOS[47] = AP_AXIMM_47_ARQOS;
            assign ap_ARVALID[47] = AP_AXIMM_47_ARVALID;
            assign AP_AXIMM_47_ARREADY = ap_ARREADY[47];
            assign AP_AXIMM_47_RDATA = ap_RDATA[47][M_AXIMM_47_DATA_WIDTH-1:0];
            assign AP_AXIMM_47_RRESP = ap_RRESP[47];
            assign AP_AXIMM_47_RLAST = ap_RLAST[47];
            assign AP_AXIMM_47_RVALID = ap_RVALID[47];
            assign ap_RREADY[47] = AP_AXIMM_47_RREADY;
            assign M_AXIMM_47_AWADDR = dm_AWADDR[47][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_47_AWLEN = dm_AWLEN[47];
            assign M_AXIMM_47_AWSIZE = dm_AWSIZE[47];
            assign M_AXIMM_47_AWBURST = dm_AWBURST[47];
            assign M_AXIMM_47_AWLOCK = dm_AWLOCK[47];
            assign M_AXIMM_47_AWCACHE = dm_AWCACHE[47];
            assign M_AXIMM_47_AWPROT = dm_AWPROT[47];
            assign M_AXIMM_47_AWREGION = dm_AWREGION[47];
            assign M_AXIMM_47_AWQOS = dm_AWQOS[47];
            assign M_AXIMM_47_AWVALID = dm_AWVALID[47];
            assign dm_AWREADY[47] = M_AXIMM_47_AWREADY;
            assign M_AXIMM_47_WDATA = dm_WDATA[47][M_AXIMM_47_DATA_WIDTH-1:0];
            assign M_AXIMM_47_WSTRB = dm_WSTRB[47][M_AXIMM_47_DATA_WIDTH/8-1:0];
            assign M_AXIMM_47_WLAST = dm_WLAST[47];
            assign M_AXIMM_47_WVALID = dm_WVALID[47];
            assign dm_WREADY[47] = M_AXIMM_47_WREADY;
            assign dm_BRESP[47] = M_AXIMM_47_BRESP;
            assign dm_BVALID[47] = M_AXIMM_47_BVALID;
            assign M_AXIMM_47_BREADY = dm_BREADY[47];
            assign M_AXIMM_47_ARADDR = dm_ARADDR[47][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_47_ARLEN = dm_ARLEN[47];
            assign M_AXIMM_47_ARSIZE = dm_ARSIZE[47];
            assign M_AXIMM_47_ARBURST = dm_ARBURST[47];
            assign M_AXIMM_47_ARLOCK = dm_ARLOCK[47];
            assign M_AXIMM_47_ARCACHE = dm_ARCACHE[47];
            assign M_AXIMM_47_ARPROT = dm_ARPROT[47];
            assign M_AXIMM_47_ARREGION = dm_ARREGION[47];
            assign M_AXIMM_47_ARQOS = dm_ARQOS[47];
            assign M_AXIMM_47_ARVALID = dm_ARVALID[47];
            assign dm_ARREADY[47] = M_AXIMM_47_ARREADY;
            assign dm_RDATA[47][M_AXIMM_47_DATA_WIDTH-1:0] = M_AXIMM_47_RDATA;
            assign dm_RRESP[47] = M_AXIMM_47_RRESP;
            assign dm_RLAST[47] = M_AXIMM_47_RLAST;
            assign dm_RVALID[47] = M_AXIMM_47_RVALID;
            assign M_AXIMM_47_RREADY = dm_RREADY[47];
        end
        if(C_NUM_AXIMMs > 48) begin
            assign ap_AWADDR[48][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_48_AWADDR;
            assign ap_AWLEN[48] = AP_AXIMM_48_AWLEN;
            assign ap_AWSIZE[48] = AP_AXIMM_48_AWSIZE;
            assign ap_AWBURST[48] = AP_AXIMM_48_AWBURST;
            assign ap_AWLOCK[48] = AP_AXIMM_48_AWLOCK;
            assign ap_AWCACHE[48] = AP_AXIMM_48_AWCACHE;
            assign ap_AWPROT[48] = AP_AXIMM_48_AWPROT;
            assign ap_AWREGION[48] = AP_AXIMM_48_AWREGION;
            assign ap_AWQOS[48] = AP_AXIMM_48_AWQOS;
            assign ap_AWVALID[48] = AP_AXIMM_48_AWVALID;
            assign AP_AXIMM_48_AWREADY = ap_AWREADY[48];
            assign ap_WDATA[48][M_AXIMM_48_DATA_WIDTH-1:0] = AP_AXIMM_48_WDATA;
            assign ap_WSTRB[48][M_AXIMM_48_DATA_WIDTH/8-1:0] = AP_AXIMM_48_WSTRB;
            assign ap_WLAST[48] = AP_AXIMM_48_WLAST;
            assign ap_WVALID[48] = AP_AXIMM_48_WVALID;
            assign AP_AXIMM_48_WREADY = ap_WREADY[48];
            assign AP_AXIMM_48_BRESP = ap_BRESP[48];
            assign AP_AXIMM_48_BVALID = ap_BVALID[48];
            assign ap_BREADY[48] = AP_AXIMM_48_BREADY;
            assign ap_ARADDR[48][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_48_ARADDR;
            assign ap_ARLEN[48] = AP_AXIMM_48_ARLEN;
            assign ap_ARSIZE[48] = AP_AXIMM_48_ARSIZE;
            assign ap_ARBURST[48] = AP_AXIMM_48_ARBURST;
            assign ap_ARLOCK[48] = AP_AXIMM_48_ARLOCK;
            assign ap_ARCACHE[48] = AP_AXIMM_48_ARCACHE;
            assign ap_ARPROT[48] = AP_AXIMM_48_ARPROT;
            assign ap_ARREGION[48] = AP_AXIMM_48_ARREGION;
            assign ap_ARQOS[48] = AP_AXIMM_48_ARQOS;
            assign ap_ARVALID[48] = AP_AXIMM_48_ARVALID;
            assign AP_AXIMM_48_ARREADY = ap_ARREADY[48];
            assign AP_AXIMM_48_RDATA = ap_RDATA[48][M_AXIMM_48_DATA_WIDTH-1:0];
            assign AP_AXIMM_48_RRESP = ap_RRESP[48];
            assign AP_AXIMM_48_RLAST = ap_RLAST[48];
            assign AP_AXIMM_48_RVALID = ap_RVALID[48];
            assign ap_RREADY[48] = AP_AXIMM_48_RREADY;
            assign M_AXIMM_48_AWADDR = dm_AWADDR[48][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_48_AWLEN = dm_AWLEN[48];
            assign M_AXIMM_48_AWSIZE = dm_AWSIZE[48];
            assign M_AXIMM_48_AWBURST = dm_AWBURST[48];
            assign M_AXIMM_48_AWLOCK = dm_AWLOCK[48];
            assign M_AXIMM_48_AWCACHE = dm_AWCACHE[48];
            assign M_AXIMM_48_AWPROT = dm_AWPROT[48];
            assign M_AXIMM_48_AWREGION = dm_AWREGION[48];
            assign M_AXIMM_48_AWQOS = dm_AWQOS[48];
            assign M_AXIMM_48_AWVALID = dm_AWVALID[48];
            assign dm_AWREADY[48] = M_AXIMM_48_AWREADY;
            assign M_AXIMM_48_WDATA = dm_WDATA[48][M_AXIMM_48_DATA_WIDTH-1:0];
            assign M_AXIMM_48_WSTRB = dm_WSTRB[48][M_AXIMM_48_DATA_WIDTH/8-1:0];
            assign M_AXIMM_48_WLAST = dm_WLAST[48];
            assign M_AXIMM_48_WVALID = dm_WVALID[48];
            assign dm_WREADY[48] = M_AXIMM_48_WREADY;
            assign dm_BRESP[48] = M_AXIMM_48_BRESP;
            assign dm_BVALID[48] = M_AXIMM_48_BVALID;
            assign M_AXIMM_48_BREADY = dm_BREADY[48];
            assign M_AXIMM_48_ARADDR = dm_ARADDR[48][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_48_ARLEN = dm_ARLEN[48];
            assign M_AXIMM_48_ARSIZE = dm_ARSIZE[48];
            assign M_AXIMM_48_ARBURST = dm_ARBURST[48];
            assign M_AXIMM_48_ARLOCK = dm_ARLOCK[48];
            assign M_AXIMM_48_ARCACHE = dm_ARCACHE[48];
            assign M_AXIMM_48_ARPROT = dm_ARPROT[48];
            assign M_AXIMM_48_ARREGION = dm_ARREGION[48];
            assign M_AXIMM_48_ARQOS = dm_ARQOS[48];
            assign M_AXIMM_48_ARVALID = dm_ARVALID[48];
            assign dm_ARREADY[48] = M_AXIMM_48_ARREADY;
            assign dm_RDATA[48][M_AXIMM_48_DATA_WIDTH-1:0] = M_AXIMM_48_RDATA;
            assign dm_RRESP[48] = M_AXIMM_48_RRESP;
            assign dm_RLAST[48] = M_AXIMM_48_RLAST;
            assign dm_RVALID[48] = M_AXIMM_48_RVALID;
            assign M_AXIMM_48_RREADY = dm_RREADY[48];
        end
        if(C_NUM_AXIMMs > 49) begin
            assign ap_AWADDR[49][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_49_AWADDR;
            assign ap_AWLEN[49] = AP_AXIMM_49_AWLEN;
            assign ap_AWSIZE[49] = AP_AXIMM_49_AWSIZE;
            assign ap_AWBURST[49] = AP_AXIMM_49_AWBURST;
            assign ap_AWLOCK[49] = AP_AXIMM_49_AWLOCK;
            assign ap_AWCACHE[49] = AP_AXIMM_49_AWCACHE;
            assign ap_AWPROT[49] = AP_AXIMM_49_AWPROT;
            assign ap_AWREGION[49] = AP_AXIMM_49_AWREGION;
            assign ap_AWQOS[49] = AP_AXIMM_49_AWQOS;
            assign ap_AWVALID[49] = AP_AXIMM_49_AWVALID;
            assign AP_AXIMM_49_AWREADY = ap_AWREADY[49];
            assign ap_WDATA[49][M_AXIMM_49_DATA_WIDTH-1:0] = AP_AXIMM_49_WDATA;
            assign ap_WSTRB[49][M_AXIMM_49_DATA_WIDTH/8-1:0] = AP_AXIMM_49_WSTRB;
            assign ap_WLAST[49] = AP_AXIMM_49_WLAST;
            assign ap_WVALID[49] = AP_AXIMM_49_WVALID;
            assign AP_AXIMM_49_WREADY = ap_WREADY[49];
            assign AP_AXIMM_49_BRESP = ap_BRESP[49];
            assign AP_AXIMM_49_BVALID = ap_BVALID[49];
            assign ap_BREADY[49] = AP_AXIMM_49_BREADY;
            assign ap_ARADDR[49][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_49_ARADDR;
            assign ap_ARLEN[49] = AP_AXIMM_49_ARLEN;
            assign ap_ARSIZE[49] = AP_AXIMM_49_ARSIZE;
            assign ap_ARBURST[49] = AP_AXIMM_49_ARBURST;
            assign ap_ARLOCK[49] = AP_AXIMM_49_ARLOCK;
            assign ap_ARCACHE[49] = AP_AXIMM_49_ARCACHE;
            assign ap_ARPROT[49] = AP_AXIMM_49_ARPROT;
            assign ap_ARREGION[49] = AP_AXIMM_49_ARREGION;
            assign ap_ARQOS[49] = AP_AXIMM_49_ARQOS;
            assign ap_ARVALID[49] = AP_AXIMM_49_ARVALID;
            assign AP_AXIMM_49_ARREADY = ap_ARREADY[49];
            assign AP_AXIMM_49_RDATA = ap_RDATA[49][M_AXIMM_49_DATA_WIDTH-1:0];
            assign AP_AXIMM_49_RRESP = ap_RRESP[49];
            assign AP_AXIMM_49_RLAST = ap_RLAST[49];
            assign AP_AXIMM_49_RVALID = ap_RVALID[49];
            assign ap_RREADY[49] = AP_AXIMM_49_RREADY;
            assign M_AXIMM_49_AWADDR = dm_AWADDR[49][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_49_AWLEN = dm_AWLEN[49];
            assign M_AXIMM_49_AWSIZE = dm_AWSIZE[49];
            assign M_AXIMM_49_AWBURST = dm_AWBURST[49];
            assign M_AXIMM_49_AWLOCK = dm_AWLOCK[49];
            assign M_AXIMM_49_AWCACHE = dm_AWCACHE[49];
            assign M_AXIMM_49_AWPROT = dm_AWPROT[49];
            assign M_AXIMM_49_AWREGION = dm_AWREGION[49];
            assign M_AXIMM_49_AWQOS = dm_AWQOS[49];
            assign M_AXIMM_49_AWVALID = dm_AWVALID[49];
            assign dm_AWREADY[49] = M_AXIMM_49_AWREADY;
            assign M_AXIMM_49_WDATA = dm_WDATA[49][M_AXIMM_49_DATA_WIDTH-1:0];
            assign M_AXIMM_49_WSTRB = dm_WSTRB[49][M_AXIMM_49_DATA_WIDTH/8-1:0];
            assign M_AXIMM_49_WLAST = dm_WLAST[49];
            assign M_AXIMM_49_WVALID = dm_WVALID[49];
            assign dm_WREADY[49] = M_AXIMM_49_WREADY;
            assign dm_BRESP[49] = M_AXIMM_49_BRESP;
            assign dm_BVALID[49] = M_AXIMM_49_BVALID;
            assign M_AXIMM_49_BREADY = dm_BREADY[49];
            assign M_AXIMM_49_ARADDR = dm_ARADDR[49][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_49_ARLEN = dm_ARLEN[49];
            assign M_AXIMM_49_ARSIZE = dm_ARSIZE[49];
            assign M_AXIMM_49_ARBURST = dm_ARBURST[49];
            assign M_AXIMM_49_ARLOCK = dm_ARLOCK[49];
            assign M_AXIMM_49_ARCACHE = dm_ARCACHE[49];
            assign M_AXIMM_49_ARPROT = dm_ARPROT[49];
            assign M_AXIMM_49_ARREGION = dm_ARREGION[49];
            assign M_AXIMM_49_ARQOS = dm_ARQOS[49];
            assign M_AXIMM_49_ARVALID = dm_ARVALID[49];
            assign dm_ARREADY[49] = M_AXIMM_49_ARREADY;
            assign dm_RDATA[49][M_AXIMM_49_DATA_WIDTH-1:0] = M_AXIMM_49_RDATA;
            assign dm_RRESP[49] = M_AXIMM_49_RRESP;
            assign dm_RLAST[49] = M_AXIMM_49_RLAST;
            assign dm_RVALID[49] = M_AXIMM_49_RVALID;
            assign M_AXIMM_49_RREADY = dm_RREADY[49];
        end
        if(C_NUM_AXIMMs > 50) begin
            assign ap_AWADDR[50][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_50_AWADDR;
            assign ap_AWLEN[50] = AP_AXIMM_50_AWLEN;
            assign ap_AWSIZE[50] = AP_AXIMM_50_AWSIZE;
            assign ap_AWBURST[50] = AP_AXIMM_50_AWBURST;
            assign ap_AWLOCK[50] = AP_AXIMM_50_AWLOCK;
            assign ap_AWCACHE[50] = AP_AXIMM_50_AWCACHE;
            assign ap_AWPROT[50] = AP_AXIMM_50_AWPROT;
            assign ap_AWREGION[50] = AP_AXIMM_50_AWREGION;
            assign ap_AWQOS[50] = AP_AXIMM_50_AWQOS;
            assign ap_AWVALID[50] = AP_AXIMM_50_AWVALID;
            assign AP_AXIMM_50_AWREADY = ap_AWREADY[50];
            assign ap_WDATA[50][M_AXIMM_50_DATA_WIDTH-1:0] = AP_AXIMM_50_WDATA;
            assign ap_WSTRB[50][M_AXIMM_50_DATA_WIDTH/8-1:0] = AP_AXIMM_50_WSTRB;
            assign ap_WLAST[50] = AP_AXIMM_50_WLAST;
            assign ap_WVALID[50] = AP_AXIMM_50_WVALID;
            assign AP_AXIMM_50_WREADY = ap_WREADY[50];
            assign AP_AXIMM_50_BRESP = ap_BRESP[50];
            assign AP_AXIMM_50_BVALID = ap_BVALID[50];
            assign ap_BREADY[50] = AP_AXIMM_50_BREADY;
            assign ap_ARADDR[50][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_50_ARADDR;
            assign ap_ARLEN[50] = AP_AXIMM_50_ARLEN;
            assign ap_ARSIZE[50] = AP_AXIMM_50_ARSIZE;
            assign ap_ARBURST[50] = AP_AXIMM_50_ARBURST;
            assign ap_ARLOCK[50] = AP_AXIMM_50_ARLOCK;
            assign ap_ARCACHE[50] = AP_AXIMM_50_ARCACHE;
            assign ap_ARPROT[50] = AP_AXIMM_50_ARPROT;
            assign ap_ARREGION[50] = AP_AXIMM_50_ARREGION;
            assign ap_ARQOS[50] = AP_AXIMM_50_ARQOS;
            assign ap_ARVALID[50] = AP_AXIMM_50_ARVALID;
            assign AP_AXIMM_50_ARREADY = ap_ARREADY[50];
            assign AP_AXIMM_50_RDATA = ap_RDATA[50][M_AXIMM_50_DATA_WIDTH-1:0];
            assign AP_AXIMM_50_RRESP = ap_RRESP[50];
            assign AP_AXIMM_50_RLAST = ap_RLAST[50];
            assign AP_AXIMM_50_RVALID = ap_RVALID[50];
            assign ap_RREADY[50] = AP_AXIMM_50_RREADY;
            assign M_AXIMM_50_AWADDR = dm_AWADDR[50][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_50_AWLEN = dm_AWLEN[50];
            assign M_AXIMM_50_AWSIZE = dm_AWSIZE[50];
            assign M_AXIMM_50_AWBURST = dm_AWBURST[50];
            assign M_AXIMM_50_AWLOCK = dm_AWLOCK[50];
            assign M_AXIMM_50_AWCACHE = dm_AWCACHE[50];
            assign M_AXIMM_50_AWPROT = dm_AWPROT[50];
            assign M_AXIMM_50_AWREGION = dm_AWREGION[50];
            assign M_AXIMM_50_AWQOS = dm_AWQOS[50];
            assign M_AXIMM_50_AWVALID = dm_AWVALID[50];
            assign dm_AWREADY[50] = M_AXIMM_50_AWREADY;
            assign M_AXIMM_50_WDATA = dm_WDATA[50][M_AXIMM_50_DATA_WIDTH-1:0];
            assign M_AXIMM_50_WSTRB = dm_WSTRB[50][M_AXIMM_50_DATA_WIDTH/8-1:0];
            assign M_AXIMM_50_WLAST = dm_WLAST[50];
            assign M_AXIMM_50_WVALID = dm_WVALID[50];
            assign dm_WREADY[50] = M_AXIMM_50_WREADY;
            assign dm_BRESP[50] = M_AXIMM_50_BRESP;
            assign dm_BVALID[50] = M_AXIMM_50_BVALID;
            assign M_AXIMM_50_BREADY = dm_BREADY[50];
            assign M_AXIMM_50_ARADDR = dm_ARADDR[50][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_50_ARLEN = dm_ARLEN[50];
            assign M_AXIMM_50_ARSIZE = dm_ARSIZE[50];
            assign M_AXIMM_50_ARBURST = dm_ARBURST[50];
            assign M_AXIMM_50_ARLOCK = dm_ARLOCK[50];
            assign M_AXIMM_50_ARCACHE = dm_ARCACHE[50];
            assign M_AXIMM_50_ARPROT = dm_ARPROT[50];
            assign M_AXIMM_50_ARREGION = dm_ARREGION[50];
            assign M_AXIMM_50_ARQOS = dm_ARQOS[50];
            assign M_AXIMM_50_ARVALID = dm_ARVALID[50];
            assign dm_ARREADY[50] = M_AXIMM_50_ARREADY;
            assign dm_RDATA[50][M_AXIMM_50_DATA_WIDTH-1:0] = M_AXIMM_50_RDATA;
            assign dm_RRESP[50] = M_AXIMM_50_RRESP;
            assign dm_RLAST[50] = M_AXIMM_50_RLAST;
            assign dm_RVALID[50] = M_AXIMM_50_RVALID;
            assign M_AXIMM_50_RREADY = dm_RREADY[50];
        end
        if(C_NUM_AXIMMs > 51) begin
            assign ap_AWADDR[51][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_51_AWADDR;
            assign ap_AWLEN[51] = AP_AXIMM_51_AWLEN;
            assign ap_AWSIZE[51] = AP_AXIMM_51_AWSIZE;
            assign ap_AWBURST[51] = AP_AXIMM_51_AWBURST;
            assign ap_AWLOCK[51] = AP_AXIMM_51_AWLOCK;
            assign ap_AWCACHE[51] = AP_AXIMM_51_AWCACHE;
            assign ap_AWPROT[51] = AP_AXIMM_51_AWPROT;
            assign ap_AWREGION[51] = AP_AXIMM_51_AWREGION;
            assign ap_AWQOS[51] = AP_AXIMM_51_AWQOS;
            assign ap_AWVALID[51] = AP_AXIMM_51_AWVALID;
            assign AP_AXIMM_51_AWREADY = ap_AWREADY[51];
            assign ap_WDATA[51][M_AXIMM_51_DATA_WIDTH-1:0] = AP_AXIMM_51_WDATA;
            assign ap_WSTRB[51][M_AXIMM_51_DATA_WIDTH/8-1:0] = AP_AXIMM_51_WSTRB;
            assign ap_WLAST[51] = AP_AXIMM_51_WLAST;
            assign ap_WVALID[51] = AP_AXIMM_51_WVALID;
            assign AP_AXIMM_51_WREADY = ap_WREADY[51];
            assign AP_AXIMM_51_BRESP = ap_BRESP[51];
            assign AP_AXIMM_51_BVALID = ap_BVALID[51];
            assign ap_BREADY[51] = AP_AXIMM_51_BREADY;
            assign ap_ARADDR[51][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_51_ARADDR;
            assign ap_ARLEN[51] = AP_AXIMM_51_ARLEN;
            assign ap_ARSIZE[51] = AP_AXIMM_51_ARSIZE;
            assign ap_ARBURST[51] = AP_AXIMM_51_ARBURST;
            assign ap_ARLOCK[51] = AP_AXIMM_51_ARLOCK;
            assign ap_ARCACHE[51] = AP_AXIMM_51_ARCACHE;
            assign ap_ARPROT[51] = AP_AXIMM_51_ARPROT;
            assign ap_ARREGION[51] = AP_AXIMM_51_ARREGION;
            assign ap_ARQOS[51] = AP_AXIMM_51_ARQOS;
            assign ap_ARVALID[51] = AP_AXIMM_51_ARVALID;
            assign AP_AXIMM_51_ARREADY = ap_ARREADY[51];
            assign AP_AXIMM_51_RDATA = ap_RDATA[51][M_AXIMM_51_DATA_WIDTH-1:0];
            assign AP_AXIMM_51_RRESP = ap_RRESP[51];
            assign AP_AXIMM_51_RLAST = ap_RLAST[51];
            assign AP_AXIMM_51_RVALID = ap_RVALID[51];
            assign ap_RREADY[51] = AP_AXIMM_51_RREADY;
            assign M_AXIMM_51_AWADDR = dm_AWADDR[51][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_51_AWLEN = dm_AWLEN[51];
            assign M_AXIMM_51_AWSIZE = dm_AWSIZE[51];
            assign M_AXIMM_51_AWBURST = dm_AWBURST[51];
            assign M_AXIMM_51_AWLOCK = dm_AWLOCK[51];
            assign M_AXIMM_51_AWCACHE = dm_AWCACHE[51];
            assign M_AXIMM_51_AWPROT = dm_AWPROT[51];
            assign M_AXIMM_51_AWREGION = dm_AWREGION[51];
            assign M_AXIMM_51_AWQOS = dm_AWQOS[51];
            assign M_AXIMM_51_AWVALID = dm_AWVALID[51];
            assign dm_AWREADY[51] = M_AXIMM_51_AWREADY;
            assign M_AXIMM_51_WDATA = dm_WDATA[51][M_AXIMM_51_DATA_WIDTH-1:0];
            assign M_AXIMM_51_WSTRB = dm_WSTRB[51][M_AXIMM_51_DATA_WIDTH/8-1:0];
            assign M_AXIMM_51_WLAST = dm_WLAST[51];
            assign M_AXIMM_51_WVALID = dm_WVALID[51];
            assign dm_WREADY[51] = M_AXIMM_51_WREADY;
            assign dm_BRESP[51] = M_AXIMM_51_BRESP;
            assign dm_BVALID[51] = M_AXIMM_51_BVALID;
            assign M_AXIMM_51_BREADY = dm_BREADY[51];
            assign M_AXIMM_51_ARADDR = dm_ARADDR[51][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_51_ARLEN = dm_ARLEN[51];
            assign M_AXIMM_51_ARSIZE = dm_ARSIZE[51];
            assign M_AXIMM_51_ARBURST = dm_ARBURST[51];
            assign M_AXIMM_51_ARLOCK = dm_ARLOCK[51];
            assign M_AXIMM_51_ARCACHE = dm_ARCACHE[51];
            assign M_AXIMM_51_ARPROT = dm_ARPROT[51];
            assign M_AXIMM_51_ARREGION = dm_ARREGION[51];
            assign M_AXIMM_51_ARQOS = dm_ARQOS[51];
            assign M_AXIMM_51_ARVALID = dm_ARVALID[51];
            assign dm_ARREADY[51] = M_AXIMM_51_ARREADY;
            assign dm_RDATA[51][M_AXIMM_51_DATA_WIDTH-1:0] = M_AXIMM_51_RDATA;
            assign dm_RRESP[51] = M_AXIMM_51_RRESP;
            assign dm_RLAST[51] = M_AXIMM_51_RLAST;
            assign dm_RVALID[51] = M_AXIMM_51_RVALID;
            assign M_AXIMM_51_RREADY = dm_RREADY[51];
        end
        if(C_NUM_AXIMMs > 52) begin
            assign ap_AWADDR[52][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_52_AWADDR;
            assign ap_AWLEN[52] = AP_AXIMM_52_AWLEN;
            assign ap_AWSIZE[52] = AP_AXIMM_52_AWSIZE;
            assign ap_AWBURST[52] = AP_AXIMM_52_AWBURST;
            assign ap_AWLOCK[52] = AP_AXIMM_52_AWLOCK;
            assign ap_AWCACHE[52] = AP_AXIMM_52_AWCACHE;
            assign ap_AWPROT[52] = AP_AXIMM_52_AWPROT;
            assign ap_AWREGION[52] = AP_AXIMM_52_AWREGION;
            assign ap_AWQOS[52] = AP_AXIMM_52_AWQOS;
            assign ap_AWVALID[52] = AP_AXIMM_52_AWVALID;
            assign AP_AXIMM_52_AWREADY = ap_AWREADY[52];
            assign ap_WDATA[52][M_AXIMM_52_DATA_WIDTH-1:0] = AP_AXIMM_52_WDATA;
            assign ap_WSTRB[52][M_AXIMM_52_DATA_WIDTH/8-1:0] = AP_AXIMM_52_WSTRB;
            assign ap_WLAST[52] = AP_AXIMM_52_WLAST;
            assign ap_WVALID[52] = AP_AXIMM_52_WVALID;
            assign AP_AXIMM_52_WREADY = ap_WREADY[52];
            assign AP_AXIMM_52_BRESP = ap_BRESP[52];
            assign AP_AXIMM_52_BVALID = ap_BVALID[52];
            assign ap_BREADY[52] = AP_AXIMM_52_BREADY;
            assign ap_ARADDR[52][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_52_ARADDR;
            assign ap_ARLEN[52] = AP_AXIMM_52_ARLEN;
            assign ap_ARSIZE[52] = AP_AXIMM_52_ARSIZE;
            assign ap_ARBURST[52] = AP_AXIMM_52_ARBURST;
            assign ap_ARLOCK[52] = AP_AXIMM_52_ARLOCK;
            assign ap_ARCACHE[52] = AP_AXIMM_52_ARCACHE;
            assign ap_ARPROT[52] = AP_AXIMM_52_ARPROT;
            assign ap_ARREGION[52] = AP_AXIMM_52_ARREGION;
            assign ap_ARQOS[52] = AP_AXIMM_52_ARQOS;
            assign ap_ARVALID[52] = AP_AXIMM_52_ARVALID;
            assign AP_AXIMM_52_ARREADY = ap_ARREADY[52];
            assign AP_AXIMM_52_RDATA = ap_RDATA[52][M_AXIMM_52_DATA_WIDTH-1:0];
            assign AP_AXIMM_52_RRESP = ap_RRESP[52];
            assign AP_AXIMM_52_RLAST = ap_RLAST[52];
            assign AP_AXIMM_52_RVALID = ap_RVALID[52];
            assign ap_RREADY[52] = AP_AXIMM_52_RREADY;
            assign M_AXIMM_52_AWADDR = dm_AWADDR[52][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_52_AWLEN = dm_AWLEN[52];
            assign M_AXIMM_52_AWSIZE = dm_AWSIZE[52];
            assign M_AXIMM_52_AWBURST = dm_AWBURST[52];
            assign M_AXIMM_52_AWLOCK = dm_AWLOCK[52];
            assign M_AXIMM_52_AWCACHE = dm_AWCACHE[52];
            assign M_AXIMM_52_AWPROT = dm_AWPROT[52];
            assign M_AXIMM_52_AWREGION = dm_AWREGION[52];
            assign M_AXIMM_52_AWQOS = dm_AWQOS[52];
            assign M_AXIMM_52_AWVALID = dm_AWVALID[52];
            assign dm_AWREADY[52] = M_AXIMM_52_AWREADY;
            assign M_AXIMM_52_WDATA = dm_WDATA[52][M_AXIMM_52_DATA_WIDTH-1:0];
            assign M_AXIMM_52_WSTRB = dm_WSTRB[52][M_AXIMM_52_DATA_WIDTH/8-1:0];
            assign M_AXIMM_52_WLAST = dm_WLAST[52];
            assign M_AXIMM_52_WVALID = dm_WVALID[52];
            assign dm_WREADY[52] = M_AXIMM_52_WREADY;
            assign dm_BRESP[52] = M_AXIMM_52_BRESP;
            assign dm_BVALID[52] = M_AXIMM_52_BVALID;
            assign M_AXIMM_52_BREADY = dm_BREADY[52];
            assign M_AXIMM_52_ARADDR = dm_ARADDR[52][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_52_ARLEN = dm_ARLEN[52];
            assign M_AXIMM_52_ARSIZE = dm_ARSIZE[52];
            assign M_AXIMM_52_ARBURST = dm_ARBURST[52];
            assign M_AXIMM_52_ARLOCK = dm_ARLOCK[52];
            assign M_AXIMM_52_ARCACHE = dm_ARCACHE[52];
            assign M_AXIMM_52_ARPROT = dm_ARPROT[52];
            assign M_AXIMM_52_ARREGION = dm_ARREGION[52];
            assign M_AXIMM_52_ARQOS = dm_ARQOS[52];
            assign M_AXIMM_52_ARVALID = dm_ARVALID[52];
            assign dm_ARREADY[52] = M_AXIMM_52_ARREADY;
            assign dm_RDATA[52][M_AXIMM_52_DATA_WIDTH-1:0] = M_AXIMM_52_RDATA;
            assign dm_RRESP[52] = M_AXIMM_52_RRESP;
            assign dm_RLAST[52] = M_AXIMM_52_RLAST;
            assign dm_RVALID[52] = M_AXIMM_52_RVALID;
            assign M_AXIMM_52_RREADY = dm_RREADY[52];
        end
        if(C_NUM_AXIMMs > 53) begin
            assign ap_AWADDR[53][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_53_AWADDR;
            assign ap_AWLEN[53] = AP_AXIMM_53_AWLEN;
            assign ap_AWSIZE[53] = AP_AXIMM_53_AWSIZE;
            assign ap_AWBURST[53] = AP_AXIMM_53_AWBURST;
            assign ap_AWLOCK[53] = AP_AXIMM_53_AWLOCK;
            assign ap_AWCACHE[53] = AP_AXIMM_53_AWCACHE;
            assign ap_AWPROT[53] = AP_AXIMM_53_AWPROT;
            assign ap_AWREGION[53] = AP_AXIMM_53_AWREGION;
            assign ap_AWQOS[53] = AP_AXIMM_53_AWQOS;
            assign ap_AWVALID[53] = AP_AXIMM_53_AWVALID;
            assign AP_AXIMM_53_AWREADY = ap_AWREADY[53];
            assign ap_WDATA[53][M_AXIMM_53_DATA_WIDTH-1:0] = AP_AXIMM_53_WDATA;
            assign ap_WSTRB[53][M_AXIMM_53_DATA_WIDTH/8-1:0] = AP_AXIMM_53_WSTRB;
            assign ap_WLAST[53] = AP_AXIMM_53_WLAST;
            assign ap_WVALID[53] = AP_AXIMM_53_WVALID;
            assign AP_AXIMM_53_WREADY = ap_WREADY[53];
            assign AP_AXIMM_53_BRESP = ap_BRESP[53];
            assign AP_AXIMM_53_BVALID = ap_BVALID[53];
            assign ap_BREADY[53] = AP_AXIMM_53_BREADY;
            assign ap_ARADDR[53][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_53_ARADDR;
            assign ap_ARLEN[53] = AP_AXIMM_53_ARLEN;
            assign ap_ARSIZE[53] = AP_AXIMM_53_ARSIZE;
            assign ap_ARBURST[53] = AP_AXIMM_53_ARBURST;
            assign ap_ARLOCK[53] = AP_AXIMM_53_ARLOCK;
            assign ap_ARCACHE[53] = AP_AXIMM_53_ARCACHE;
            assign ap_ARPROT[53] = AP_AXIMM_53_ARPROT;
            assign ap_ARREGION[53] = AP_AXIMM_53_ARREGION;
            assign ap_ARQOS[53] = AP_AXIMM_53_ARQOS;
            assign ap_ARVALID[53] = AP_AXIMM_53_ARVALID;
            assign AP_AXIMM_53_ARREADY = ap_ARREADY[53];
            assign AP_AXIMM_53_RDATA = ap_RDATA[53][M_AXIMM_53_DATA_WIDTH-1:0];
            assign AP_AXIMM_53_RRESP = ap_RRESP[53];
            assign AP_AXIMM_53_RLAST = ap_RLAST[53];
            assign AP_AXIMM_53_RVALID = ap_RVALID[53];
            assign ap_RREADY[53] = AP_AXIMM_53_RREADY;
            assign M_AXIMM_53_AWADDR = dm_AWADDR[53][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_53_AWLEN = dm_AWLEN[53];
            assign M_AXIMM_53_AWSIZE = dm_AWSIZE[53];
            assign M_AXIMM_53_AWBURST = dm_AWBURST[53];
            assign M_AXIMM_53_AWLOCK = dm_AWLOCK[53];
            assign M_AXIMM_53_AWCACHE = dm_AWCACHE[53];
            assign M_AXIMM_53_AWPROT = dm_AWPROT[53];
            assign M_AXIMM_53_AWREGION = dm_AWREGION[53];
            assign M_AXIMM_53_AWQOS = dm_AWQOS[53];
            assign M_AXIMM_53_AWVALID = dm_AWVALID[53];
            assign dm_AWREADY[53] = M_AXIMM_53_AWREADY;
            assign M_AXIMM_53_WDATA = dm_WDATA[53][M_AXIMM_53_DATA_WIDTH-1:0];
            assign M_AXIMM_53_WSTRB = dm_WSTRB[53][M_AXIMM_53_DATA_WIDTH/8-1:0];
            assign M_AXIMM_53_WLAST = dm_WLAST[53];
            assign M_AXIMM_53_WVALID = dm_WVALID[53];
            assign dm_WREADY[53] = M_AXIMM_53_WREADY;
            assign dm_BRESP[53] = M_AXIMM_53_BRESP;
            assign dm_BVALID[53] = M_AXIMM_53_BVALID;
            assign M_AXIMM_53_BREADY = dm_BREADY[53];
            assign M_AXIMM_53_ARADDR = dm_ARADDR[53][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_53_ARLEN = dm_ARLEN[53];
            assign M_AXIMM_53_ARSIZE = dm_ARSIZE[53];
            assign M_AXIMM_53_ARBURST = dm_ARBURST[53];
            assign M_AXIMM_53_ARLOCK = dm_ARLOCK[53];
            assign M_AXIMM_53_ARCACHE = dm_ARCACHE[53];
            assign M_AXIMM_53_ARPROT = dm_ARPROT[53];
            assign M_AXIMM_53_ARREGION = dm_ARREGION[53];
            assign M_AXIMM_53_ARQOS = dm_ARQOS[53];
            assign M_AXIMM_53_ARVALID = dm_ARVALID[53];
            assign dm_ARREADY[53] = M_AXIMM_53_ARREADY;
            assign dm_RDATA[53][M_AXIMM_53_DATA_WIDTH-1:0] = M_AXIMM_53_RDATA;
            assign dm_RRESP[53] = M_AXIMM_53_RRESP;
            assign dm_RLAST[53] = M_AXIMM_53_RLAST;
            assign dm_RVALID[53] = M_AXIMM_53_RVALID;
            assign M_AXIMM_53_RREADY = dm_RREADY[53];
        end
        if(C_NUM_AXIMMs > 54) begin
            assign ap_AWADDR[54][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_54_AWADDR;
            assign ap_AWLEN[54] = AP_AXIMM_54_AWLEN;
            assign ap_AWSIZE[54] = AP_AXIMM_54_AWSIZE;
            assign ap_AWBURST[54] = AP_AXIMM_54_AWBURST;
            assign ap_AWLOCK[54] = AP_AXIMM_54_AWLOCK;
            assign ap_AWCACHE[54] = AP_AXIMM_54_AWCACHE;
            assign ap_AWPROT[54] = AP_AXIMM_54_AWPROT;
            assign ap_AWREGION[54] = AP_AXIMM_54_AWREGION;
            assign ap_AWQOS[54] = AP_AXIMM_54_AWQOS;
            assign ap_AWVALID[54] = AP_AXIMM_54_AWVALID;
            assign AP_AXIMM_54_AWREADY = ap_AWREADY[54];
            assign ap_WDATA[54][M_AXIMM_54_DATA_WIDTH-1:0] = AP_AXIMM_54_WDATA;
            assign ap_WSTRB[54][M_AXIMM_54_DATA_WIDTH/8-1:0] = AP_AXIMM_54_WSTRB;
            assign ap_WLAST[54] = AP_AXIMM_54_WLAST;
            assign ap_WVALID[54] = AP_AXIMM_54_WVALID;
            assign AP_AXIMM_54_WREADY = ap_WREADY[54];
            assign AP_AXIMM_54_BRESP = ap_BRESP[54];
            assign AP_AXIMM_54_BVALID = ap_BVALID[54];
            assign ap_BREADY[54] = AP_AXIMM_54_BREADY;
            assign ap_ARADDR[54][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_54_ARADDR;
            assign ap_ARLEN[54] = AP_AXIMM_54_ARLEN;
            assign ap_ARSIZE[54] = AP_AXIMM_54_ARSIZE;
            assign ap_ARBURST[54] = AP_AXIMM_54_ARBURST;
            assign ap_ARLOCK[54] = AP_AXIMM_54_ARLOCK;
            assign ap_ARCACHE[54] = AP_AXIMM_54_ARCACHE;
            assign ap_ARPROT[54] = AP_AXIMM_54_ARPROT;
            assign ap_ARREGION[54] = AP_AXIMM_54_ARREGION;
            assign ap_ARQOS[54] = AP_AXIMM_54_ARQOS;
            assign ap_ARVALID[54] = AP_AXIMM_54_ARVALID;
            assign AP_AXIMM_54_ARREADY = ap_ARREADY[54];
            assign AP_AXIMM_54_RDATA = ap_RDATA[54][M_AXIMM_54_DATA_WIDTH-1:0];
            assign AP_AXIMM_54_RRESP = ap_RRESP[54];
            assign AP_AXIMM_54_RLAST = ap_RLAST[54];
            assign AP_AXIMM_54_RVALID = ap_RVALID[54];
            assign ap_RREADY[54] = AP_AXIMM_54_RREADY;
            assign M_AXIMM_54_AWADDR = dm_AWADDR[54][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_54_AWLEN = dm_AWLEN[54];
            assign M_AXIMM_54_AWSIZE = dm_AWSIZE[54];
            assign M_AXIMM_54_AWBURST = dm_AWBURST[54];
            assign M_AXIMM_54_AWLOCK = dm_AWLOCK[54];
            assign M_AXIMM_54_AWCACHE = dm_AWCACHE[54];
            assign M_AXIMM_54_AWPROT = dm_AWPROT[54];
            assign M_AXIMM_54_AWREGION = dm_AWREGION[54];
            assign M_AXIMM_54_AWQOS = dm_AWQOS[54];
            assign M_AXIMM_54_AWVALID = dm_AWVALID[54];
            assign dm_AWREADY[54] = M_AXIMM_54_AWREADY;
            assign M_AXIMM_54_WDATA = dm_WDATA[54][M_AXIMM_54_DATA_WIDTH-1:0];
            assign M_AXIMM_54_WSTRB = dm_WSTRB[54][M_AXIMM_54_DATA_WIDTH/8-1:0];
            assign M_AXIMM_54_WLAST = dm_WLAST[54];
            assign M_AXIMM_54_WVALID = dm_WVALID[54];
            assign dm_WREADY[54] = M_AXIMM_54_WREADY;
            assign dm_BRESP[54] = M_AXIMM_54_BRESP;
            assign dm_BVALID[54] = M_AXIMM_54_BVALID;
            assign M_AXIMM_54_BREADY = dm_BREADY[54];
            assign M_AXIMM_54_ARADDR = dm_ARADDR[54][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_54_ARLEN = dm_ARLEN[54];
            assign M_AXIMM_54_ARSIZE = dm_ARSIZE[54];
            assign M_AXIMM_54_ARBURST = dm_ARBURST[54];
            assign M_AXIMM_54_ARLOCK = dm_ARLOCK[54];
            assign M_AXIMM_54_ARCACHE = dm_ARCACHE[54];
            assign M_AXIMM_54_ARPROT = dm_ARPROT[54];
            assign M_AXIMM_54_ARREGION = dm_ARREGION[54];
            assign M_AXIMM_54_ARQOS = dm_ARQOS[54];
            assign M_AXIMM_54_ARVALID = dm_ARVALID[54];
            assign dm_ARREADY[54] = M_AXIMM_54_ARREADY;
            assign dm_RDATA[54][M_AXIMM_54_DATA_WIDTH-1:0] = M_AXIMM_54_RDATA;
            assign dm_RRESP[54] = M_AXIMM_54_RRESP;
            assign dm_RLAST[54] = M_AXIMM_54_RLAST;
            assign dm_RVALID[54] = M_AXIMM_54_RVALID;
            assign M_AXIMM_54_RREADY = dm_RREADY[54];
        end
        if(C_NUM_AXIMMs > 55) begin
            assign ap_AWADDR[55][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_55_AWADDR;
            assign ap_AWLEN[55] = AP_AXIMM_55_AWLEN;
            assign ap_AWSIZE[55] = AP_AXIMM_55_AWSIZE;
            assign ap_AWBURST[55] = AP_AXIMM_55_AWBURST;
            assign ap_AWLOCK[55] = AP_AXIMM_55_AWLOCK;
            assign ap_AWCACHE[55] = AP_AXIMM_55_AWCACHE;
            assign ap_AWPROT[55] = AP_AXIMM_55_AWPROT;
            assign ap_AWREGION[55] = AP_AXIMM_55_AWREGION;
            assign ap_AWQOS[55] = AP_AXIMM_55_AWQOS;
            assign ap_AWVALID[55] = AP_AXIMM_55_AWVALID;
            assign AP_AXIMM_55_AWREADY = ap_AWREADY[55];
            assign ap_WDATA[55][M_AXIMM_55_DATA_WIDTH-1:0] = AP_AXIMM_55_WDATA;
            assign ap_WSTRB[55][M_AXIMM_55_DATA_WIDTH/8-1:0] = AP_AXIMM_55_WSTRB;
            assign ap_WLAST[55] = AP_AXIMM_55_WLAST;
            assign ap_WVALID[55] = AP_AXIMM_55_WVALID;
            assign AP_AXIMM_55_WREADY = ap_WREADY[55];
            assign AP_AXIMM_55_BRESP = ap_BRESP[55];
            assign AP_AXIMM_55_BVALID = ap_BVALID[55];
            assign ap_BREADY[55] = AP_AXIMM_55_BREADY;
            assign ap_ARADDR[55][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_55_ARADDR;
            assign ap_ARLEN[55] = AP_AXIMM_55_ARLEN;
            assign ap_ARSIZE[55] = AP_AXIMM_55_ARSIZE;
            assign ap_ARBURST[55] = AP_AXIMM_55_ARBURST;
            assign ap_ARLOCK[55] = AP_AXIMM_55_ARLOCK;
            assign ap_ARCACHE[55] = AP_AXIMM_55_ARCACHE;
            assign ap_ARPROT[55] = AP_AXIMM_55_ARPROT;
            assign ap_ARREGION[55] = AP_AXIMM_55_ARREGION;
            assign ap_ARQOS[55] = AP_AXIMM_55_ARQOS;
            assign ap_ARVALID[55] = AP_AXIMM_55_ARVALID;
            assign AP_AXIMM_55_ARREADY = ap_ARREADY[55];
            assign AP_AXIMM_55_RDATA = ap_RDATA[55][M_AXIMM_55_DATA_WIDTH-1:0];
            assign AP_AXIMM_55_RRESP = ap_RRESP[55];
            assign AP_AXIMM_55_RLAST = ap_RLAST[55];
            assign AP_AXIMM_55_RVALID = ap_RVALID[55];
            assign ap_RREADY[55] = AP_AXIMM_55_RREADY;
            assign M_AXIMM_55_AWADDR = dm_AWADDR[55][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_55_AWLEN = dm_AWLEN[55];
            assign M_AXIMM_55_AWSIZE = dm_AWSIZE[55];
            assign M_AXIMM_55_AWBURST = dm_AWBURST[55];
            assign M_AXIMM_55_AWLOCK = dm_AWLOCK[55];
            assign M_AXIMM_55_AWCACHE = dm_AWCACHE[55];
            assign M_AXIMM_55_AWPROT = dm_AWPROT[55];
            assign M_AXIMM_55_AWREGION = dm_AWREGION[55];
            assign M_AXIMM_55_AWQOS = dm_AWQOS[55];
            assign M_AXIMM_55_AWVALID = dm_AWVALID[55];
            assign dm_AWREADY[55] = M_AXIMM_55_AWREADY;
            assign M_AXIMM_55_WDATA = dm_WDATA[55][M_AXIMM_55_DATA_WIDTH-1:0];
            assign M_AXIMM_55_WSTRB = dm_WSTRB[55][M_AXIMM_55_DATA_WIDTH/8-1:0];
            assign M_AXIMM_55_WLAST = dm_WLAST[55];
            assign M_AXIMM_55_WVALID = dm_WVALID[55];
            assign dm_WREADY[55] = M_AXIMM_55_WREADY;
            assign dm_BRESP[55] = M_AXIMM_55_BRESP;
            assign dm_BVALID[55] = M_AXIMM_55_BVALID;
            assign M_AXIMM_55_BREADY = dm_BREADY[55];
            assign M_AXIMM_55_ARADDR = dm_ARADDR[55][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_55_ARLEN = dm_ARLEN[55];
            assign M_AXIMM_55_ARSIZE = dm_ARSIZE[55];
            assign M_AXIMM_55_ARBURST = dm_ARBURST[55];
            assign M_AXIMM_55_ARLOCK = dm_ARLOCK[55];
            assign M_AXIMM_55_ARCACHE = dm_ARCACHE[55];
            assign M_AXIMM_55_ARPROT = dm_ARPROT[55];
            assign M_AXIMM_55_ARREGION = dm_ARREGION[55];
            assign M_AXIMM_55_ARQOS = dm_ARQOS[55];
            assign M_AXIMM_55_ARVALID = dm_ARVALID[55];
            assign dm_ARREADY[55] = M_AXIMM_55_ARREADY;
            assign dm_RDATA[55][M_AXIMM_55_DATA_WIDTH-1:0] = M_AXIMM_55_RDATA;
            assign dm_RRESP[55] = M_AXIMM_55_RRESP;
            assign dm_RLAST[55] = M_AXIMM_55_RLAST;
            assign dm_RVALID[55] = M_AXIMM_55_RVALID;
            assign M_AXIMM_55_RREADY = dm_RREADY[55];
        end
        if(C_NUM_AXIMMs > 56) begin
            assign ap_AWADDR[56][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_56_AWADDR;
            assign ap_AWLEN[56] = AP_AXIMM_56_AWLEN;
            assign ap_AWSIZE[56] = AP_AXIMM_56_AWSIZE;
            assign ap_AWBURST[56] = AP_AXIMM_56_AWBURST;
            assign ap_AWLOCK[56] = AP_AXIMM_56_AWLOCK;
            assign ap_AWCACHE[56] = AP_AXIMM_56_AWCACHE;
            assign ap_AWPROT[56] = AP_AXIMM_56_AWPROT;
            assign ap_AWREGION[56] = AP_AXIMM_56_AWREGION;
            assign ap_AWQOS[56] = AP_AXIMM_56_AWQOS;
            assign ap_AWVALID[56] = AP_AXIMM_56_AWVALID;
            assign AP_AXIMM_56_AWREADY = ap_AWREADY[56];
            assign ap_WDATA[56][M_AXIMM_56_DATA_WIDTH-1:0] = AP_AXIMM_56_WDATA;
            assign ap_WSTRB[56][M_AXIMM_56_DATA_WIDTH/8-1:0] = AP_AXIMM_56_WSTRB;
            assign ap_WLAST[56] = AP_AXIMM_56_WLAST;
            assign ap_WVALID[56] = AP_AXIMM_56_WVALID;
            assign AP_AXIMM_56_WREADY = ap_WREADY[56];
            assign AP_AXIMM_56_BRESP = ap_BRESP[56];
            assign AP_AXIMM_56_BVALID = ap_BVALID[56];
            assign ap_BREADY[56] = AP_AXIMM_56_BREADY;
            assign ap_ARADDR[56][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_56_ARADDR;
            assign ap_ARLEN[56] = AP_AXIMM_56_ARLEN;
            assign ap_ARSIZE[56] = AP_AXIMM_56_ARSIZE;
            assign ap_ARBURST[56] = AP_AXIMM_56_ARBURST;
            assign ap_ARLOCK[56] = AP_AXIMM_56_ARLOCK;
            assign ap_ARCACHE[56] = AP_AXIMM_56_ARCACHE;
            assign ap_ARPROT[56] = AP_AXIMM_56_ARPROT;
            assign ap_ARREGION[56] = AP_AXIMM_56_ARREGION;
            assign ap_ARQOS[56] = AP_AXIMM_56_ARQOS;
            assign ap_ARVALID[56] = AP_AXIMM_56_ARVALID;
            assign AP_AXIMM_56_ARREADY = ap_ARREADY[56];
            assign AP_AXIMM_56_RDATA = ap_RDATA[56][M_AXIMM_56_DATA_WIDTH-1:0];
            assign AP_AXIMM_56_RRESP = ap_RRESP[56];
            assign AP_AXIMM_56_RLAST = ap_RLAST[56];
            assign AP_AXIMM_56_RVALID = ap_RVALID[56];
            assign ap_RREADY[56] = AP_AXIMM_56_RREADY;
            assign M_AXIMM_56_AWADDR = dm_AWADDR[56][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_56_AWLEN = dm_AWLEN[56];
            assign M_AXIMM_56_AWSIZE = dm_AWSIZE[56];
            assign M_AXIMM_56_AWBURST = dm_AWBURST[56];
            assign M_AXIMM_56_AWLOCK = dm_AWLOCK[56];
            assign M_AXIMM_56_AWCACHE = dm_AWCACHE[56];
            assign M_AXIMM_56_AWPROT = dm_AWPROT[56];
            assign M_AXIMM_56_AWREGION = dm_AWREGION[56];
            assign M_AXIMM_56_AWQOS = dm_AWQOS[56];
            assign M_AXIMM_56_AWVALID = dm_AWVALID[56];
            assign dm_AWREADY[56] = M_AXIMM_56_AWREADY;
            assign M_AXIMM_56_WDATA = dm_WDATA[56][M_AXIMM_56_DATA_WIDTH-1:0];
            assign M_AXIMM_56_WSTRB = dm_WSTRB[56][M_AXIMM_56_DATA_WIDTH/8-1:0];
            assign M_AXIMM_56_WLAST = dm_WLAST[56];
            assign M_AXIMM_56_WVALID = dm_WVALID[56];
            assign dm_WREADY[56] = M_AXIMM_56_WREADY;
            assign dm_BRESP[56] = M_AXIMM_56_BRESP;
            assign dm_BVALID[56] = M_AXIMM_56_BVALID;
            assign M_AXIMM_56_BREADY = dm_BREADY[56];
            assign M_AXIMM_56_ARADDR = dm_ARADDR[56][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_56_ARLEN = dm_ARLEN[56];
            assign M_AXIMM_56_ARSIZE = dm_ARSIZE[56];
            assign M_AXIMM_56_ARBURST = dm_ARBURST[56];
            assign M_AXIMM_56_ARLOCK = dm_ARLOCK[56];
            assign M_AXIMM_56_ARCACHE = dm_ARCACHE[56];
            assign M_AXIMM_56_ARPROT = dm_ARPROT[56];
            assign M_AXIMM_56_ARREGION = dm_ARREGION[56];
            assign M_AXIMM_56_ARQOS = dm_ARQOS[56];
            assign M_AXIMM_56_ARVALID = dm_ARVALID[56];
            assign dm_ARREADY[56] = M_AXIMM_56_ARREADY;
            assign dm_RDATA[56][M_AXIMM_56_DATA_WIDTH-1:0] = M_AXIMM_56_RDATA;
            assign dm_RRESP[56] = M_AXIMM_56_RRESP;
            assign dm_RLAST[56] = M_AXIMM_56_RLAST;
            assign dm_RVALID[56] = M_AXIMM_56_RVALID;
            assign M_AXIMM_56_RREADY = dm_RREADY[56];
        end
        if(C_NUM_AXIMMs > 57) begin
            assign ap_AWADDR[57][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_57_AWADDR;
            assign ap_AWLEN[57] = AP_AXIMM_57_AWLEN;
            assign ap_AWSIZE[57] = AP_AXIMM_57_AWSIZE;
            assign ap_AWBURST[57] = AP_AXIMM_57_AWBURST;
            assign ap_AWLOCK[57] = AP_AXIMM_57_AWLOCK;
            assign ap_AWCACHE[57] = AP_AXIMM_57_AWCACHE;
            assign ap_AWPROT[57] = AP_AXIMM_57_AWPROT;
            assign ap_AWREGION[57] = AP_AXIMM_57_AWREGION;
            assign ap_AWQOS[57] = AP_AXIMM_57_AWQOS;
            assign ap_AWVALID[57] = AP_AXIMM_57_AWVALID;
            assign AP_AXIMM_57_AWREADY = ap_AWREADY[57];
            assign ap_WDATA[57][M_AXIMM_57_DATA_WIDTH-1:0] = AP_AXIMM_57_WDATA;
            assign ap_WSTRB[57][M_AXIMM_57_DATA_WIDTH/8-1:0] = AP_AXIMM_57_WSTRB;
            assign ap_WLAST[57] = AP_AXIMM_57_WLAST;
            assign ap_WVALID[57] = AP_AXIMM_57_WVALID;
            assign AP_AXIMM_57_WREADY = ap_WREADY[57];
            assign AP_AXIMM_57_BRESP = ap_BRESP[57];
            assign AP_AXIMM_57_BVALID = ap_BVALID[57];
            assign ap_BREADY[57] = AP_AXIMM_57_BREADY;
            assign ap_ARADDR[57][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_57_ARADDR;
            assign ap_ARLEN[57] = AP_AXIMM_57_ARLEN;
            assign ap_ARSIZE[57] = AP_AXIMM_57_ARSIZE;
            assign ap_ARBURST[57] = AP_AXIMM_57_ARBURST;
            assign ap_ARLOCK[57] = AP_AXIMM_57_ARLOCK;
            assign ap_ARCACHE[57] = AP_AXIMM_57_ARCACHE;
            assign ap_ARPROT[57] = AP_AXIMM_57_ARPROT;
            assign ap_ARREGION[57] = AP_AXIMM_57_ARREGION;
            assign ap_ARQOS[57] = AP_AXIMM_57_ARQOS;
            assign ap_ARVALID[57] = AP_AXIMM_57_ARVALID;
            assign AP_AXIMM_57_ARREADY = ap_ARREADY[57];
            assign AP_AXIMM_57_RDATA = ap_RDATA[57][M_AXIMM_57_DATA_WIDTH-1:0];
            assign AP_AXIMM_57_RRESP = ap_RRESP[57];
            assign AP_AXIMM_57_RLAST = ap_RLAST[57];
            assign AP_AXIMM_57_RVALID = ap_RVALID[57];
            assign ap_RREADY[57] = AP_AXIMM_57_RREADY;
            assign M_AXIMM_57_AWADDR = dm_AWADDR[57][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_57_AWLEN = dm_AWLEN[57];
            assign M_AXIMM_57_AWSIZE = dm_AWSIZE[57];
            assign M_AXIMM_57_AWBURST = dm_AWBURST[57];
            assign M_AXIMM_57_AWLOCK = dm_AWLOCK[57];
            assign M_AXIMM_57_AWCACHE = dm_AWCACHE[57];
            assign M_AXIMM_57_AWPROT = dm_AWPROT[57];
            assign M_AXIMM_57_AWREGION = dm_AWREGION[57];
            assign M_AXIMM_57_AWQOS = dm_AWQOS[57];
            assign M_AXIMM_57_AWVALID = dm_AWVALID[57];
            assign dm_AWREADY[57] = M_AXIMM_57_AWREADY;
            assign M_AXIMM_57_WDATA = dm_WDATA[57][M_AXIMM_57_DATA_WIDTH-1:0];
            assign M_AXIMM_57_WSTRB = dm_WSTRB[57][M_AXIMM_57_DATA_WIDTH/8-1:0];
            assign M_AXIMM_57_WLAST = dm_WLAST[57];
            assign M_AXIMM_57_WVALID = dm_WVALID[57];
            assign dm_WREADY[57] = M_AXIMM_57_WREADY;
            assign dm_BRESP[57] = M_AXIMM_57_BRESP;
            assign dm_BVALID[57] = M_AXIMM_57_BVALID;
            assign M_AXIMM_57_BREADY = dm_BREADY[57];
            assign M_AXIMM_57_ARADDR = dm_ARADDR[57][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_57_ARLEN = dm_ARLEN[57];
            assign M_AXIMM_57_ARSIZE = dm_ARSIZE[57];
            assign M_AXIMM_57_ARBURST = dm_ARBURST[57];
            assign M_AXIMM_57_ARLOCK = dm_ARLOCK[57];
            assign M_AXIMM_57_ARCACHE = dm_ARCACHE[57];
            assign M_AXIMM_57_ARPROT = dm_ARPROT[57];
            assign M_AXIMM_57_ARREGION = dm_ARREGION[57];
            assign M_AXIMM_57_ARQOS = dm_ARQOS[57];
            assign M_AXIMM_57_ARVALID = dm_ARVALID[57];
            assign dm_ARREADY[57] = M_AXIMM_57_ARREADY;
            assign dm_RDATA[57][M_AXIMM_57_DATA_WIDTH-1:0] = M_AXIMM_57_RDATA;
            assign dm_RRESP[57] = M_AXIMM_57_RRESP;
            assign dm_RLAST[57] = M_AXIMM_57_RLAST;
            assign dm_RVALID[57] = M_AXIMM_57_RVALID;
            assign M_AXIMM_57_RREADY = dm_RREADY[57];
        end
        if(C_NUM_AXIMMs > 58) begin
            assign ap_AWADDR[58][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_58_AWADDR;
            assign ap_AWLEN[58] = AP_AXIMM_58_AWLEN;
            assign ap_AWSIZE[58] = AP_AXIMM_58_AWSIZE;
            assign ap_AWBURST[58] = AP_AXIMM_58_AWBURST;
            assign ap_AWLOCK[58] = AP_AXIMM_58_AWLOCK;
            assign ap_AWCACHE[58] = AP_AXIMM_58_AWCACHE;
            assign ap_AWPROT[58] = AP_AXIMM_58_AWPROT;
            assign ap_AWREGION[58] = AP_AXIMM_58_AWREGION;
            assign ap_AWQOS[58] = AP_AXIMM_58_AWQOS;
            assign ap_AWVALID[58] = AP_AXIMM_58_AWVALID;
            assign AP_AXIMM_58_AWREADY = ap_AWREADY[58];
            assign ap_WDATA[58][M_AXIMM_58_DATA_WIDTH-1:0] = AP_AXIMM_58_WDATA;
            assign ap_WSTRB[58][M_AXIMM_58_DATA_WIDTH/8-1:0] = AP_AXIMM_58_WSTRB;
            assign ap_WLAST[58] = AP_AXIMM_58_WLAST;
            assign ap_WVALID[58] = AP_AXIMM_58_WVALID;
            assign AP_AXIMM_58_WREADY = ap_WREADY[58];
            assign AP_AXIMM_58_BRESP = ap_BRESP[58];
            assign AP_AXIMM_58_BVALID = ap_BVALID[58];
            assign ap_BREADY[58] = AP_AXIMM_58_BREADY;
            assign ap_ARADDR[58][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_58_ARADDR;
            assign ap_ARLEN[58] = AP_AXIMM_58_ARLEN;
            assign ap_ARSIZE[58] = AP_AXIMM_58_ARSIZE;
            assign ap_ARBURST[58] = AP_AXIMM_58_ARBURST;
            assign ap_ARLOCK[58] = AP_AXIMM_58_ARLOCK;
            assign ap_ARCACHE[58] = AP_AXIMM_58_ARCACHE;
            assign ap_ARPROT[58] = AP_AXIMM_58_ARPROT;
            assign ap_ARREGION[58] = AP_AXIMM_58_ARREGION;
            assign ap_ARQOS[58] = AP_AXIMM_58_ARQOS;
            assign ap_ARVALID[58] = AP_AXIMM_58_ARVALID;
            assign AP_AXIMM_58_ARREADY = ap_ARREADY[58];
            assign AP_AXIMM_58_RDATA = ap_RDATA[58][M_AXIMM_58_DATA_WIDTH-1:0];
            assign AP_AXIMM_58_RRESP = ap_RRESP[58];
            assign AP_AXIMM_58_RLAST = ap_RLAST[58];
            assign AP_AXIMM_58_RVALID = ap_RVALID[58];
            assign ap_RREADY[58] = AP_AXIMM_58_RREADY;
            assign M_AXIMM_58_AWADDR = dm_AWADDR[58][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_58_AWLEN = dm_AWLEN[58];
            assign M_AXIMM_58_AWSIZE = dm_AWSIZE[58];
            assign M_AXIMM_58_AWBURST = dm_AWBURST[58];
            assign M_AXIMM_58_AWLOCK = dm_AWLOCK[58];
            assign M_AXIMM_58_AWCACHE = dm_AWCACHE[58];
            assign M_AXIMM_58_AWPROT = dm_AWPROT[58];
            assign M_AXIMM_58_AWREGION = dm_AWREGION[58];
            assign M_AXIMM_58_AWQOS = dm_AWQOS[58];
            assign M_AXIMM_58_AWVALID = dm_AWVALID[58];
            assign dm_AWREADY[58] = M_AXIMM_58_AWREADY;
            assign M_AXIMM_58_WDATA = dm_WDATA[58][M_AXIMM_58_DATA_WIDTH-1:0];
            assign M_AXIMM_58_WSTRB = dm_WSTRB[58][M_AXIMM_58_DATA_WIDTH/8-1:0];
            assign M_AXIMM_58_WLAST = dm_WLAST[58];
            assign M_AXIMM_58_WVALID = dm_WVALID[58];
            assign dm_WREADY[58] = M_AXIMM_58_WREADY;
            assign dm_BRESP[58] = M_AXIMM_58_BRESP;
            assign dm_BVALID[58] = M_AXIMM_58_BVALID;
            assign M_AXIMM_58_BREADY = dm_BREADY[58];
            assign M_AXIMM_58_ARADDR = dm_ARADDR[58][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_58_ARLEN = dm_ARLEN[58];
            assign M_AXIMM_58_ARSIZE = dm_ARSIZE[58];
            assign M_AXIMM_58_ARBURST = dm_ARBURST[58];
            assign M_AXIMM_58_ARLOCK = dm_ARLOCK[58];
            assign M_AXIMM_58_ARCACHE = dm_ARCACHE[58];
            assign M_AXIMM_58_ARPROT = dm_ARPROT[58];
            assign M_AXIMM_58_ARREGION = dm_ARREGION[58];
            assign M_AXIMM_58_ARQOS = dm_ARQOS[58];
            assign M_AXIMM_58_ARVALID = dm_ARVALID[58];
            assign dm_ARREADY[58] = M_AXIMM_58_ARREADY;
            assign dm_RDATA[58][M_AXIMM_58_DATA_WIDTH-1:0] = M_AXIMM_58_RDATA;
            assign dm_RRESP[58] = M_AXIMM_58_RRESP;
            assign dm_RLAST[58] = M_AXIMM_58_RLAST;
            assign dm_RVALID[58] = M_AXIMM_58_RVALID;
            assign M_AXIMM_58_RREADY = dm_RREADY[58];
        end
        if(C_NUM_AXIMMs > 59) begin
            assign ap_AWADDR[59][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_59_AWADDR;
            assign ap_AWLEN[59] = AP_AXIMM_59_AWLEN;
            assign ap_AWSIZE[59] = AP_AXIMM_59_AWSIZE;
            assign ap_AWBURST[59] = AP_AXIMM_59_AWBURST;
            assign ap_AWLOCK[59] = AP_AXIMM_59_AWLOCK;
            assign ap_AWCACHE[59] = AP_AXIMM_59_AWCACHE;
            assign ap_AWPROT[59] = AP_AXIMM_59_AWPROT;
            assign ap_AWREGION[59] = AP_AXIMM_59_AWREGION;
            assign ap_AWQOS[59] = AP_AXIMM_59_AWQOS;
            assign ap_AWVALID[59] = AP_AXIMM_59_AWVALID;
            assign AP_AXIMM_59_AWREADY = ap_AWREADY[59];
            assign ap_WDATA[59][M_AXIMM_59_DATA_WIDTH-1:0] = AP_AXIMM_59_WDATA;
            assign ap_WSTRB[59][M_AXIMM_59_DATA_WIDTH/8-1:0] = AP_AXIMM_59_WSTRB;
            assign ap_WLAST[59] = AP_AXIMM_59_WLAST;
            assign ap_WVALID[59] = AP_AXIMM_59_WVALID;
            assign AP_AXIMM_59_WREADY = ap_WREADY[59];
            assign AP_AXIMM_59_BRESP = ap_BRESP[59];
            assign AP_AXIMM_59_BVALID = ap_BVALID[59];
            assign ap_BREADY[59] = AP_AXIMM_59_BREADY;
            assign ap_ARADDR[59][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_59_ARADDR;
            assign ap_ARLEN[59] = AP_AXIMM_59_ARLEN;
            assign ap_ARSIZE[59] = AP_AXIMM_59_ARSIZE;
            assign ap_ARBURST[59] = AP_AXIMM_59_ARBURST;
            assign ap_ARLOCK[59] = AP_AXIMM_59_ARLOCK;
            assign ap_ARCACHE[59] = AP_AXIMM_59_ARCACHE;
            assign ap_ARPROT[59] = AP_AXIMM_59_ARPROT;
            assign ap_ARREGION[59] = AP_AXIMM_59_ARREGION;
            assign ap_ARQOS[59] = AP_AXIMM_59_ARQOS;
            assign ap_ARVALID[59] = AP_AXIMM_59_ARVALID;
            assign AP_AXIMM_59_ARREADY = ap_ARREADY[59];
            assign AP_AXIMM_59_RDATA = ap_RDATA[59][M_AXIMM_59_DATA_WIDTH-1:0];
            assign AP_AXIMM_59_RRESP = ap_RRESP[59];
            assign AP_AXIMM_59_RLAST = ap_RLAST[59];
            assign AP_AXIMM_59_RVALID = ap_RVALID[59];
            assign ap_RREADY[59] = AP_AXIMM_59_RREADY;
            assign M_AXIMM_59_AWADDR = dm_AWADDR[59][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_59_AWLEN = dm_AWLEN[59];
            assign M_AXIMM_59_AWSIZE = dm_AWSIZE[59];
            assign M_AXIMM_59_AWBURST = dm_AWBURST[59];
            assign M_AXIMM_59_AWLOCK = dm_AWLOCK[59];
            assign M_AXIMM_59_AWCACHE = dm_AWCACHE[59];
            assign M_AXIMM_59_AWPROT = dm_AWPROT[59];
            assign M_AXIMM_59_AWREGION = dm_AWREGION[59];
            assign M_AXIMM_59_AWQOS = dm_AWQOS[59];
            assign M_AXIMM_59_AWVALID = dm_AWVALID[59];
            assign dm_AWREADY[59] = M_AXIMM_59_AWREADY;
            assign M_AXIMM_59_WDATA = dm_WDATA[59][M_AXIMM_59_DATA_WIDTH-1:0];
            assign M_AXIMM_59_WSTRB = dm_WSTRB[59][M_AXIMM_59_DATA_WIDTH/8-1:0];
            assign M_AXIMM_59_WLAST = dm_WLAST[59];
            assign M_AXIMM_59_WVALID = dm_WVALID[59];
            assign dm_WREADY[59] = M_AXIMM_59_WREADY;
            assign dm_BRESP[59] = M_AXIMM_59_BRESP;
            assign dm_BVALID[59] = M_AXIMM_59_BVALID;
            assign M_AXIMM_59_BREADY = dm_BREADY[59];
            assign M_AXIMM_59_ARADDR = dm_ARADDR[59][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_59_ARLEN = dm_ARLEN[59];
            assign M_AXIMM_59_ARSIZE = dm_ARSIZE[59];
            assign M_AXIMM_59_ARBURST = dm_ARBURST[59];
            assign M_AXIMM_59_ARLOCK = dm_ARLOCK[59];
            assign M_AXIMM_59_ARCACHE = dm_ARCACHE[59];
            assign M_AXIMM_59_ARPROT = dm_ARPROT[59];
            assign M_AXIMM_59_ARREGION = dm_ARREGION[59];
            assign M_AXIMM_59_ARQOS = dm_ARQOS[59];
            assign M_AXIMM_59_ARVALID = dm_ARVALID[59];
            assign dm_ARREADY[59] = M_AXIMM_59_ARREADY;
            assign dm_RDATA[59][M_AXIMM_59_DATA_WIDTH-1:0] = M_AXIMM_59_RDATA;
            assign dm_RRESP[59] = M_AXIMM_59_RRESP;
            assign dm_RLAST[59] = M_AXIMM_59_RLAST;
            assign dm_RVALID[59] = M_AXIMM_59_RVALID;
            assign M_AXIMM_59_RREADY = dm_RREADY[59];
        end
        if(C_NUM_AXIMMs > 60) begin
            assign ap_AWADDR[60][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_60_AWADDR;
            assign ap_AWLEN[60] = AP_AXIMM_60_AWLEN;
            assign ap_AWSIZE[60] = AP_AXIMM_60_AWSIZE;
            assign ap_AWBURST[60] = AP_AXIMM_60_AWBURST;
            assign ap_AWLOCK[60] = AP_AXIMM_60_AWLOCK;
            assign ap_AWCACHE[60] = AP_AXIMM_60_AWCACHE;
            assign ap_AWPROT[60] = AP_AXIMM_60_AWPROT;
            assign ap_AWREGION[60] = AP_AXIMM_60_AWREGION;
            assign ap_AWQOS[60] = AP_AXIMM_60_AWQOS;
            assign ap_AWVALID[60] = AP_AXIMM_60_AWVALID;
            assign AP_AXIMM_60_AWREADY = ap_AWREADY[60];
            assign ap_WDATA[60][M_AXIMM_60_DATA_WIDTH-1:0] = AP_AXIMM_60_WDATA;
            assign ap_WSTRB[60][M_AXIMM_60_DATA_WIDTH/8-1:0] = AP_AXIMM_60_WSTRB;
            assign ap_WLAST[60] = AP_AXIMM_60_WLAST;
            assign ap_WVALID[60] = AP_AXIMM_60_WVALID;
            assign AP_AXIMM_60_WREADY = ap_WREADY[60];
            assign AP_AXIMM_60_BRESP = ap_BRESP[60];
            assign AP_AXIMM_60_BVALID = ap_BVALID[60];
            assign ap_BREADY[60] = AP_AXIMM_60_BREADY;
            assign ap_ARADDR[60][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_60_ARADDR;
            assign ap_ARLEN[60] = AP_AXIMM_60_ARLEN;
            assign ap_ARSIZE[60] = AP_AXIMM_60_ARSIZE;
            assign ap_ARBURST[60] = AP_AXIMM_60_ARBURST;
            assign ap_ARLOCK[60] = AP_AXIMM_60_ARLOCK;
            assign ap_ARCACHE[60] = AP_AXIMM_60_ARCACHE;
            assign ap_ARPROT[60] = AP_AXIMM_60_ARPROT;
            assign ap_ARREGION[60] = AP_AXIMM_60_ARREGION;
            assign ap_ARQOS[60] = AP_AXIMM_60_ARQOS;
            assign ap_ARVALID[60] = AP_AXIMM_60_ARVALID;
            assign AP_AXIMM_60_ARREADY = ap_ARREADY[60];
            assign AP_AXIMM_60_RDATA = ap_RDATA[60][M_AXIMM_60_DATA_WIDTH-1:0];
            assign AP_AXIMM_60_RRESP = ap_RRESP[60];
            assign AP_AXIMM_60_RLAST = ap_RLAST[60];
            assign AP_AXIMM_60_RVALID = ap_RVALID[60];
            assign ap_RREADY[60] = AP_AXIMM_60_RREADY;
            assign M_AXIMM_60_AWADDR = dm_AWADDR[60][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_60_AWLEN = dm_AWLEN[60];
            assign M_AXIMM_60_AWSIZE = dm_AWSIZE[60];
            assign M_AXIMM_60_AWBURST = dm_AWBURST[60];
            assign M_AXIMM_60_AWLOCK = dm_AWLOCK[60];
            assign M_AXIMM_60_AWCACHE = dm_AWCACHE[60];
            assign M_AXIMM_60_AWPROT = dm_AWPROT[60];
            assign M_AXIMM_60_AWREGION = dm_AWREGION[60];
            assign M_AXIMM_60_AWQOS = dm_AWQOS[60];
            assign M_AXIMM_60_AWVALID = dm_AWVALID[60];
            assign dm_AWREADY[60] = M_AXIMM_60_AWREADY;
            assign M_AXIMM_60_WDATA = dm_WDATA[60][M_AXIMM_60_DATA_WIDTH-1:0];
            assign M_AXIMM_60_WSTRB = dm_WSTRB[60][M_AXIMM_60_DATA_WIDTH/8-1:0];
            assign M_AXIMM_60_WLAST = dm_WLAST[60];
            assign M_AXIMM_60_WVALID = dm_WVALID[60];
            assign dm_WREADY[60] = M_AXIMM_60_WREADY;
            assign dm_BRESP[60] = M_AXIMM_60_BRESP;
            assign dm_BVALID[60] = M_AXIMM_60_BVALID;
            assign M_AXIMM_60_BREADY = dm_BREADY[60];
            assign M_AXIMM_60_ARADDR = dm_ARADDR[60][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_60_ARLEN = dm_ARLEN[60];
            assign M_AXIMM_60_ARSIZE = dm_ARSIZE[60];
            assign M_AXIMM_60_ARBURST = dm_ARBURST[60];
            assign M_AXIMM_60_ARLOCK = dm_ARLOCK[60];
            assign M_AXIMM_60_ARCACHE = dm_ARCACHE[60];
            assign M_AXIMM_60_ARPROT = dm_ARPROT[60];
            assign M_AXIMM_60_ARREGION = dm_ARREGION[60];
            assign M_AXIMM_60_ARQOS = dm_ARQOS[60];
            assign M_AXIMM_60_ARVALID = dm_ARVALID[60];
            assign dm_ARREADY[60] = M_AXIMM_60_ARREADY;
            assign dm_RDATA[60][M_AXIMM_60_DATA_WIDTH-1:0] = M_AXIMM_60_RDATA;
            assign dm_RRESP[60] = M_AXIMM_60_RRESP;
            assign dm_RLAST[60] = M_AXIMM_60_RLAST;
            assign dm_RVALID[60] = M_AXIMM_60_RVALID;
            assign M_AXIMM_60_RREADY = dm_RREADY[60];
        end
        if(C_NUM_AXIMMs > 61) begin
            assign ap_AWADDR[61][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_61_AWADDR;
            assign ap_AWLEN[61] = AP_AXIMM_61_AWLEN;
            assign ap_AWSIZE[61] = AP_AXIMM_61_AWSIZE;
            assign ap_AWBURST[61] = AP_AXIMM_61_AWBURST;
            assign ap_AWLOCK[61] = AP_AXIMM_61_AWLOCK;
            assign ap_AWCACHE[61] = AP_AXIMM_61_AWCACHE;
            assign ap_AWPROT[61] = AP_AXIMM_61_AWPROT;
            assign ap_AWREGION[61] = AP_AXIMM_61_AWREGION;
            assign ap_AWQOS[61] = AP_AXIMM_61_AWQOS;
            assign ap_AWVALID[61] = AP_AXIMM_61_AWVALID;
            assign AP_AXIMM_61_AWREADY = ap_AWREADY[61];
            assign ap_WDATA[61][M_AXIMM_61_DATA_WIDTH-1:0] = AP_AXIMM_61_WDATA;
            assign ap_WSTRB[61][M_AXIMM_61_DATA_WIDTH/8-1:0] = AP_AXIMM_61_WSTRB;
            assign ap_WLAST[61] = AP_AXIMM_61_WLAST;
            assign ap_WVALID[61] = AP_AXIMM_61_WVALID;
            assign AP_AXIMM_61_WREADY = ap_WREADY[61];
            assign AP_AXIMM_61_BRESP = ap_BRESP[61];
            assign AP_AXIMM_61_BVALID = ap_BVALID[61];
            assign ap_BREADY[61] = AP_AXIMM_61_BREADY;
            assign ap_ARADDR[61][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_61_ARADDR;
            assign ap_ARLEN[61] = AP_AXIMM_61_ARLEN;
            assign ap_ARSIZE[61] = AP_AXIMM_61_ARSIZE;
            assign ap_ARBURST[61] = AP_AXIMM_61_ARBURST;
            assign ap_ARLOCK[61] = AP_AXIMM_61_ARLOCK;
            assign ap_ARCACHE[61] = AP_AXIMM_61_ARCACHE;
            assign ap_ARPROT[61] = AP_AXIMM_61_ARPROT;
            assign ap_ARREGION[61] = AP_AXIMM_61_ARREGION;
            assign ap_ARQOS[61] = AP_AXIMM_61_ARQOS;
            assign ap_ARVALID[61] = AP_AXIMM_61_ARVALID;
            assign AP_AXIMM_61_ARREADY = ap_ARREADY[61];
            assign AP_AXIMM_61_RDATA = ap_RDATA[61][M_AXIMM_61_DATA_WIDTH-1:0];
            assign AP_AXIMM_61_RRESP = ap_RRESP[61];
            assign AP_AXIMM_61_RLAST = ap_RLAST[61];
            assign AP_AXIMM_61_RVALID = ap_RVALID[61];
            assign ap_RREADY[61] = AP_AXIMM_61_RREADY;
            assign M_AXIMM_61_AWADDR = dm_AWADDR[61][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_61_AWLEN = dm_AWLEN[61];
            assign M_AXIMM_61_AWSIZE = dm_AWSIZE[61];
            assign M_AXIMM_61_AWBURST = dm_AWBURST[61];
            assign M_AXIMM_61_AWLOCK = dm_AWLOCK[61];
            assign M_AXIMM_61_AWCACHE = dm_AWCACHE[61];
            assign M_AXIMM_61_AWPROT = dm_AWPROT[61];
            assign M_AXIMM_61_AWREGION = dm_AWREGION[61];
            assign M_AXIMM_61_AWQOS = dm_AWQOS[61];
            assign M_AXIMM_61_AWVALID = dm_AWVALID[61];
            assign dm_AWREADY[61] = M_AXIMM_61_AWREADY;
            assign M_AXIMM_61_WDATA = dm_WDATA[61][M_AXIMM_61_DATA_WIDTH-1:0];
            assign M_AXIMM_61_WSTRB = dm_WSTRB[61][M_AXIMM_61_DATA_WIDTH/8-1:0];
            assign M_AXIMM_61_WLAST = dm_WLAST[61];
            assign M_AXIMM_61_WVALID = dm_WVALID[61];
            assign dm_WREADY[61] = M_AXIMM_61_WREADY;
            assign dm_BRESP[61] = M_AXIMM_61_BRESP;
            assign dm_BVALID[61] = M_AXIMM_61_BVALID;
            assign M_AXIMM_61_BREADY = dm_BREADY[61];
            assign M_AXIMM_61_ARADDR = dm_ARADDR[61][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_61_ARLEN = dm_ARLEN[61];
            assign M_AXIMM_61_ARSIZE = dm_ARSIZE[61];
            assign M_AXIMM_61_ARBURST = dm_ARBURST[61];
            assign M_AXIMM_61_ARLOCK = dm_ARLOCK[61];
            assign M_AXIMM_61_ARCACHE = dm_ARCACHE[61];
            assign M_AXIMM_61_ARPROT = dm_ARPROT[61];
            assign M_AXIMM_61_ARREGION = dm_ARREGION[61];
            assign M_AXIMM_61_ARQOS = dm_ARQOS[61];
            assign M_AXIMM_61_ARVALID = dm_ARVALID[61];
            assign dm_ARREADY[61] = M_AXIMM_61_ARREADY;
            assign dm_RDATA[61][M_AXIMM_61_DATA_WIDTH-1:0] = M_AXIMM_61_RDATA;
            assign dm_RRESP[61] = M_AXIMM_61_RRESP;
            assign dm_RLAST[61] = M_AXIMM_61_RLAST;
            assign dm_RVALID[61] = M_AXIMM_61_RVALID;
            assign M_AXIMM_61_RREADY = dm_RREADY[61];
        end
        if(C_NUM_AXIMMs > 62) begin
            assign ap_AWADDR[62][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_62_AWADDR;
            assign ap_AWLEN[62] = AP_AXIMM_62_AWLEN;
            assign ap_AWSIZE[62] = AP_AXIMM_62_AWSIZE;
            assign ap_AWBURST[62] = AP_AXIMM_62_AWBURST;
            assign ap_AWLOCK[62] = AP_AXIMM_62_AWLOCK;
            assign ap_AWCACHE[62] = AP_AXIMM_62_AWCACHE;
            assign ap_AWPROT[62] = AP_AXIMM_62_AWPROT;
            assign ap_AWREGION[62] = AP_AXIMM_62_AWREGION;
            assign ap_AWQOS[62] = AP_AXIMM_62_AWQOS;
            assign ap_AWVALID[62] = AP_AXIMM_62_AWVALID;
            assign AP_AXIMM_62_AWREADY = ap_AWREADY[62];
            assign ap_WDATA[62][M_AXIMM_62_DATA_WIDTH-1:0] = AP_AXIMM_62_WDATA;
            assign ap_WSTRB[62][M_AXIMM_62_DATA_WIDTH/8-1:0] = AP_AXIMM_62_WSTRB;
            assign ap_WLAST[62] = AP_AXIMM_62_WLAST;
            assign ap_WVALID[62] = AP_AXIMM_62_WVALID;
            assign AP_AXIMM_62_WREADY = ap_WREADY[62];
            assign AP_AXIMM_62_BRESP = ap_BRESP[62];
            assign AP_AXIMM_62_BVALID = ap_BVALID[62];
            assign ap_BREADY[62] = AP_AXIMM_62_BREADY;
            assign ap_ARADDR[62][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_62_ARADDR;
            assign ap_ARLEN[62] = AP_AXIMM_62_ARLEN;
            assign ap_ARSIZE[62] = AP_AXIMM_62_ARSIZE;
            assign ap_ARBURST[62] = AP_AXIMM_62_ARBURST;
            assign ap_ARLOCK[62] = AP_AXIMM_62_ARLOCK;
            assign ap_ARCACHE[62] = AP_AXIMM_62_ARCACHE;
            assign ap_ARPROT[62] = AP_AXIMM_62_ARPROT;
            assign ap_ARREGION[62] = AP_AXIMM_62_ARREGION;
            assign ap_ARQOS[62] = AP_AXIMM_62_ARQOS;
            assign ap_ARVALID[62] = AP_AXIMM_62_ARVALID;
            assign AP_AXIMM_62_ARREADY = ap_ARREADY[62];
            assign AP_AXIMM_62_RDATA = ap_RDATA[62][M_AXIMM_62_DATA_WIDTH-1:0];
            assign AP_AXIMM_62_RRESP = ap_RRESP[62];
            assign AP_AXIMM_62_RLAST = ap_RLAST[62];
            assign AP_AXIMM_62_RVALID = ap_RVALID[62];
            assign ap_RREADY[62] = AP_AXIMM_62_RREADY;
            assign M_AXIMM_62_AWADDR = dm_AWADDR[62][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_62_AWLEN = dm_AWLEN[62];
            assign M_AXIMM_62_AWSIZE = dm_AWSIZE[62];
            assign M_AXIMM_62_AWBURST = dm_AWBURST[62];
            assign M_AXIMM_62_AWLOCK = dm_AWLOCK[62];
            assign M_AXIMM_62_AWCACHE = dm_AWCACHE[62];
            assign M_AXIMM_62_AWPROT = dm_AWPROT[62];
            assign M_AXIMM_62_AWREGION = dm_AWREGION[62];
            assign M_AXIMM_62_AWQOS = dm_AWQOS[62];
            assign M_AXIMM_62_AWVALID = dm_AWVALID[62];
            assign dm_AWREADY[62] = M_AXIMM_62_AWREADY;
            assign M_AXIMM_62_WDATA = dm_WDATA[62][M_AXIMM_62_DATA_WIDTH-1:0];
            assign M_AXIMM_62_WSTRB = dm_WSTRB[62][M_AXIMM_62_DATA_WIDTH/8-1:0];
            assign M_AXIMM_62_WLAST = dm_WLAST[62];
            assign M_AXIMM_62_WVALID = dm_WVALID[62];
            assign dm_WREADY[62] = M_AXIMM_62_WREADY;
            assign dm_BRESP[62] = M_AXIMM_62_BRESP;
            assign dm_BVALID[62] = M_AXIMM_62_BVALID;
            assign M_AXIMM_62_BREADY = dm_BREADY[62];
            assign M_AXIMM_62_ARADDR = dm_ARADDR[62][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_62_ARLEN = dm_ARLEN[62];
            assign M_AXIMM_62_ARSIZE = dm_ARSIZE[62];
            assign M_AXIMM_62_ARBURST = dm_ARBURST[62];
            assign M_AXIMM_62_ARLOCK = dm_ARLOCK[62];
            assign M_AXIMM_62_ARCACHE = dm_ARCACHE[62];
            assign M_AXIMM_62_ARPROT = dm_ARPROT[62];
            assign M_AXIMM_62_ARREGION = dm_ARREGION[62];
            assign M_AXIMM_62_ARQOS = dm_ARQOS[62];
            assign M_AXIMM_62_ARVALID = dm_ARVALID[62];
            assign dm_ARREADY[62] = M_AXIMM_62_ARREADY;
            assign dm_RDATA[62][M_AXIMM_62_DATA_WIDTH-1:0] = M_AXIMM_62_RDATA;
            assign dm_RRESP[62] = M_AXIMM_62_RRESP;
            assign dm_RLAST[62] = M_AXIMM_62_RLAST;
            assign dm_RVALID[62] = M_AXIMM_62_RVALID;
            assign M_AXIMM_62_RREADY = dm_RREADY[62];
        end
        if(C_NUM_AXIMMs > 63) begin
            assign ap_AWADDR[63][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_63_AWADDR;
            assign ap_AWLEN[63] = AP_AXIMM_63_AWLEN;
            assign ap_AWSIZE[63] = AP_AXIMM_63_AWSIZE;
            assign ap_AWBURST[63] = AP_AXIMM_63_AWBURST;
            assign ap_AWLOCK[63] = AP_AXIMM_63_AWLOCK;
            assign ap_AWCACHE[63] = AP_AXIMM_63_AWCACHE;
            assign ap_AWPROT[63] = AP_AXIMM_63_AWPROT;
            assign ap_AWREGION[63] = AP_AXIMM_63_AWREGION;
            assign ap_AWQOS[63] = AP_AXIMM_63_AWQOS;
            assign ap_AWVALID[63] = AP_AXIMM_63_AWVALID;
            assign AP_AXIMM_63_AWREADY = ap_AWREADY[63];
            assign ap_WDATA[63][M_AXIMM_63_DATA_WIDTH-1:0] = AP_AXIMM_63_WDATA;
            assign ap_WSTRB[63][M_AXIMM_63_DATA_WIDTH/8-1:0] = AP_AXIMM_63_WSTRB;
            assign ap_WLAST[63] = AP_AXIMM_63_WLAST;
            assign ap_WVALID[63] = AP_AXIMM_63_WVALID;
            assign AP_AXIMM_63_WREADY = ap_WREADY[63];
            assign AP_AXIMM_63_BRESP = ap_BRESP[63];
            assign AP_AXIMM_63_BVALID = ap_BVALID[63];
            assign ap_BREADY[63] = AP_AXIMM_63_BREADY;
            assign ap_ARADDR[63][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_63_ARADDR;
            assign ap_ARLEN[63] = AP_AXIMM_63_ARLEN;
            assign ap_ARSIZE[63] = AP_AXIMM_63_ARSIZE;
            assign ap_ARBURST[63] = AP_AXIMM_63_ARBURST;
            assign ap_ARLOCK[63] = AP_AXIMM_63_ARLOCK;
            assign ap_ARCACHE[63] = AP_AXIMM_63_ARCACHE;
            assign ap_ARPROT[63] = AP_AXIMM_63_ARPROT;
            assign ap_ARREGION[63] = AP_AXIMM_63_ARREGION;
            assign ap_ARQOS[63] = AP_AXIMM_63_ARQOS;
            assign ap_ARVALID[63] = AP_AXIMM_63_ARVALID;
            assign AP_AXIMM_63_ARREADY = ap_ARREADY[63];
            assign AP_AXIMM_63_RDATA = ap_RDATA[63][M_AXIMM_63_DATA_WIDTH-1:0];
            assign AP_AXIMM_63_RRESP = ap_RRESP[63];
            assign AP_AXIMM_63_RLAST = ap_RLAST[63];
            assign AP_AXIMM_63_RVALID = ap_RVALID[63];
            assign ap_RREADY[63] = AP_AXIMM_63_RREADY;
            assign M_AXIMM_63_AWADDR = dm_AWADDR[63][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_63_AWLEN = dm_AWLEN[63];
            assign M_AXIMM_63_AWSIZE = dm_AWSIZE[63];
            assign M_AXIMM_63_AWBURST = dm_AWBURST[63];
            assign M_AXIMM_63_AWLOCK = dm_AWLOCK[63];
            assign M_AXIMM_63_AWCACHE = dm_AWCACHE[63];
            assign M_AXIMM_63_AWPROT = dm_AWPROT[63];
            assign M_AXIMM_63_AWREGION = dm_AWREGION[63];
            assign M_AXIMM_63_AWQOS = dm_AWQOS[63];
            assign M_AXIMM_63_AWVALID = dm_AWVALID[63];
            assign dm_AWREADY[63] = M_AXIMM_63_AWREADY;
            assign M_AXIMM_63_WDATA = dm_WDATA[63][M_AXIMM_63_DATA_WIDTH-1:0];
            assign M_AXIMM_63_WSTRB = dm_WSTRB[63][M_AXIMM_63_DATA_WIDTH/8-1:0];
            assign M_AXIMM_63_WLAST = dm_WLAST[63];
            assign M_AXIMM_63_WVALID = dm_WVALID[63];
            assign dm_WREADY[63] = M_AXIMM_63_WREADY;
            assign dm_BRESP[63] = M_AXIMM_63_BRESP;
            assign dm_BVALID[63] = M_AXIMM_63_BVALID;
            assign M_AXIMM_63_BREADY = dm_BREADY[63];
            assign M_AXIMM_63_ARADDR = dm_ARADDR[63][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_63_ARLEN = dm_ARLEN[63];
            assign M_AXIMM_63_ARSIZE = dm_ARSIZE[63];
            assign M_AXIMM_63_ARBURST = dm_ARBURST[63];
            assign M_AXIMM_63_ARLOCK = dm_ARLOCK[63];
            assign M_AXIMM_63_ARCACHE = dm_ARCACHE[63];
            assign M_AXIMM_63_ARPROT = dm_ARPROT[63];
            assign M_AXIMM_63_ARREGION = dm_ARREGION[63];
            assign M_AXIMM_63_ARQOS = dm_ARQOS[63];
            assign M_AXIMM_63_ARVALID = dm_ARVALID[63];
            assign dm_ARREADY[63] = M_AXIMM_63_ARREADY;
            assign dm_RDATA[63][M_AXIMM_63_DATA_WIDTH-1:0] = M_AXIMM_63_RDATA;
            assign dm_RRESP[63] = M_AXIMM_63_RRESP;
            assign dm_RLAST[63] = M_AXIMM_63_RLAST;
            assign dm_RVALID[63] = M_AXIMM_63_RVALID;
            assign M_AXIMM_63_RREADY = dm_RREADY[63];
        end
        if(C_NUM_AXIMMs > 64) begin
            assign ap_AWADDR[64][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_64_AWADDR;
            assign ap_AWLEN[64] = AP_AXIMM_64_AWLEN;
            assign ap_AWSIZE[64] = AP_AXIMM_64_AWSIZE;
            assign ap_AWBURST[64] = AP_AXIMM_64_AWBURST;
            assign ap_AWLOCK[64] = AP_AXIMM_64_AWLOCK;
            assign ap_AWCACHE[64] = AP_AXIMM_64_AWCACHE;
            assign ap_AWPROT[64] = AP_AXIMM_64_AWPROT;
            assign ap_AWREGION[64] = AP_AXIMM_64_AWREGION;
            assign ap_AWQOS[64] = AP_AXIMM_64_AWQOS;
            assign ap_AWVALID[64] = AP_AXIMM_64_AWVALID;
            assign AP_AXIMM_64_AWREADY = ap_AWREADY[64];
            assign ap_WDATA[64][M_AXIMM_64_DATA_WIDTH-1:0] = AP_AXIMM_64_WDATA;
            assign ap_WSTRB[64][M_AXIMM_64_DATA_WIDTH/8-1:0] = AP_AXIMM_64_WSTRB;
            assign ap_WLAST[64] = AP_AXIMM_64_WLAST;
            assign ap_WVALID[64] = AP_AXIMM_64_WVALID;
            assign AP_AXIMM_64_WREADY = ap_WREADY[64];
            assign AP_AXIMM_64_BRESP = ap_BRESP[64];
            assign AP_AXIMM_64_BVALID = ap_BVALID[64];
            assign ap_BREADY[64] = AP_AXIMM_64_BREADY;
            assign ap_ARADDR[64][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_64_ARADDR;
            assign ap_ARLEN[64] = AP_AXIMM_64_ARLEN;
            assign ap_ARSIZE[64] = AP_AXIMM_64_ARSIZE;
            assign ap_ARBURST[64] = AP_AXIMM_64_ARBURST;
            assign ap_ARLOCK[64] = AP_AXIMM_64_ARLOCK;
            assign ap_ARCACHE[64] = AP_AXIMM_64_ARCACHE;
            assign ap_ARPROT[64] = AP_AXIMM_64_ARPROT;
            assign ap_ARREGION[64] = AP_AXIMM_64_ARREGION;
            assign ap_ARQOS[64] = AP_AXIMM_64_ARQOS;
            assign ap_ARVALID[64] = AP_AXIMM_64_ARVALID;
            assign AP_AXIMM_64_ARREADY = ap_ARREADY[64];
            assign AP_AXIMM_64_RDATA = ap_RDATA[64][M_AXIMM_64_DATA_WIDTH-1:0];
            assign AP_AXIMM_64_RRESP = ap_RRESP[64];
            assign AP_AXIMM_64_RLAST = ap_RLAST[64];
            assign AP_AXIMM_64_RVALID = ap_RVALID[64];
            assign ap_RREADY[64] = AP_AXIMM_64_RREADY;
            assign M_AXIMM_64_AWADDR = dm_AWADDR[64][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_64_AWLEN = dm_AWLEN[64];
            assign M_AXIMM_64_AWSIZE = dm_AWSIZE[64];
            assign M_AXIMM_64_AWBURST = dm_AWBURST[64];
            assign M_AXIMM_64_AWLOCK = dm_AWLOCK[64];
            assign M_AXIMM_64_AWCACHE = dm_AWCACHE[64];
            assign M_AXIMM_64_AWPROT = dm_AWPROT[64];
            assign M_AXIMM_64_AWREGION = dm_AWREGION[64];
            assign M_AXIMM_64_AWQOS = dm_AWQOS[64];
            assign M_AXIMM_64_AWVALID = dm_AWVALID[64];
            assign dm_AWREADY[64] = M_AXIMM_64_AWREADY;
            assign M_AXIMM_64_WDATA = dm_WDATA[64][M_AXIMM_64_DATA_WIDTH-1:0];
            assign M_AXIMM_64_WSTRB = dm_WSTRB[64][M_AXIMM_64_DATA_WIDTH/8-1:0];
            assign M_AXIMM_64_WLAST = dm_WLAST[64];
            assign M_AXIMM_64_WVALID = dm_WVALID[64];
            assign dm_WREADY[64] = M_AXIMM_64_WREADY;
            assign dm_BRESP[64] = M_AXIMM_64_BRESP;
            assign dm_BVALID[64] = M_AXIMM_64_BVALID;
            assign M_AXIMM_64_BREADY = dm_BREADY[64];
            assign M_AXIMM_64_ARADDR = dm_ARADDR[64][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_64_ARLEN = dm_ARLEN[64];
            assign M_AXIMM_64_ARSIZE = dm_ARSIZE[64];
            assign M_AXIMM_64_ARBURST = dm_ARBURST[64];
            assign M_AXIMM_64_ARLOCK = dm_ARLOCK[64];
            assign M_AXIMM_64_ARCACHE = dm_ARCACHE[64];
            assign M_AXIMM_64_ARPROT = dm_ARPROT[64];
            assign M_AXIMM_64_ARREGION = dm_ARREGION[64];
            assign M_AXIMM_64_ARQOS = dm_ARQOS[64];
            assign M_AXIMM_64_ARVALID = dm_ARVALID[64];
            assign dm_ARREADY[64] = M_AXIMM_64_ARREADY;
            assign dm_RDATA[64][M_AXIMM_64_DATA_WIDTH-1:0] = M_AXIMM_64_RDATA;
            assign dm_RRESP[64] = M_AXIMM_64_RRESP;
            assign dm_RLAST[64] = M_AXIMM_64_RLAST;
            assign dm_RVALID[64] = M_AXIMM_64_RVALID;
            assign M_AXIMM_64_RREADY = dm_RREADY[64];
        end
        if(C_NUM_AXIMMs > 65) begin
            assign ap_AWADDR[65][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_65_AWADDR;
            assign ap_AWLEN[65] = AP_AXIMM_65_AWLEN;
            assign ap_AWSIZE[65] = AP_AXIMM_65_AWSIZE;
            assign ap_AWBURST[65] = AP_AXIMM_65_AWBURST;
            assign ap_AWLOCK[65] = AP_AXIMM_65_AWLOCK;
            assign ap_AWCACHE[65] = AP_AXIMM_65_AWCACHE;
            assign ap_AWPROT[65] = AP_AXIMM_65_AWPROT;
            assign ap_AWREGION[65] = AP_AXIMM_65_AWREGION;
            assign ap_AWQOS[65] = AP_AXIMM_65_AWQOS;
            assign ap_AWVALID[65] = AP_AXIMM_65_AWVALID;
            assign AP_AXIMM_65_AWREADY = ap_AWREADY[65];
            assign ap_WDATA[65][M_AXIMM_65_DATA_WIDTH-1:0] = AP_AXIMM_65_WDATA;
            assign ap_WSTRB[65][M_AXIMM_65_DATA_WIDTH/8-1:0] = AP_AXIMM_65_WSTRB;
            assign ap_WLAST[65] = AP_AXIMM_65_WLAST;
            assign ap_WVALID[65] = AP_AXIMM_65_WVALID;
            assign AP_AXIMM_65_WREADY = ap_WREADY[65];
            assign AP_AXIMM_65_BRESP = ap_BRESP[65];
            assign AP_AXIMM_65_BVALID = ap_BVALID[65];
            assign ap_BREADY[65] = AP_AXIMM_65_BREADY;
            assign ap_ARADDR[65][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_65_ARADDR;
            assign ap_ARLEN[65] = AP_AXIMM_65_ARLEN;
            assign ap_ARSIZE[65] = AP_AXIMM_65_ARSIZE;
            assign ap_ARBURST[65] = AP_AXIMM_65_ARBURST;
            assign ap_ARLOCK[65] = AP_AXIMM_65_ARLOCK;
            assign ap_ARCACHE[65] = AP_AXIMM_65_ARCACHE;
            assign ap_ARPROT[65] = AP_AXIMM_65_ARPROT;
            assign ap_ARREGION[65] = AP_AXIMM_65_ARREGION;
            assign ap_ARQOS[65] = AP_AXIMM_65_ARQOS;
            assign ap_ARVALID[65] = AP_AXIMM_65_ARVALID;
            assign AP_AXIMM_65_ARREADY = ap_ARREADY[65];
            assign AP_AXIMM_65_RDATA = ap_RDATA[65][M_AXIMM_65_DATA_WIDTH-1:0];
            assign AP_AXIMM_65_RRESP = ap_RRESP[65];
            assign AP_AXIMM_65_RLAST = ap_RLAST[65];
            assign AP_AXIMM_65_RVALID = ap_RVALID[65];
            assign ap_RREADY[65] = AP_AXIMM_65_RREADY;
            assign M_AXIMM_65_AWADDR = dm_AWADDR[65][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_65_AWLEN = dm_AWLEN[65];
            assign M_AXIMM_65_AWSIZE = dm_AWSIZE[65];
            assign M_AXIMM_65_AWBURST = dm_AWBURST[65];
            assign M_AXIMM_65_AWLOCK = dm_AWLOCK[65];
            assign M_AXIMM_65_AWCACHE = dm_AWCACHE[65];
            assign M_AXIMM_65_AWPROT = dm_AWPROT[65];
            assign M_AXIMM_65_AWREGION = dm_AWREGION[65];
            assign M_AXIMM_65_AWQOS = dm_AWQOS[65];
            assign M_AXIMM_65_AWVALID = dm_AWVALID[65];
            assign dm_AWREADY[65] = M_AXIMM_65_AWREADY;
            assign M_AXIMM_65_WDATA = dm_WDATA[65][M_AXIMM_65_DATA_WIDTH-1:0];
            assign M_AXIMM_65_WSTRB = dm_WSTRB[65][M_AXIMM_65_DATA_WIDTH/8-1:0];
            assign M_AXIMM_65_WLAST = dm_WLAST[65];
            assign M_AXIMM_65_WVALID = dm_WVALID[65];
            assign dm_WREADY[65] = M_AXIMM_65_WREADY;
            assign dm_BRESP[65] = M_AXIMM_65_BRESP;
            assign dm_BVALID[65] = M_AXIMM_65_BVALID;
            assign M_AXIMM_65_BREADY = dm_BREADY[65];
            assign M_AXIMM_65_ARADDR = dm_ARADDR[65][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_65_ARLEN = dm_ARLEN[65];
            assign M_AXIMM_65_ARSIZE = dm_ARSIZE[65];
            assign M_AXIMM_65_ARBURST = dm_ARBURST[65];
            assign M_AXIMM_65_ARLOCK = dm_ARLOCK[65];
            assign M_AXIMM_65_ARCACHE = dm_ARCACHE[65];
            assign M_AXIMM_65_ARPROT = dm_ARPROT[65];
            assign M_AXIMM_65_ARREGION = dm_ARREGION[65];
            assign M_AXIMM_65_ARQOS = dm_ARQOS[65];
            assign M_AXIMM_65_ARVALID = dm_ARVALID[65];
            assign dm_ARREADY[65] = M_AXIMM_65_ARREADY;
            assign dm_RDATA[65][M_AXIMM_65_DATA_WIDTH-1:0] = M_AXIMM_65_RDATA;
            assign dm_RRESP[65] = M_AXIMM_65_RRESP;
            assign dm_RLAST[65] = M_AXIMM_65_RLAST;
            assign dm_RVALID[65] = M_AXIMM_65_RVALID;
            assign M_AXIMM_65_RREADY = dm_RREADY[65];
        end
        if(C_NUM_AXIMMs > 66) begin
            assign ap_AWADDR[66][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_66_AWADDR;
            assign ap_AWLEN[66] = AP_AXIMM_66_AWLEN;
            assign ap_AWSIZE[66] = AP_AXIMM_66_AWSIZE;
            assign ap_AWBURST[66] = AP_AXIMM_66_AWBURST;
            assign ap_AWLOCK[66] = AP_AXIMM_66_AWLOCK;
            assign ap_AWCACHE[66] = AP_AXIMM_66_AWCACHE;
            assign ap_AWPROT[66] = AP_AXIMM_66_AWPROT;
            assign ap_AWREGION[66] = AP_AXIMM_66_AWREGION;
            assign ap_AWQOS[66] = AP_AXIMM_66_AWQOS;
            assign ap_AWVALID[66] = AP_AXIMM_66_AWVALID;
            assign AP_AXIMM_66_AWREADY = ap_AWREADY[66];
            assign ap_WDATA[66][M_AXIMM_66_DATA_WIDTH-1:0] = AP_AXIMM_66_WDATA;
            assign ap_WSTRB[66][M_AXIMM_66_DATA_WIDTH/8-1:0] = AP_AXIMM_66_WSTRB;
            assign ap_WLAST[66] = AP_AXIMM_66_WLAST;
            assign ap_WVALID[66] = AP_AXIMM_66_WVALID;
            assign AP_AXIMM_66_WREADY = ap_WREADY[66];
            assign AP_AXIMM_66_BRESP = ap_BRESP[66];
            assign AP_AXIMM_66_BVALID = ap_BVALID[66];
            assign ap_BREADY[66] = AP_AXIMM_66_BREADY;
            assign ap_ARADDR[66][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_66_ARADDR;
            assign ap_ARLEN[66] = AP_AXIMM_66_ARLEN;
            assign ap_ARSIZE[66] = AP_AXIMM_66_ARSIZE;
            assign ap_ARBURST[66] = AP_AXIMM_66_ARBURST;
            assign ap_ARLOCK[66] = AP_AXIMM_66_ARLOCK;
            assign ap_ARCACHE[66] = AP_AXIMM_66_ARCACHE;
            assign ap_ARPROT[66] = AP_AXIMM_66_ARPROT;
            assign ap_ARREGION[66] = AP_AXIMM_66_ARREGION;
            assign ap_ARQOS[66] = AP_AXIMM_66_ARQOS;
            assign ap_ARVALID[66] = AP_AXIMM_66_ARVALID;
            assign AP_AXIMM_66_ARREADY = ap_ARREADY[66];
            assign AP_AXIMM_66_RDATA = ap_RDATA[66][M_AXIMM_66_DATA_WIDTH-1:0];
            assign AP_AXIMM_66_RRESP = ap_RRESP[66];
            assign AP_AXIMM_66_RLAST = ap_RLAST[66];
            assign AP_AXIMM_66_RVALID = ap_RVALID[66];
            assign ap_RREADY[66] = AP_AXIMM_66_RREADY;
            assign M_AXIMM_66_AWADDR = dm_AWADDR[66][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_66_AWLEN = dm_AWLEN[66];
            assign M_AXIMM_66_AWSIZE = dm_AWSIZE[66];
            assign M_AXIMM_66_AWBURST = dm_AWBURST[66];
            assign M_AXIMM_66_AWLOCK = dm_AWLOCK[66];
            assign M_AXIMM_66_AWCACHE = dm_AWCACHE[66];
            assign M_AXIMM_66_AWPROT = dm_AWPROT[66];
            assign M_AXIMM_66_AWREGION = dm_AWREGION[66];
            assign M_AXIMM_66_AWQOS = dm_AWQOS[66];
            assign M_AXIMM_66_AWVALID = dm_AWVALID[66];
            assign dm_AWREADY[66] = M_AXIMM_66_AWREADY;
            assign M_AXIMM_66_WDATA = dm_WDATA[66][M_AXIMM_66_DATA_WIDTH-1:0];
            assign M_AXIMM_66_WSTRB = dm_WSTRB[66][M_AXIMM_66_DATA_WIDTH/8-1:0];
            assign M_AXIMM_66_WLAST = dm_WLAST[66];
            assign M_AXIMM_66_WVALID = dm_WVALID[66];
            assign dm_WREADY[66] = M_AXIMM_66_WREADY;
            assign dm_BRESP[66] = M_AXIMM_66_BRESP;
            assign dm_BVALID[66] = M_AXIMM_66_BVALID;
            assign M_AXIMM_66_BREADY = dm_BREADY[66];
            assign M_AXIMM_66_ARADDR = dm_ARADDR[66][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_66_ARLEN = dm_ARLEN[66];
            assign M_AXIMM_66_ARSIZE = dm_ARSIZE[66];
            assign M_AXIMM_66_ARBURST = dm_ARBURST[66];
            assign M_AXIMM_66_ARLOCK = dm_ARLOCK[66];
            assign M_AXIMM_66_ARCACHE = dm_ARCACHE[66];
            assign M_AXIMM_66_ARPROT = dm_ARPROT[66];
            assign M_AXIMM_66_ARREGION = dm_ARREGION[66];
            assign M_AXIMM_66_ARQOS = dm_ARQOS[66];
            assign M_AXIMM_66_ARVALID = dm_ARVALID[66];
            assign dm_ARREADY[66] = M_AXIMM_66_ARREADY;
            assign dm_RDATA[66][M_AXIMM_66_DATA_WIDTH-1:0] = M_AXIMM_66_RDATA;
            assign dm_RRESP[66] = M_AXIMM_66_RRESP;
            assign dm_RLAST[66] = M_AXIMM_66_RLAST;
            assign dm_RVALID[66] = M_AXIMM_66_RVALID;
            assign M_AXIMM_66_RREADY = dm_RREADY[66];
        end
        if(C_NUM_AXIMMs > 67) begin
            assign ap_AWADDR[67][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_67_AWADDR;
            assign ap_AWLEN[67] = AP_AXIMM_67_AWLEN;
            assign ap_AWSIZE[67] = AP_AXIMM_67_AWSIZE;
            assign ap_AWBURST[67] = AP_AXIMM_67_AWBURST;
            assign ap_AWLOCK[67] = AP_AXIMM_67_AWLOCK;
            assign ap_AWCACHE[67] = AP_AXIMM_67_AWCACHE;
            assign ap_AWPROT[67] = AP_AXIMM_67_AWPROT;
            assign ap_AWREGION[67] = AP_AXIMM_67_AWREGION;
            assign ap_AWQOS[67] = AP_AXIMM_67_AWQOS;
            assign ap_AWVALID[67] = AP_AXIMM_67_AWVALID;
            assign AP_AXIMM_67_AWREADY = ap_AWREADY[67];
            assign ap_WDATA[67][M_AXIMM_67_DATA_WIDTH-1:0] = AP_AXIMM_67_WDATA;
            assign ap_WSTRB[67][M_AXIMM_67_DATA_WIDTH/8-1:0] = AP_AXIMM_67_WSTRB;
            assign ap_WLAST[67] = AP_AXIMM_67_WLAST;
            assign ap_WVALID[67] = AP_AXIMM_67_WVALID;
            assign AP_AXIMM_67_WREADY = ap_WREADY[67];
            assign AP_AXIMM_67_BRESP = ap_BRESP[67];
            assign AP_AXIMM_67_BVALID = ap_BVALID[67];
            assign ap_BREADY[67] = AP_AXIMM_67_BREADY;
            assign ap_ARADDR[67][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_67_ARADDR;
            assign ap_ARLEN[67] = AP_AXIMM_67_ARLEN;
            assign ap_ARSIZE[67] = AP_AXIMM_67_ARSIZE;
            assign ap_ARBURST[67] = AP_AXIMM_67_ARBURST;
            assign ap_ARLOCK[67] = AP_AXIMM_67_ARLOCK;
            assign ap_ARCACHE[67] = AP_AXIMM_67_ARCACHE;
            assign ap_ARPROT[67] = AP_AXIMM_67_ARPROT;
            assign ap_ARREGION[67] = AP_AXIMM_67_ARREGION;
            assign ap_ARQOS[67] = AP_AXIMM_67_ARQOS;
            assign ap_ARVALID[67] = AP_AXIMM_67_ARVALID;
            assign AP_AXIMM_67_ARREADY = ap_ARREADY[67];
            assign AP_AXIMM_67_RDATA = ap_RDATA[67][M_AXIMM_67_DATA_WIDTH-1:0];
            assign AP_AXIMM_67_RRESP = ap_RRESP[67];
            assign AP_AXIMM_67_RLAST = ap_RLAST[67];
            assign AP_AXIMM_67_RVALID = ap_RVALID[67];
            assign ap_RREADY[67] = AP_AXIMM_67_RREADY;
            assign M_AXIMM_67_AWADDR = dm_AWADDR[67][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_67_AWLEN = dm_AWLEN[67];
            assign M_AXIMM_67_AWSIZE = dm_AWSIZE[67];
            assign M_AXIMM_67_AWBURST = dm_AWBURST[67];
            assign M_AXIMM_67_AWLOCK = dm_AWLOCK[67];
            assign M_AXIMM_67_AWCACHE = dm_AWCACHE[67];
            assign M_AXIMM_67_AWPROT = dm_AWPROT[67];
            assign M_AXIMM_67_AWREGION = dm_AWREGION[67];
            assign M_AXIMM_67_AWQOS = dm_AWQOS[67];
            assign M_AXIMM_67_AWVALID = dm_AWVALID[67];
            assign dm_AWREADY[67] = M_AXIMM_67_AWREADY;
            assign M_AXIMM_67_WDATA = dm_WDATA[67][M_AXIMM_67_DATA_WIDTH-1:0];
            assign M_AXIMM_67_WSTRB = dm_WSTRB[67][M_AXIMM_67_DATA_WIDTH/8-1:0];
            assign M_AXIMM_67_WLAST = dm_WLAST[67];
            assign M_AXIMM_67_WVALID = dm_WVALID[67];
            assign dm_WREADY[67] = M_AXIMM_67_WREADY;
            assign dm_BRESP[67] = M_AXIMM_67_BRESP;
            assign dm_BVALID[67] = M_AXIMM_67_BVALID;
            assign M_AXIMM_67_BREADY = dm_BREADY[67];
            assign M_AXIMM_67_ARADDR = dm_ARADDR[67][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_67_ARLEN = dm_ARLEN[67];
            assign M_AXIMM_67_ARSIZE = dm_ARSIZE[67];
            assign M_AXIMM_67_ARBURST = dm_ARBURST[67];
            assign M_AXIMM_67_ARLOCK = dm_ARLOCK[67];
            assign M_AXIMM_67_ARCACHE = dm_ARCACHE[67];
            assign M_AXIMM_67_ARPROT = dm_ARPROT[67];
            assign M_AXIMM_67_ARREGION = dm_ARREGION[67];
            assign M_AXIMM_67_ARQOS = dm_ARQOS[67];
            assign M_AXIMM_67_ARVALID = dm_ARVALID[67];
            assign dm_ARREADY[67] = M_AXIMM_67_ARREADY;
            assign dm_RDATA[67][M_AXIMM_67_DATA_WIDTH-1:0] = M_AXIMM_67_RDATA;
            assign dm_RRESP[67] = M_AXIMM_67_RRESP;
            assign dm_RLAST[67] = M_AXIMM_67_RLAST;
            assign dm_RVALID[67] = M_AXIMM_67_RVALID;
            assign M_AXIMM_67_RREADY = dm_RREADY[67];
        end
        if(C_NUM_AXIMMs > 68) begin
            assign ap_AWADDR[68][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_68_AWADDR;
            assign ap_AWLEN[68] = AP_AXIMM_68_AWLEN;
            assign ap_AWSIZE[68] = AP_AXIMM_68_AWSIZE;
            assign ap_AWBURST[68] = AP_AXIMM_68_AWBURST;
            assign ap_AWLOCK[68] = AP_AXIMM_68_AWLOCK;
            assign ap_AWCACHE[68] = AP_AXIMM_68_AWCACHE;
            assign ap_AWPROT[68] = AP_AXIMM_68_AWPROT;
            assign ap_AWREGION[68] = AP_AXIMM_68_AWREGION;
            assign ap_AWQOS[68] = AP_AXIMM_68_AWQOS;
            assign ap_AWVALID[68] = AP_AXIMM_68_AWVALID;
            assign AP_AXIMM_68_AWREADY = ap_AWREADY[68];
            assign ap_WDATA[68][M_AXIMM_68_DATA_WIDTH-1:0] = AP_AXIMM_68_WDATA;
            assign ap_WSTRB[68][M_AXIMM_68_DATA_WIDTH/8-1:0] = AP_AXIMM_68_WSTRB;
            assign ap_WLAST[68] = AP_AXIMM_68_WLAST;
            assign ap_WVALID[68] = AP_AXIMM_68_WVALID;
            assign AP_AXIMM_68_WREADY = ap_WREADY[68];
            assign AP_AXIMM_68_BRESP = ap_BRESP[68];
            assign AP_AXIMM_68_BVALID = ap_BVALID[68];
            assign ap_BREADY[68] = AP_AXIMM_68_BREADY;
            assign ap_ARADDR[68][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_68_ARADDR;
            assign ap_ARLEN[68] = AP_AXIMM_68_ARLEN;
            assign ap_ARSIZE[68] = AP_AXIMM_68_ARSIZE;
            assign ap_ARBURST[68] = AP_AXIMM_68_ARBURST;
            assign ap_ARLOCK[68] = AP_AXIMM_68_ARLOCK;
            assign ap_ARCACHE[68] = AP_AXIMM_68_ARCACHE;
            assign ap_ARPROT[68] = AP_AXIMM_68_ARPROT;
            assign ap_ARREGION[68] = AP_AXIMM_68_ARREGION;
            assign ap_ARQOS[68] = AP_AXIMM_68_ARQOS;
            assign ap_ARVALID[68] = AP_AXIMM_68_ARVALID;
            assign AP_AXIMM_68_ARREADY = ap_ARREADY[68];
            assign AP_AXIMM_68_RDATA = ap_RDATA[68][M_AXIMM_68_DATA_WIDTH-1:0];
            assign AP_AXIMM_68_RRESP = ap_RRESP[68];
            assign AP_AXIMM_68_RLAST = ap_RLAST[68];
            assign AP_AXIMM_68_RVALID = ap_RVALID[68];
            assign ap_RREADY[68] = AP_AXIMM_68_RREADY;
            assign M_AXIMM_68_AWADDR = dm_AWADDR[68][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_68_AWLEN = dm_AWLEN[68];
            assign M_AXIMM_68_AWSIZE = dm_AWSIZE[68];
            assign M_AXIMM_68_AWBURST = dm_AWBURST[68];
            assign M_AXIMM_68_AWLOCK = dm_AWLOCK[68];
            assign M_AXIMM_68_AWCACHE = dm_AWCACHE[68];
            assign M_AXIMM_68_AWPROT = dm_AWPROT[68];
            assign M_AXIMM_68_AWREGION = dm_AWREGION[68];
            assign M_AXIMM_68_AWQOS = dm_AWQOS[68];
            assign M_AXIMM_68_AWVALID = dm_AWVALID[68];
            assign dm_AWREADY[68] = M_AXIMM_68_AWREADY;
            assign M_AXIMM_68_WDATA = dm_WDATA[68][M_AXIMM_68_DATA_WIDTH-1:0];
            assign M_AXIMM_68_WSTRB = dm_WSTRB[68][M_AXIMM_68_DATA_WIDTH/8-1:0];
            assign M_AXIMM_68_WLAST = dm_WLAST[68];
            assign M_AXIMM_68_WVALID = dm_WVALID[68];
            assign dm_WREADY[68] = M_AXIMM_68_WREADY;
            assign dm_BRESP[68] = M_AXIMM_68_BRESP;
            assign dm_BVALID[68] = M_AXIMM_68_BVALID;
            assign M_AXIMM_68_BREADY = dm_BREADY[68];
            assign M_AXIMM_68_ARADDR = dm_ARADDR[68][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_68_ARLEN = dm_ARLEN[68];
            assign M_AXIMM_68_ARSIZE = dm_ARSIZE[68];
            assign M_AXIMM_68_ARBURST = dm_ARBURST[68];
            assign M_AXIMM_68_ARLOCK = dm_ARLOCK[68];
            assign M_AXIMM_68_ARCACHE = dm_ARCACHE[68];
            assign M_AXIMM_68_ARPROT = dm_ARPROT[68];
            assign M_AXIMM_68_ARREGION = dm_ARREGION[68];
            assign M_AXIMM_68_ARQOS = dm_ARQOS[68];
            assign M_AXIMM_68_ARVALID = dm_ARVALID[68];
            assign dm_ARREADY[68] = M_AXIMM_68_ARREADY;
            assign dm_RDATA[68][M_AXIMM_68_DATA_WIDTH-1:0] = M_AXIMM_68_RDATA;
            assign dm_RRESP[68] = M_AXIMM_68_RRESP;
            assign dm_RLAST[68] = M_AXIMM_68_RLAST;
            assign dm_RVALID[68] = M_AXIMM_68_RVALID;
            assign M_AXIMM_68_RREADY = dm_RREADY[68];
        end
        if(C_NUM_AXIMMs > 69) begin
            assign ap_AWADDR[69][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_69_AWADDR;
            assign ap_AWLEN[69] = AP_AXIMM_69_AWLEN;
            assign ap_AWSIZE[69] = AP_AXIMM_69_AWSIZE;
            assign ap_AWBURST[69] = AP_AXIMM_69_AWBURST;
            assign ap_AWLOCK[69] = AP_AXIMM_69_AWLOCK;
            assign ap_AWCACHE[69] = AP_AXIMM_69_AWCACHE;
            assign ap_AWPROT[69] = AP_AXIMM_69_AWPROT;
            assign ap_AWREGION[69] = AP_AXIMM_69_AWREGION;
            assign ap_AWQOS[69] = AP_AXIMM_69_AWQOS;
            assign ap_AWVALID[69] = AP_AXIMM_69_AWVALID;
            assign AP_AXIMM_69_AWREADY = ap_AWREADY[69];
            assign ap_WDATA[69][M_AXIMM_69_DATA_WIDTH-1:0] = AP_AXIMM_69_WDATA;
            assign ap_WSTRB[69][M_AXIMM_69_DATA_WIDTH/8-1:0] = AP_AXIMM_69_WSTRB;
            assign ap_WLAST[69] = AP_AXIMM_69_WLAST;
            assign ap_WVALID[69] = AP_AXIMM_69_WVALID;
            assign AP_AXIMM_69_WREADY = ap_WREADY[69];
            assign AP_AXIMM_69_BRESP = ap_BRESP[69];
            assign AP_AXIMM_69_BVALID = ap_BVALID[69];
            assign ap_BREADY[69] = AP_AXIMM_69_BREADY;
            assign ap_ARADDR[69][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_69_ARADDR;
            assign ap_ARLEN[69] = AP_AXIMM_69_ARLEN;
            assign ap_ARSIZE[69] = AP_AXIMM_69_ARSIZE;
            assign ap_ARBURST[69] = AP_AXIMM_69_ARBURST;
            assign ap_ARLOCK[69] = AP_AXIMM_69_ARLOCK;
            assign ap_ARCACHE[69] = AP_AXIMM_69_ARCACHE;
            assign ap_ARPROT[69] = AP_AXIMM_69_ARPROT;
            assign ap_ARREGION[69] = AP_AXIMM_69_ARREGION;
            assign ap_ARQOS[69] = AP_AXIMM_69_ARQOS;
            assign ap_ARVALID[69] = AP_AXIMM_69_ARVALID;
            assign AP_AXIMM_69_ARREADY = ap_ARREADY[69];
            assign AP_AXIMM_69_RDATA = ap_RDATA[69][M_AXIMM_69_DATA_WIDTH-1:0];
            assign AP_AXIMM_69_RRESP = ap_RRESP[69];
            assign AP_AXIMM_69_RLAST = ap_RLAST[69];
            assign AP_AXIMM_69_RVALID = ap_RVALID[69];
            assign ap_RREADY[69] = AP_AXIMM_69_RREADY;
            assign M_AXIMM_69_AWADDR = dm_AWADDR[69][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_69_AWLEN = dm_AWLEN[69];
            assign M_AXIMM_69_AWSIZE = dm_AWSIZE[69];
            assign M_AXIMM_69_AWBURST = dm_AWBURST[69];
            assign M_AXIMM_69_AWLOCK = dm_AWLOCK[69];
            assign M_AXIMM_69_AWCACHE = dm_AWCACHE[69];
            assign M_AXIMM_69_AWPROT = dm_AWPROT[69];
            assign M_AXIMM_69_AWREGION = dm_AWREGION[69];
            assign M_AXIMM_69_AWQOS = dm_AWQOS[69];
            assign M_AXIMM_69_AWVALID = dm_AWVALID[69];
            assign dm_AWREADY[69] = M_AXIMM_69_AWREADY;
            assign M_AXIMM_69_WDATA = dm_WDATA[69][M_AXIMM_69_DATA_WIDTH-1:0];
            assign M_AXIMM_69_WSTRB = dm_WSTRB[69][M_AXIMM_69_DATA_WIDTH/8-1:0];
            assign M_AXIMM_69_WLAST = dm_WLAST[69];
            assign M_AXIMM_69_WVALID = dm_WVALID[69];
            assign dm_WREADY[69] = M_AXIMM_69_WREADY;
            assign dm_BRESP[69] = M_AXIMM_69_BRESP;
            assign dm_BVALID[69] = M_AXIMM_69_BVALID;
            assign M_AXIMM_69_BREADY = dm_BREADY[69];
            assign M_AXIMM_69_ARADDR = dm_ARADDR[69][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_69_ARLEN = dm_ARLEN[69];
            assign M_AXIMM_69_ARSIZE = dm_ARSIZE[69];
            assign M_AXIMM_69_ARBURST = dm_ARBURST[69];
            assign M_AXIMM_69_ARLOCK = dm_ARLOCK[69];
            assign M_AXIMM_69_ARCACHE = dm_ARCACHE[69];
            assign M_AXIMM_69_ARPROT = dm_ARPROT[69];
            assign M_AXIMM_69_ARREGION = dm_ARREGION[69];
            assign M_AXIMM_69_ARQOS = dm_ARQOS[69];
            assign M_AXIMM_69_ARVALID = dm_ARVALID[69];
            assign dm_ARREADY[69] = M_AXIMM_69_ARREADY;
            assign dm_RDATA[69][M_AXIMM_69_DATA_WIDTH-1:0] = M_AXIMM_69_RDATA;
            assign dm_RRESP[69] = M_AXIMM_69_RRESP;
            assign dm_RLAST[69] = M_AXIMM_69_RLAST;
            assign dm_RVALID[69] = M_AXIMM_69_RVALID;
            assign M_AXIMM_69_RREADY = dm_RREADY[69];
        end
        if(C_NUM_AXIMMs > 70) begin
            assign ap_AWADDR[70][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_70_AWADDR;
            assign ap_AWLEN[70] = AP_AXIMM_70_AWLEN;
            assign ap_AWSIZE[70] = AP_AXIMM_70_AWSIZE;
            assign ap_AWBURST[70] = AP_AXIMM_70_AWBURST;
            assign ap_AWLOCK[70] = AP_AXIMM_70_AWLOCK;
            assign ap_AWCACHE[70] = AP_AXIMM_70_AWCACHE;
            assign ap_AWPROT[70] = AP_AXIMM_70_AWPROT;
            assign ap_AWREGION[70] = AP_AXIMM_70_AWREGION;
            assign ap_AWQOS[70] = AP_AXIMM_70_AWQOS;
            assign ap_AWVALID[70] = AP_AXIMM_70_AWVALID;
            assign AP_AXIMM_70_AWREADY = ap_AWREADY[70];
            assign ap_WDATA[70][M_AXIMM_70_DATA_WIDTH-1:0] = AP_AXIMM_70_WDATA;
            assign ap_WSTRB[70][M_AXIMM_70_DATA_WIDTH/8-1:0] = AP_AXIMM_70_WSTRB;
            assign ap_WLAST[70] = AP_AXIMM_70_WLAST;
            assign ap_WVALID[70] = AP_AXIMM_70_WVALID;
            assign AP_AXIMM_70_WREADY = ap_WREADY[70];
            assign AP_AXIMM_70_BRESP = ap_BRESP[70];
            assign AP_AXIMM_70_BVALID = ap_BVALID[70];
            assign ap_BREADY[70] = AP_AXIMM_70_BREADY;
            assign ap_ARADDR[70][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_70_ARADDR;
            assign ap_ARLEN[70] = AP_AXIMM_70_ARLEN;
            assign ap_ARSIZE[70] = AP_AXIMM_70_ARSIZE;
            assign ap_ARBURST[70] = AP_AXIMM_70_ARBURST;
            assign ap_ARLOCK[70] = AP_AXIMM_70_ARLOCK;
            assign ap_ARCACHE[70] = AP_AXIMM_70_ARCACHE;
            assign ap_ARPROT[70] = AP_AXIMM_70_ARPROT;
            assign ap_ARREGION[70] = AP_AXIMM_70_ARREGION;
            assign ap_ARQOS[70] = AP_AXIMM_70_ARQOS;
            assign ap_ARVALID[70] = AP_AXIMM_70_ARVALID;
            assign AP_AXIMM_70_ARREADY = ap_ARREADY[70];
            assign AP_AXIMM_70_RDATA = ap_RDATA[70][M_AXIMM_70_DATA_WIDTH-1:0];
            assign AP_AXIMM_70_RRESP = ap_RRESP[70];
            assign AP_AXIMM_70_RLAST = ap_RLAST[70];
            assign AP_AXIMM_70_RVALID = ap_RVALID[70];
            assign ap_RREADY[70] = AP_AXIMM_70_RREADY;
            assign M_AXIMM_70_AWADDR = dm_AWADDR[70][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_70_AWLEN = dm_AWLEN[70];
            assign M_AXIMM_70_AWSIZE = dm_AWSIZE[70];
            assign M_AXIMM_70_AWBURST = dm_AWBURST[70];
            assign M_AXIMM_70_AWLOCK = dm_AWLOCK[70];
            assign M_AXIMM_70_AWCACHE = dm_AWCACHE[70];
            assign M_AXIMM_70_AWPROT = dm_AWPROT[70];
            assign M_AXIMM_70_AWREGION = dm_AWREGION[70];
            assign M_AXIMM_70_AWQOS = dm_AWQOS[70];
            assign M_AXIMM_70_AWVALID = dm_AWVALID[70];
            assign dm_AWREADY[70] = M_AXIMM_70_AWREADY;
            assign M_AXIMM_70_WDATA = dm_WDATA[70][M_AXIMM_70_DATA_WIDTH-1:0];
            assign M_AXIMM_70_WSTRB = dm_WSTRB[70][M_AXIMM_70_DATA_WIDTH/8-1:0];
            assign M_AXIMM_70_WLAST = dm_WLAST[70];
            assign M_AXIMM_70_WVALID = dm_WVALID[70];
            assign dm_WREADY[70] = M_AXIMM_70_WREADY;
            assign dm_BRESP[70] = M_AXIMM_70_BRESP;
            assign dm_BVALID[70] = M_AXIMM_70_BVALID;
            assign M_AXIMM_70_BREADY = dm_BREADY[70];
            assign M_AXIMM_70_ARADDR = dm_ARADDR[70][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_70_ARLEN = dm_ARLEN[70];
            assign M_AXIMM_70_ARSIZE = dm_ARSIZE[70];
            assign M_AXIMM_70_ARBURST = dm_ARBURST[70];
            assign M_AXIMM_70_ARLOCK = dm_ARLOCK[70];
            assign M_AXIMM_70_ARCACHE = dm_ARCACHE[70];
            assign M_AXIMM_70_ARPROT = dm_ARPROT[70];
            assign M_AXIMM_70_ARREGION = dm_ARREGION[70];
            assign M_AXIMM_70_ARQOS = dm_ARQOS[70];
            assign M_AXIMM_70_ARVALID = dm_ARVALID[70];
            assign dm_ARREADY[70] = M_AXIMM_70_ARREADY;
            assign dm_RDATA[70][M_AXIMM_70_DATA_WIDTH-1:0] = M_AXIMM_70_RDATA;
            assign dm_RRESP[70] = M_AXIMM_70_RRESP;
            assign dm_RLAST[70] = M_AXIMM_70_RLAST;
            assign dm_RVALID[70] = M_AXIMM_70_RVALID;
            assign M_AXIMM_70_RREADY = dm_RREADY[70];
        end
        if(C_NUM_AXIMMs > 71) begin
            assign ap_AWADDR[71][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_71_AWADDR;
            assign ap_AWLEN[71] = AP_AXIMM_71_AWLEN;
            assign ap_AWSIZE[71] = AP_AXIMM_71_AWSIZE;
            assign ap_AWBURST[71] = AP_AXIMM_71_AWBURST;
            assign ap_AWLOCK[71] = AP_AXIMM_71_AWLOCK;
            assign ap_AWCACHE[71] = AP_AXIMM_71_AWCACHE;
            assign ap_AWPROT[71] = AP_AXIMM_71_AWPROT;
            assign ap_AWREGION[71] = AP_AXIMM_71_AWREGION;
            assign ap_AWQOS[71] = AP_AXIMM_71_AWQOS;
            assign ap_AWVALID[71] = AP_AXIMM_71_AWVALID;
            assign AP_AXIMM_71_AWREADY = ap_AWREADY[71];
            assign ap_WDATA[71][M_AXIMM_71_DATA_WIDTH-1:0] = AP_AXIMM_71_WDATA;
            assign ap_WSTRB[71][M_AXIMM_71_DATA_WIDTH/8-1:0] = AP_AXIMM_71_WSTRB;
            assign ap_WLAST[71] = AP_AXIMM_71_WLAST;
            assign ap_WVALID[71] = AP_AXIMM_71_WVALID;
            assign AP_AXIMM_71_WREADY = ap_WREADY[71];
            assign AP_AXIMM_71_BRESP = ap_BRESP[71];
            assign AP_AXIMM_71_BVALID = ap_BVALID[71];
            assign ap_BREADY[71] = AP_AXIMM_71_BREADY;
            assign ap_ARADDR[71][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_71_ARADDR;
            assign ap_ARLEN[71] = AP_AXIMM_71_ARLEN;
            assign ap_ARSIZE[71] = AP_AXIMM_71_ARSIZE;
            assign ap_ARBURST[71] = AP_AXIMM_71_ARBURST;
            assign ap_ARLOCK[71] = AP_AXIMM_71_ARLOCK;
            assign ap_ARCACHE[71] = AP_AXIMM_71_ARCACHE;
            assign ap_ARPROT[71] = AP_AXIMM_71_ARPROT;
            assign ap_ARREGION[71] = AP_AXIMM_71_ARREGION;
            assign ap_ARQOS[71] = AP_AXIMM_71_ARQOS;
            assign ap_ARVALID[71] = AP_AXIMM_71_ARVALID;
            assign AP_AXIMM_71_ARREADY = ap_ARREADY[71];
            assign AP_AXIMM_71_RDATA = ap_RDATA[71][M_AXIMM_71_DATA_WIDTH-1:0];
            assign AP_AXIMM_71_RRESP = ap_RRESP[71];
            assign AP_AXIMM_71_RLAST = ap_RLAST[71];
            assign AP_AXIMM_71_RVALID = ap_RVALID[71];
            assign ap_RREADY[71] = AP_AXIMM_71_RREADY;
            assign M_AXIMM_71_AWADDR = dm_AWADDR[71][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_71_AWLEN = dm_AWLEN[71];
            assign M_AXIMM_71_AWSIZE = dm_AWSIZE[71];
            assign M_AXIMM_71_AWBURST = dm_AWBURST[71];
            assign M_AXIMM_71_AWLOCK = dm_AWLOCK[71];
            assign M_AXIMM_71_AWCACHE = dm_AWCACHE[71];
            assign M_AXIMM_71_AWPROT = dm_AWPROT[71];
            assign M_AXIMM_71_AWREGION = dm_AWREGION[71];
            assign M_AXIMM_71_AWQOS = dm_AWQOS[71];
            assign M_AXIMM_71_AWVALID = dm_AWVALID[71];
            assign dm_AWREADY[71] = M_AXIMM_71_AWREADY;
            assign M_AXIMM_71_WDATA = dm_WDATA[71][M_AXIMM_71_DATA_WIDTH-1:0];
            assign M_AXIMM_71_WSTRB = dm_WSTRB[71][M_AXIMM_71_DATA_WIDTH/8-1:0];
            assign M_AXIMM_71_WLAST = dm_WLAST[71];
            assign M_AXIMM_71_WVALID = dm_WVALID[71];
            assign dm_WREADY[71] = M_AXIMM_71_WREADY;
            assign dm_BRESP[71] = M_AXIMM_71_BRESP;
            assign dm_BVALID[71] = M_AXIMM_71_BVALID;
            assign M_AXIMM_71_BREADY = dm_BREADY[71];
            assign M_AXIMM_71_ARADDR = dm_ARADDR[71][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_71_ARLEN = dm_ARLEN[71];
            assign M_AXIMM_71_ARSIZE = dm_ARSIZE[71];
            assign M_AXIMM_71_ARBURST = dm_ARBURST[71];
            assign M_AXIMM_71_ARLOCK = dm_ARLOCK[71];
            assign M_AXIMM_71_ARCACHE = dm_ARCACHE[71];
            assign M_AXIMM_71_ARPROT = dm_ARPROT[71];
            assign M_AXIMM_71_ARREGION = dm_ARREGION[71];
            assign M_AXIMM_71_ARQOS = dm_ARQOS[71];
            assign M_AXIMM_71_ARVALID = dm_ARVALID[71];
            assign dm_ARREADY[71] = M_AXIMM_71_ARREADY;
            assign dm_RDATA[71][M_AXIMM_71_DATA_WIDTH-1:0] = M_AXIMM_71_RDATA;
            assign dm_RRESP[71] = M_AXIMM_71_RRESP;
            assign dm_RLAST[71] = M_AXIMM_71_RLAST;
            assign dm_RVALID[71] = M_AXIMM_71_RVALID;
            assign M_AXIMM_71_RREADY = dm_RREADY[71];
        end
        if(C_NUM_AXIMMs > 72) begin
            assign ap_AWADDR[72][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_72_AWADDR;
            assign ap_AWLEN[72] = AP_AXIMM_72_AWLEN;
            assign ap_AWSIZE[72] = AP_AXIMM_72_AWSIZE;
            assign ap_AWBURST[72] = AP_AXIMM_72_AWBURST;
            assign ap_AWLOCK[72] = AP_AXIMM_72_AWLOCK;
            assign ap_AWCACHE[72] = AP_AXIMM_72_AWCACHE;
            assign ap_AWPROT[72] = AP_AXIMM_72_AWPROT;
            assign ap_AWREGION[72] = AP_AXIMM_72_AWREGION;
            assign ap_AWQOS[72] = AP_AXIMM_72_AWQOS;
            assign ap_AWVALID[72] = AP_AXIMM_72_AWVALID;
            assign AP_AXIMM_72_AWREADY = ap_AWREADY[72];
            assign ap_WDATA[72][M_AXIMM_72_DATA_WIDTH-1:0] = AP_AXIMM_72_WDATA;
            assign ap_WSTRB[72][M_AXIMM_72_DATA_WIDTH/8-1:0] = AP_AXIMM_72_WSTRB;
            assign ap_WLAST[72] = AP_AXIMM_72_WLAST;
            assign ap_WVALID[72] = AP_AXIMM_72_WVALID;
            assign AP_AXIMM_72_WREADY = ap_WREADY[72];
            assign AP_AXIMM_72_BRESP = ap_BRESP[72];
            assign AP_AXIMM_72_BVALID = ap_BVALID[72];
            assign ap_BREADY[72] = AP_AXIMM_72_BREADY;
            assign ap_ARADDR[72][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_72_ARADDR;
            assign ap_ARLEN[72] = AP_AXIMM_72_ARLEN;
            assign ap_ARSIZE[72] = AP_AXIMM_72_ARSIZE;
            assign ap_ARBURST[72] = AP_AXIMM_72_ARBURST;
            assign ap_ARLOCK[72] = AP_AXIMM_72_ARLOCK;
            assign ap_ARCACHE[72] = AP_AXIMM_72_ARCACHE;
            assign ap_ARPROT[72] = AP_AXIMM_72_ARPROT;
            assign ap_ARREGION[72] = AP_AXIMM_72_ARREGION;
            assign ap_ARQOS[72] = AP_AXIMM_72_ARQOS;
            assign ap_ARVALID[72] = AP_AXIMM_72_ARVALID;
            assign AP_AXIMM_72_ARREADY = ap_ARREADY[72];
            assign AP_AXIMM_72_RDATA = ap_RDATA[72][M_AXIMM_72_DATA_WIDTH-1:0];
            assign AP_AXIMM_72_RRESP = ap_RRESP[72];
            assign AP_AXIMM_72_RLAST = ap_RLAST[72];
            assign AP_AXIMM_72_RVALID = ap_RVALID[72];
            assign ap_RREADY[72] = AP_AXIMM_72_RREADY;
            assign M_AXIMM_72_AWADDR = dm_AWADDR[72][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_72_AWLEN = dm_AWLEN[72];
            assign M_AXIMM_72_AWSIZE = dm_AWSIZE[72];
            assign M_AXIMM_72_AWBURST = dm_AWBURST[72];
            assign M_AXIMM_72_AWLOCK = dm_AWLOCK[72];
            assign M_AXIMM_72_AWCACHE = dm_AWCACHE[72];
            assign M_AXIMM_72_AWPROT = dm_AWPROT[72];
            assign M_AXIMM_72_AWREGION = dm_AWREGION[72];
            assign M_AXIMM_72_AWQOS = dm_AWQOS[72];
            assign M_AXIMM_72_AWVALID = dm_AWVALID[72];
            assign dm_AWREADY[72] = M_AXIMM_72_AWREADY;
            assign M_AXIMM_72_WDATA = dm_WDATA[72][M_AXIMM_72_DATA_WIDTH-1:0];
            assign M_AXIMM_72_WSTRB = dm_WSTRB[72][M_AXIMM_72_DATA_WIDTH/8-1:0];
            assign M_AXIMM_72_WLAST = dm_WLAST[72];
            assign M_AXIMM_72_WVALID = dm_WVALID[72];
            assign dm_WREADY[72] = M_AXIMM_72_WREADY;
            assign dm_BRESP[72] = M_AXIMM_72_BRESP;
            assign dm_BVALID[72] = M_AXIMM_72_BVALID;
            assign M_AXIMM_72_BREADY = dm_BREADY[72];
            assign M_AXIMM_72_ARADDR = dm_ARADDR[72][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_72_ARLEN = dm_ARLEN[72];
            assign M_AXIMM_72_ARSIZE = dm_ARSIZE[72];
            assign M_AXIMM_72_ARBURST = dm_ARBURST[72];
            assign M_AXIMM_72_ARLOCK = dm_ARLOCK[72];
            assign M_AXIMM_72_ARCACHE = dm_ARCACHE[72];
            assign M_AXIMM_72_ARPROT = dm_ARPROT[72];
            assign M_AXIMM_72_ARREGION = dm_ARREGION[72];
            assign M_AXIMM_72_ARQOS = dm_ARQOS[72];
            assign M_AXIMM_72_ARVALID = dm_ARVALID[72];
            assign dm_ARREADY[72] = M_AXIMM_72_ARREADY;
            assign dm_RDATA[72][M_AXIMM_72_DATA_WIDTH-1:0] = M_AXIMM_72_RDATA;
            assign dm_RRESP[72] = M_AXIMM_72_RRESP;
            assign dm_RLAST[72] = M_AXIMM_72_RLAST;
            assign dm_RVALID[72] = M_AXIMM_72_RVALID;
            assign M_AXIMM_72_RREADY = dm_RREADY[72];
        end
        if(C_NUM_AXIMMs > 73) begin
            assign ap_AWADDR[73][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_73_AWADDR;
            assign ap_AWLEN[73] = AP_AXIMM_73_AWLEN;
            assign ap_AWSIZE[73] = AP_AXIMM_73_AWSIZE;
            assign ap_AWBURST[73] = AP_AXIMM_73_AWBURST;
            assign ap_AWLOCK[73] = AP_AXIMM_73_AWLOCK;
            assign ap_AWCACHE[73] = AP_AXIMM_73_AWCACHE;
            assign ap_AWPROT[73] = AP_AXIMM_73_AWPROT;
            assign ap_AWREGION[73] = AP_AXIMM_73_AWREGION;
            assign ap_AWQOS[73] = AP_AXIMM_73_AWQOS;
            assign ap_AWVALID[73] = AP_AXIMM_73_AWVALID;
            assign AP_AXIMM_73_AWREADY = ap_AWREADY[73];
            assign ap_WDATA[73][M_AXIMM_73_DATA_WIDTH-1:0] = AP_AXIMM_73_WDATA;
            assign ap_WSTRB[73][M_AXIMM_73_DATA_WIDTH/8-1:0] = AP_AXIMM_73_WSTRB;
            assign ap_WLAST[73] = AP_AXIMM_73_WLAST;
            assign ap_WVALID[73] = AP_AXIMM_73_WVALID;
            assign AP_AXIMM_73_WREADY = ap_WREADY[73];
            assign AP_AXIMM_73_BRESP = ap_BRESP[73];
            assign AP_AXIMM_73_BVALID = ap_BVALID[73];
            assign ap_BREADY[73] = AP_AXIMM_73_BREADY;
            assign ap_ARADDR[73][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_73_ARADDR;
            assign ap_ARLEN[73] = AP_AXIMM_73_ARLEN;
            assign ap_ARSIZE[73] = AP_AXIMM_73_ARSIZE;
            assign ap_ARBURST[73] = AP_AXIMM_73_ARBURST;
            assign ap_ARLOCK[73] = AP_AXIMM_73_ARLOCK;
            assign ap_ARCACHE[73] = AP_AXIMM_73_ARCACHE;
            assign ap_ARPROT[73] = AP_AXIMM_73_ARPROT;
            assign ap_ARREGION[73] = AP_AXIMM_73_ARREGION;
            assign ap_ARQOS[73] = AP_AXIMM_73_ARQOS;
            assign ap_ARVALID[73] = AP_AXIMM_73_ARVALID;
            assign AP_AXIMM_73_ARREADY = ap_ARREADY[73];
            assign AP_AXIMM_73_RDATA = ap_RDATA[73][M_AXIMM_73_DATA_WIDTH-1:0];
            assign AP_AXIMM_73_RRESP = ap_RRESP[73];
            assign AP_AXIMM_73_RLAST = ap_RLAST[73];
            assign AP_AXIMM_73_RVALID = ap_RVALID[73];
            assign ap_RREADY[73] = AP_AXIMM_73_RREADY;
            assign M_AXIMM_73_AWADDR = dm_AWADDR[73][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_73_AWLEN = dm_AWLEN[73];
            assign M_AXIMM_73_AWSIZE = dm_AWSIZE[73];
            assign M_AXIMM_73_AWBURST = dm_AWBURST[73];
            assign M_AXIMM_73_AWLOCK = dm_AWLOCK[73];
            assign M_AXIMM_73_AWCACHE = dm_AWCACHE[73];
            assign M_AXIMM_73_AWPROT = dm_AWPROT[73];
            assign M_AXIMM_73_AWREGION = dm_AWREGION[73];
            assign M_AXIMM_73_AWQOS = dm_AWQOS[73];
            assign M_AXIMM_73_AWVALID = dm_AWVALID[73];
            assign dm_AWREADY[73] = M_AXIMM_73_AWREADY;
            assign M_AXIMM_73_WDATA = dm_WDATA[73][M_AXIMM_73_DATA_WIDTH-1:0];
            assign M_AXIMM_73_WSTRB = dm_WSTRB[73][M_AXIMM_73_DATA_WIDTH/8-1:0];
            assign M_AXIMM_73_WLAST = dm_WLAST[73];
            assign M_AXIMM_73_WVALID = dm_WVALID[73];
            assign dm_WREADY[73] = M_AXIMM_73_WREADY;
            assign dm_BRESP[73] = M_AXIMM_73_BRESP;
            assign dm_BVALID[73] = M_AXIMM_73_BVALID;
            assign M_AXIMM_73_BREADY = dm_BREADY[73];
            assign M_AXIMM_73_ARADDR = dm_ARADDR[73][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_73_ARLEN = dm_ARLEN[73];
            assign M_AXIMM_73_ARSIZE = dm_ARSIZE[73];
            assign M_AXIMM_73_ARBURST = dm_ARBURST[73];
            assign M_AXIMM_73_ARLOCK = dm_ARLOCK[73];
            assign M_AXIMM_73_ARCACHE = dm_ARCACHE[73];
            assign M_AXIMM_73_ARPROT = dm_ARPROT[73];
            assign M_AXIMM_73_ARREGION = dm_ARREGION[73];
            assign M_AXIMM_73_ARQOS = dm_ARQOS[73];
            assign M_AXIMM_73_ARVALID = dm_ARVALID[73];
            assign dm_ARREADY[73] = M_AXIMM_73_ARREADY;
            assign dm_RDATA[73][M_AXIMM_73_DATA_WIDTH-1:0] = M_AXIMM_73_RDATA;
            assign dm_RRESP[73] = M_AXIMM_73_RRESP;
            assign dm_RLAST[73] = M_AXIMM_73_RLAST;
            assign dm_RVALID[73] = M_AXIMM_73_RVALID;
            assign M_AXIMM_73_RREADY = dm_RREADY[73];
        end
        if(C_NUM_AXIMMs > 74) begin
            assign ap_AWADDR[74][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_74_AWADDR;
            assign ap_AWLEN[74] = AP_AXIMM_74_AWLEN;
            assign ap_AWSIZE[74] = AP_AXIMM_74_AWSIZE;
            assign ap_AWBURST[74] = AP_AXIMM_74_AWBURST;
            assign ap_AWLOCK[74] = AP_AXIMM_74_AWLOCK;
            assign ap_AWCACHE[74] = AP_AXIMM_74_AWCACHE;
            assign ap_AWPROT[74] = AP_AXIMM_74_AWPROT;
            assign ap_AWREGION[74] = AP_AXIMM_74_AWREGION;
            assign ap_AWQOS[74] = AP_AXIMM_74_AWQOS;
            assign ap_AWVALID[74] = AP_AXIMM_74_AWVALID;
            assign AP_AXIMM_74_AWREADY = ap_AWREADY[74];
            assign ap_WDATA[74][M_AXIMM_74_DATA_WIDTH-1:0] = AP_AXIMM_74_WDATA;
            assign ap_WSTRB[74][M_AXIMM_74_DATA_WIDTH/8-1:0] = AP_AXIMM_74_WSTRB;
            assign ap_WLAST[74] = AP_AXIMM_74_WLAST;
            assign ap_WVALID[74] = AP_AXIMM_74_WVALID;
            assign AP_AXIMM_74_WREADY = ap_WREADY[74];
            assign AP_AXIMM_74_BRESP = ap_BRESP[74];
            assign AP_AXIMM_74_BVALID = ap_BVALID[74];
            assign ap_BREADY[74] = AP_AXIMM_74_BREADY;
            assign ap_ARADDR[74][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_74_ARADDR;
            assign ap_ARLEN[74] = AP_AXIMM_74_ARLEN;
            assign ap_ARSIZE[74] = AP_AXIMM_74_ARSIZE;
            assign ap_ARBURST[74] = AP_AXIMM_74_ARBURST;
            assign ap_ARLOCK[74] = AP_AXIMM_74_ARLOCK;
            assign ap_ARCACHE[74] = AP_AXIMM_74_ARCACHE;
            assign ap_ARPROT[74] = AP_AXIMM_74_ARPROT;
            assign ap_ARREGION[74] = AP_AXIMM_74_ARREGION;
            assign ap_ARQOS[74] = AP_AXIMM_74_ARQOS;
            assign ap_ARVALID[74] = AP_AXIMM_74_ARVALID;
            assign AP_AXIMM_74_ARREADY = ap_ARREADY[74];
            assign AP_AXIMM_74_RDATA = ap_RDATA[74][M_AXIMM_74_DATA_WIDTH-1:0];
            assign AP_AXIMM_74_RRESP = ap_RRESP[74];
            assign AP_AXIMM_74_RLAST = ap_RLAST[74];
            assign AP_AXIMM_74_RVALID = ap_RVALID[74];
            assign ap_RREADY[74] = AP_AXIMM_74_RREADY;
            assign M_AXIMM_74_AWADDR = dm_AWADDR[74][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_74_AWLEN = dm_AWLEN[74];
            assign M_AXIMM_74_AWSIZE = dm_AWSIZE[74];
            assign M_AXIMM_74_AWBURST = dm_AWBURST[74];
            assign M_AXIMM_74_AWLOCK = dm_AWLOCK[74];
            assign M_AXIMM_74_AWCACHE = dm_AWCACHE[74];
            assign M_AXIMM_74_AWPROT = dm_AWPROT[74];
            assign M_AXIMM_74_AWREGION = dm_AWREGION[74];
            assign M_AXIMM_74_AWQOS = dm_AWQOS[74];
            assign M_AXIMM_74_AWVALID = dm_AWVALID[74];
            assign dm_AWREADY[74] = M_AXIMM_74_AWREADY;
            assign M_AXIMM_74_WDATA = dm_WDATA[74][M_AXIMM_74_DATA_WIDTH-1:0];
            assign M_AXIMM_74_WSTRB = dm_WSTRB[74][M_AXIMM_74_DATA_WIDTH/8-1:0];
            assign M_AXIMM_74_WLAST = dm_WLAST[74];
            assign M_AXIMM_74_WVALID = dm_WVALID[74];
            assign dm_WREADY[74] = M_AXIMM_74_WREADY;
            assign dm_BRESP[74] = M_AXIMM_74_BRESP;
            assign dm_BVALID[74] = M_AXIMM_74_BVALID;
            assign M_AXIMM_74_BREADY = dm_BREADY[74];
            assign M_AXIMM_74_ARADDR = dm_ARADDR[74][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_74_ARLEN = dm_ARLEN[74];
            assign M_AXIMM_74_ARSIZE = dm_ARSIZE[74];
            assign M_AXIMM_74_ARBURST = dm_ARBURST[74];
            assign M_AXIMM_74_ARLOCK = dm_ARLOCK[74];
            assign M_AXIMM_74_ARCACHE = dm_ARCACHE[74];
            assign M_AXIMM_74_ARPROT = dm_ARPROT[74];
            assign M_AXIMM_74_ARREGION = dm_ARREGION[74];
            assign M_AXIMM_74_ARQOS = dm_ARQOS[74];
            assign M_AXIMM_74_ARVALID = dm_ARVALID[74];
            assign dm_ARREADY[74] = M_AXIMM_74_ARREADY;
            assign dm_RDATA[74][M_AXIMM_74_DATA_WIDTH-1:0] = M_AXIMM_74_RDATA;
            assign dm_RRESP[74] = M_AXIMM_74_RRESP;
            assign dm_RLAST[74] = M_AXIMM_74_RLAST;
            assign dm_RVALID[74] = M_AXIMM_74_RVALID;
            assign M_AXIMM_74_RREADY = dm_RREADY[74];
        end
        if(C_NUM_AXIMMs > 75) begin
            assign ap_AWADDR[75][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_75_AWADDR;
            assign ap_AWLEN[75] = AP_AXIMM_75_AWLEN;
            assign ap_AWSIZE[75] = AP_AXIMM_75_AWSIZE;
            assign ap_AWBURST[75] = AP_AXIMM_75_AWBURST;
            assign ap_AWLOCK[75] = AP_AXIMM_75_AWLOCK;
            assign ap_AWCACHE[75] = AP_AXIMM_75_AWCACHE;
            assign ap_AWPROT[75] = AP_AXIMM_75_AWPROT;
            assign ap_AWREGION[75] = AP_AXIMM_75_AWREGION;
            assign ap_AWQOS[75] = AP_AXIMM_75_AWQOS;
            assign ap_AWVALID[75] = AP_AXIMM_75_AWVALID;
            assign AP_AXIMM_75_AWREADY = ap_AWREADY[75];
            assign ap_WDATA[75][M_AXIMM_75_DATA_WIDTH-1:0] = AP_AXIMM_75_WDATA;
            assign ap_WSTRB[75][M_AXIMM_75_DATA_WIDTH/8-1:0] = AP_AXIMM_75_WSTRB;
            assign ap_WLAST[75] = AP_AXIMM_75_WLAST;
            assign ap_WVALID[75] = AP_AXIMM_75_WVALID;
            assign AP_AXIMM_75_WREADY = ap_WREADY[75];
            assign AP_AXIMM_75_BRESP = ap_BRESP[75];
            assign AP_AXIMM_75_BVALID = ap_BVALID[75];
            assign ap_BREADY[75] = AP_AXIMM_75_BREADY;
            assign ap_ARADDR[75][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_75_ARADDR;
            assign ap_ARLEN[75] = AP_AXIMM_75_ARLEN;
            assign ap_ARSIZE[75] = AP_AXIMM_75_ARSIZE;
            assign ap_ARBURST[75] = AP_AXIMM_75_ARBURST;
            assign ap_ARLOCK[75] = AP_AXIMM_75_ARLOCK;
            assign ap_ARCACHE[75] = AP_AXIMM_75_ARCACHE;
            assign ap_ARPROT[75] = AP_AXIMM_75_ARPROT;
            assign ap_ARREGION[75] = AP_AXIMM_75_ARREGION;
            assign ap_ARQOS[75] = AP_AXIMM_75_ARQOS;
            assign ap_ARVALID[75] = AP_AXIMM_75_ARVALID;
            assign AP_AXIMM_75_ARREADY = ap_ARREADY[75];
            assign AP_AXIMM_75_RDATA = ap_RDATA[75][M_AXIMM_75_DATA_WIDTH-1:0];
            assign AP_AXIMM_75_RRESP = ap_RRESP[75];
            assign AP_AXIMM_75_RLAST = ap_RLAST[75];
            assign AP_AXIMM_75_RVALID = ap_RVALID[75];
            assign ap_RREADY[75] = AP_AXIMM_75_RREADY;
            assign M_AXIMM_75_AWADDR = dm_AWADDR[75][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_75_AWLEN = dm_AWLEN[75];
            assign M_AXIMM_75_AWSIZE = dm_AWSIZE[75];
            assign M_AXIMM_75_AWBURST = dm_AWBURST[75];
            assign M_AXIMM_75_AWLOCK = dm_AWLOCK[75];
            assign M_AXIMM_75_AWCACHE = dm_AWCACHE[75];
            assign M_AXIMM_75_AWPROT = dm_AWPROT[75];
            assign M_AXIMM_75_AWREGION = dm_AWREGION[75];
            assign M_AXIMM_75_AWQOS = dm_AWQOS[75];
            assign M_AXIMM_75_AWVALID = dm_AWVALID[75];
            assign dm_AWREADY[75] = M_AXIMM_75_AWREADY;
            assign M_AXIMM_75_WDATA = dm_WDATA[75][M_AXIMM_75_DATA_WIDTH-1:0];
            assign M_AXIMM_75_WSTRB = dm_WSTRB[75][M_AXIMM_75_DATA_WIDTH/8-1:0];
            assign M_AXIMM_75_WLAST = dm_WLAST[75];
            assign M_AXIMM_75_WVALID = dm_WVALID[75];
            assign dm_WREADY[75] = M_AXIMM_75_WREADY;
            assign dm_BRESP[75] = M_AXIMM_75_BRESP;
            assign dm_BVALID[75] = M_AXIMM_75_BVALID;
            assign M_AXIMM_75_BREADY = dm_BREADY[75];
            assign M_AXIMM_75_ARADDR = dm_ARADDR[75][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_75_ARLEN = dm_ARLEN[75];
            assign M_AXIMM_75_ARSIZE = dm_ARSIZE[75];
            assign M_AXIMM_75_ARBURST = dm_ARBURST[75];
            assign M_AXIMM_75_ARLOCK = dm_ARLOCK[75];
            assign M_AXIMM_75_ARCACHE = dm_ARCACHE[75];
            assign M_AXIMM_75_ARPROT = dm_ARPROT[75];
            assign M_AXIMM_75_ARREGION = dm_ARREGION[75];
            assign M_AXIMM_75_ARQOS = dm_ARQOS[75];
            assign M_AXIMM_75_ARVALID = dm_ARVALID[75];
            assign dm_ARREADY[75] = M_AXIMM_75_ARREADY;
            assign dm_RDATA[75][M_AXIMM_75_DATA_WIDTH-1:0] = M_AXIMM_75_RDATA;
            assign dm_RRESP[75] = M_AXIMM_75_RRESP;
            assign dm_RLAST[75] = M_AXIMM_75_RLAST;
            assign dm_RVALID[75] = M_AXIMM_75_RVALID;
            assign M_AXIMM_75_RREADY = dm_RREADY[75];
        end
        if(C_NUM_AXIMMs > 76) begin
            assign ap_AWADDR[76][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_76_AWADDR;
            assign ap_AWLEN[76] = AP_AXIMM_76_AWLEN;
            assign ap_AWSIZE[76] = AP_AXIMM_76_AWSIZE;
            assign ap_AWBURST[76] = AP_AXIMM_76_AWBURST;
            assign ap_AWLOCK[76] = AP_AXIMM_76_AWLOCK;
            assign ap_AWCACHE[76] = AP_AXIMM_76_AWCACHE;
            assign ap_AWPROT[76] = AP_AXIMM_76_AWPROT;
            assign ap_AWREGION[76] = AP_AXIMM_76_AWREGION;
            assign ap_AWQOS[76] = AP_AXIMM_76_AWQOS;
            assign ap_AWVALID[76] = AP_AXIMM_76_AWVALID;
            assign AP_AXIMM_76_AWREADY = ap_AWREADY[76];
            assign ap_WDATA[76][M_AXIMM_76_DATA_WIDTH-1:0] = AP_AXIMM_76_WDATA;
            assign ap_WSTRB[76][M_AXIMM_76_DATA_WIDTH/8-1:0] = AP_AXIMM_76_WSTRB;
            assign ap_WLAST[76] = AP_AXIMM_76_WLAST;
            assign ap_WVALID[76] = AP_AXIMM_76_WVALID;
            assign AP_AXIMM_76_WREADY = ap_WREADY[76];
            assign AP_AXIMM_76_BRESP = ap_BRESP[76];
            assign AP_AXIMM_76_BVALID = ap_BVALID[76];
            assign ap_BREADY[76] = AP_AXIMM_76_BREADY;
            assign ap_ARADDR[76][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_76_ARADDR;
            assign ap_ARLEN[76] = AP_AXIMM_76_ARLEN;
            assign ap_ARSIZE[76] = AP_AXIMM_76_ARSIZE;
            assign ap_ARBURST[76] = AP_AXIMM_76_ARBURST;
            assign ap_ARLOCK[76] = AP_AXIMM_76_ARLOCK;
            assign ap_ARCACHE[76] = AP_AXIMM_76_ARCACHE;
            assign ap_ARPROT[76] = AP_AXIMM_76_ARPROT;
            assign ap_ARREGION[76] = AP_AXIMM_76_ARREGION;
            assign ap_ARQOS[76] = AP_AXIMM_76_ARQOS;
            assign ap_ARVALID[76] = AP_AXIMM_76_ARVALID;
            assign AP_AXIMM_76_ARREADY = ap_ARREADY[76];
            assign AP_AXIMM_76_RDATA = ap_RDATA[76][M_AXIMM_76_DATA_WIDTH-1:0];
            assign AP_AXIMM_76_RRESP = ap_RRESP[76];
            assign AP_AXIMM_76_RLAST = ap_RLAST[76];
            assign AP_AXIMM_76_RVALID = ap_RVALID[76];
            assign ap_RREADY[76] = AP_AXIMM_76_RREADY;
            assign M_AXIMM_76_AWADDR = dm_AWADDR[76][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_76_AWLEN = dm_AWLEN[76];
            assign M_AXIMM_76_AWSIZE = dm_AWSIZE[76];
            assign M_AXIMM_76_AWBURST = dm_AWBURST[76];
            assign M_AXIMM_76_AWLOCK = dm_AWLOCK[76];
            assign M_AXIMM_76_AWCACHE = dm_AWCACHE[76];
            assign M_AXIMM_76_AWPROT = dm_AWPROT[76];
            assign M_AXIMM_76_AWREGION = dm_AWREGION[76];
            assign M_AXIMM_76_AWQOS = dm_AWQOS[76];
            assign M_AXIMM_76_AWVALID = dm_AWVALID[76];
            assign dm_AWREADY[76] = M_AXIMM_76_AWREADY;
            assign M_AXIMM_76_WDATA = dm_WDATA[76][M_AXIMM_76_DATA_WIDTH-1:0];
            assign M_AXIMM_76_WSTRB = dm_WSTRB[76][M_AXIMM_76_DATA_WIDTH/8-1:0];
            assign M_AXIMM_76_WLAST = dm_WLAST[76];
            assign M_AXIMM_76_WVALID = dm_WVALID[76];
            assign dm_WREADY[76] = M_AXIMM_76_WREADY;
            assign dm_BRESP[76] = M_AXIMM_76_BRESP;
            assign dm_BVALID[76] = M_AXIMM_76_BVALID;
            assign M_AXIMM_76_BREADY = dm_BREADY[76];
            assign M_AXIMM_76_ARADDR = dm_ARADDR[76][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_76_ARLEN = dm_ARLEN[76];
            assign M_AXIMM_76_ARSIZE = dm_ARSIZE[76];
            assign M_AXIMM_76_ARBURST = dm_ARBURST[76];
            assign M_AXIMM_76_ARLOCK = dm_ARLOCK[76];
            assign M_AXIMM_76_ARCACHE = dm_ARCACHE[76];
            assign M_AXIMM_76_ARPROT = dm_ARPROT[76];
            assign M_AXIMM_76_ARREGION = dm_ARREGION[76];
            assign M_AXIMM_76_ARQOS = dm_ARQOS[76];
            assign M_AXIMM_76_ARVALID = dm_ARVALID[76];
            assign dm_ARREADY[76] = M_AXIMM_76_ARREADY;
            assign dm_RDATA[76][M_AXIMM_76_DATA_WIDTH-1:0] = M_AXIMM_76_RDATA;
            assign dm_RRESP[76] = M_AXIMM_76_RRESP;
            assign dm_RLAST[76] = M_AXIMM_76_RLAST;
            assign dm_RVALID[76] = M_AXIMM_76_RVALID;
            assign M_AXIMM_76_RREADY = dm_RREADY[76];
        end
        if(C_NUM_AXIMMs > 77) begin
            assign ap_AWADDR[77][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_77_AWADDR;
            assign ap_AWLEN[77] = AP_AXIMM_77_AWLEN;
            assign ap_AWSIZE[77] = AP_AXIMM_77_AWSIZE;
            assign ap_AWBURST[77] = AP_AXIMM_77_AWBURST;
            assign ap_AWLOCK[77] = AP_AXIMM_77_AWLOCK;
            assign ap_AWCACHE[77] = AP_AXIMM_77_AWCACHE;
            assign ap_AWPROT[77] = AP_AXIMM_77_AWPROT;
            assign ap_AWREGION[77] = AP_AXIMM_77_AWREGION;
            assign ap_AWQOS[77] = AP_AXIMM_77_AWQOS;
            assign ap_AWVALID[77] = AP_AXIMM_77_AWVALID;
            assign AP_AXIMM_77_AWREADY = ap_AWREADY[77];
            assign ap_WDATA[77][M_AXIMM_77_DATA_WIDTH-1:0] = AP_AXIMM_77_WDATA;
            assign ap_WSTRB[77][M_AXIMM_77_DATA_WIDTH/8-1:0] = AP_AXIMM_77_WSTRB;
            assign ap_WLAST[77] = AP_AXIMM_77_WLAST;
            assign ap_WVALID[77] = AP_AXIMM_77_WVALID;
            assign AP_AXIMM_77_WREADY = ap_WREADY[77];
            assign AP_AXIMM_77_BRESP = ap_BRESP[77];
            assign AP_AXIMM_77_BVALID = ap_BVALID[77];
            assign ap_BREADY[77] = AP_AXIMM_77_BREADY;
            assign ap_ARADDR[77][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_77_ARADDR;
            assign ap_ARLEN[77] = AP_AXIMM_77_ARLEN;
            assign ap_ARSIZE[77] = AP_AXIMM_77_ARSIZE;
            assign ap_ARBURST[77] = AP_AXIMM_77_ARBURST;
            assign ap_ARLOCK[77] = AP_AXIMM_77_ARLOCK;
            assign ap_ARCACHE[77] = AP_AXIMM_77_ARCACHE;
            assign ap_ARPROT[77] = AP_AXIMM_77_ARPROT;
            assign ap_ARREGION[77] = AP_AXIMM_77_ARREGION;
            assign ap_ARQOS[77] = AP_AXIMM_77_ARQOS;
            assign ap_ARVALID[77] = AP_AXIMM_77_ARVALID;
            assign AP_AXIMM_77_ARREADY = ap_ARREADY[77];
            assign AP_AXIMM_77_RDATA = ap_RDATA[77][M_AXIMM_77_DATA_WIDTH-1:0];
            assign AP_AXIMM_77_RRESP = ap_RRESP[77];
            assign AP_AXIMM_77_RLAST = ap_RLAST[77];
            assign AP_AXIMM_77_RVALID = ap_RVALID[77];
            assign ap_RREADY[77] = AP_AXIMM_77_RREADY;
            assign M_AXIMM_77_AWADDR = dm_AWADDR[77][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_77_AWLEN = dm_AWLEN[77];
            assign M_AXIMM_77_AWSIZE = dm_AWSIZE[77];
            assign M_AXIMM_77_AWBURST = dm_AWBURST[77];
            assign M_AXIMM_77_AWLOCK = dm_AWLOCK[77];
            assign M_AXIMM_77_AWCACHE = dm_AWCACHE[77];
            assign M_AXIMM_77_AWPROT = dm_AWPROT[77];
            assign M_AXIMM_77_AWREGION = dm_AWREGION[77];
            assign M_AXIMM_77_AWQOS = dm_AWQOS[77];
            assign M_AXIMM_77_AWVALID = dm_AWVALID[77];
            assign dm_AWREADY[77] = M_AXIMM_77_AWREADY;
            assign M_AXIMM_77_WDATA = dm_WDATA[77][M_AXIMM_77_DATA_WIDTH-1:0];
            assign M_AXIMM_77_WSTRB = dm_WSTRB[77][M_AXIMM_77_DATA_WIDTH/8-1:0];
            assign M_AXIMM_77_WLAST = dm_WLAST[77];
            assign M_AXIMM_77_WVALID = dm_WVALID[77];
            assign dm_WREADY[77] = M_AXIMM_77_WREADY;
            assign dm_BRESP[77] = M_AXIMM_77_BRESP;
            assign dm_BVALID[77] = M_AXIMM_77_BVALID;
            assign M_AXIMM_77_BREADY = dm_BREADY[77];
            assign M_AXIMM_77_ARADDR = dm_ARADDR[77][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_77_ARLEN = dm_ARLEN[77];
            assign M_AXIMM_77_ARSIZE = dm_ARSIZE[77];
            assign M_AXIMM_77_ARBURST = dm_ARBURST[77];
            assign M_AXIMM_77_ARLOCK = dm_ARLOCK[77];
            assign M_AXIMM_77_ARCACHE = dm_ARCACHE[77];
            assign M_AXIMM_77_ARPROT = dm_ARPROT[77];
            assign M_AXIMM_77_ARREGION = dm_ARREGION[77];
            assign M_AXIMM_77_ARQOS = dm_ARQOS[77];
            assign M_AXIMM_77_ARVALID = dm_ARVALID[77];
            assign dm_ARREADY[77] = M_AXIMM_77_ARREADY;
            assign dm_RDATA[77][M_AXIMM_77_DATA_WIDTH-1:0] = M_AXIMM_77_RDATA;
            assign dm_RRESP[77] = M_AXIMM_77_RRESP;
            assign dm_RLAST[77] = M_AXIMM_77_RLAST;
            assign dm_RVALID[77] = M_AXIMM_77_RVALID;
            assign M_AXIMM_77_RREADY = dm_RREADY[77];
        end
        if(C_NUM_AXIMMs > 78) begin
            assign ap_AWADDR[78][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_78_AWADDR;
            assign ap_AWLEN[78] = AP_AXIMM_78_AWLEN;
            assign ap_AWSIZE[78] = AP_AXIMM_78_AWSIZE;
            assign ap_AWBURST[78] = AP_AXIMM_78_AWBURST;
            assign ap_AWLOCK[78] = AP_AXIMM_78_AWLOCK;
            assign ap_AWCACHE[78] = AP_AXIMM_78_AWCACHE;
            assign ap_AWPROT[78] = AP_AXIMM_78_AWPROT;
            assign ap_AWREGION[78] = AP_AXIMM_78_AWREGION;
            assign ap_AWQOS[78] = AP_AXIMM_78_AWQOS;
            assign ap_AWVALID[78] = AP_AXIMM_78_AWVALID;
            assign AP_AXIMM_78_AWREADY = ap_AWREADY[78];
            assign ap_WDATA[78][M_AXIMM_78_DATA_WIDTH-1:0] = AP_AXIMM_78_WDATA;
            assign ap_WSTRB[78][M_AXIMM_78_DATA_WIDTH/8-1:0] = AP_AXIMM_78_WSTRB;
            assign ap_WLAST[78] = AP_AXIMM_78_WLAST;
            assign ap_WVALID[78] = AP_AXIMM_78_WVALID;
            assign AP_AXIMM_78_WREADY = ap_WREADY[78];
            assign AP_AXIMM_78_BRESP = ap_BRESP[78];
            assign AP_AXIMM_78_BVALID = ap_BVALID[78];
            assign ap_BREADY[78] = AP_AXIMM_78_BREADY;
            assign ap_ARADDR[78][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_78_ARADDR;
            assign ap_ARLEN[78] = AP_AXIMM_78_ARLEN;
            assign ap_ARSIZE[78] = AP_AXIMM_78_ARSIZE;
            assign ap_ARBURST[78] = AP_AXIMM_78_ARBURST;
            assign ap_ARLOCK[78] = AP_AXIMM_78_ARLOCK;
            assign ap_ARCACHE[78] = AP_AXIMM_78_ARCACHE;
            assign ap_ARPROT[78] = AP_AXIMM_78_ARPROT;
            assign ap_ARREGION[78] = AP_AXIMM_78_ARREGION;
            assign ap_ARQOS[78] = AP_AXIMM_78_ARQOS;
            assign ap_ARVALID[78] = AP_AXIMM_78_ARVALID;
            assign AP_AXIMM_78_ARREADY = ap_ARREADY[78];
            assign AP_AXIMM_78_RDATA = ap_RDATA[78][M_AXIMM_78_DATA_WIDTH-1:0];
            assign AP_AXIMM_78_RRESP = ap_RRESP[78];
            assign AP_AXIMM_78_RLAST = ap_RLAST[78];
            assign AP_AXIMM_78_RVALID = ap_RVALID[78];
            assign ap_RREADY[78] = AP_AXIMM_78_RREADY;
            assign M_AXIMM_78_AWADDR = dm_AWADDR[78][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_78_AWLEN = dm_AWLEN[78];
            assign M_AXIMM_78_AWSIZE = dm_AWSIZE[78];
            assign M_AXIMM_78_AWBURST = dm_AWBURST[78];
            assign M_AXIMM_78_AWLOCK = dm_AWLOCK[78];
            assign M_AXIMM_78_AWCACHE = dm_AWCACHE[78];
            assign M_AXIMM_78_AWPROT = dm_AWPROT[78];
            assign M_AXIMM_78_AWREGION = dm_AWREGION[78];
            assign M_AXIMM_78_AWQOS = dm_AWQOS[78];
            assign M_AXIMM_78_AWVALID = dm_AWVALID[78];
            assign dm_AWREADY[78] = M_AXIMM_78_AWREADY;
            assign M_AXIMM_78_WDATA = dm_WDATA[78][M_AXIMM_78_DATA_WIDTH-1:0];
            assign M_AXIMM_78_WSTRB = dm_WSTRB[78][M_AXIMM_78_DATA_WIDTH/8-1:0];
            assign M_AXIMM_78_WLAST = dm_WLAST[78];
            assign M_AXIMM_78_WVALID = dm_WVALID[78];
            assign dm_WREADY[78] = M_AXIMM_78_WREADY;
            assign dm_BRESP[78] = M_AXIMM_78_BRESP;
            assign dm_BVALID[78] = M_AXIMM_78_BVALID;
            assign M_AXIMM_78_BREADY = dm_BREADY[78];
            assign M_AXIMM_78_ARADDR = dm_ARADDR[78][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_78_ARLEN = dm_ARLEN[78];
            assign M_AXIMM_78_ARSIZE = dm_ARSIZE[78];
            assign M_AXIMM_78_ARBURST = dm_ARBURST[78];
            assign M_AXIMM_78_ARLOCK = dm_ARLOCK[78];
            assign M_AXIMM_78_ARCACHE = dm_ARCACHE[78];
            assign M_AXIMM_78_ARPROT = dm_ARPROT[78];
            assign M_AXIMM_78_ARREGION = dm_ARREGION[78];
            assign M_AXIMM_78_ARQOS = dm_ARQOS[78];
            assign M_AXIMM_78_ARVALID = dm_ARVALID[78];
            assign dm_ARREADY[78] = M_AXIMM_78_ARREADY;
            assign dm_RDATA[78][M_AXIMM_78_DATA_WIDTH-1:0] = M_AXIMM_78_RDATA;
            assign dm_RRESP[78] = M_AXIMM_78_RRESP;
            assign dm_RLAST[78] = M_AXIMM_78_RLAST;
            assign dm_RVALID[78] = M_AXIMM_78_RVALID;
            assign M_AXIMM_78_RREADY = dm_RREADY[78];
        end
        if(C_NUM_AXIMMs > 79) begin
            assign ap_AWADDR[79][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_79_AWADDR;
            assign ap_AWLEN[79] = AP_AXIMM_79_AWLEN;
            assign ap_AWSIZE[79] = AP_AXIMM_79_AWSIZE;
            assign ap_AWBURST[79] = AP_AXIMM_79_AWBURST;
            assign ap_AWLOCK[79] = AP_AXIMM_79_AWLOCK;
            assign ap_AWCACHE[79] = AP_AXIMM_79_AWCACHE;
            assign ap_AWPROT[79] = AP_AXIMM_79_AWPROT;
            assign ap_AWREGION[79] = AP_AXIMM_79_AWREGION;
            assign ap_AWQOS[79] = AP_AXIMM_79_AWQOS;
            assign ap_AWVALID[79] = AP_AXIMM_79_AWVALID;
            assign AP_AXIMM_79_AWREADY = ap_AWREADY[79];
            assign ap_WDATA[79][M_AXIMM_79_DATA_WIDTH-1:0] = AP_AXIMM_79_WDATA;
            assign ap_WSTRB[79][M_AXIMM_79_DATA_WIDTH/8-1:0] = AP_AXIMM_79_WSTRB;
            assign ap_WLAST[79] = AP_AXIMM_79_WLAST;
            assign ap_WVALID[79] = AP_AXIMM_79_WVALID;
            assign AP_AXIMM_79_WREADY = ap_WREADY[79];
            assign AP_AXIMM_79_BRESP = ap_BRESP[79];
            assign AP_AXIMM_79_BVALID = ap_BVALID[79];
            assign ap_BREADY[79] = AP_AXIMM_79_BREADY;
            assign ap_ARADDR[79][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_79_ARADDR;
            assign ap_ARLEN[79] = AP_AXIMM_79_ARLEN;
            assign ap_ARSIZE[79] = AP_AXIMM_79_ARSIZE;
            assign ap_ARBURST[79] = AP_AXIMM_79_ARBURST;
            assign ap_ARLOCK[79] = AP_AXIMM_79_ARLOCK;
            assign ap_ARCACHE[79] = AP_AXIMM_79_ARCACHE;
            assign ap_ARPROT[79] = AP_AXIMM_79_ARPROT;
            assign ap_ARREGION[79] = AP_AXIMM_79_ARREGION;
            assign ap_ARQOS[79] = AP_AXIMM_79_ARQOS;
            assign ap_ARVALID[79] = AP_AXIMM_79_ARVALID;
            assign AP_AXIMM_79_ARREADY = ap_ARREADY[79];
            assign AP_AXIMM_79_RDATA = ap_RDATA[79][M_AXIMM_79_DATA_WIDTH-1:0];
            assign AP_AXIMM_79_RRESP = ap_RRESP[79];
            assign AP_AXIMM_79_RLAST = ap_RLAST[79];
            assign AP_AXIMM_79_RVALID = ap_RVALID[79];
            assign ap_RREADY[79] = AP_AXIMM_79_RREADY;
            assign M_AXIMM_79_AWADDR = dm_AWADDR[79][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_79_AWLEN = dm_AWLEN[79];
            assign M_AXIMM_79_AWSIZE = dm_AWSIZE[79];
            assign M_AXIMM_79_AWBURST = dm_AWBURST[79];
            assign M_AXIMM_79_AWLOCK = dm_AWLOCK[79];
            assign M_AXIMM_79_AWCACHE = dm_AWCACHE[79];
            assign M_AXIMM_79_AWPROT = dm_AWPROT[79];
            assign M_AXIMM_79_AWREGION = dm_AWREGION[79];
            assign M_AXIMM_79_AWQOS = dm_AWQOS[79];
            assign M_AXIMM_79_AWVALID = dm_AWVALID[79];
            assign dm_AWREADY[79] = M_AXIMM_79_AWREADY;
            assign M_AXIMM_79_WDATA = dm_WDATA[79][M_AXIMM_79_DATA_WIDTH-1:0];
            assign M_AXIMM_79_WSTRB = dm_WSTRB[79][M_AXIMM_79_DATA_WIDTH/8-1:0];
            assign M_AXIMM_79_WLAST = dm_WLAST[79];
            assign M_AXIMM_79_WVALID = dm_WVALID[79];
            assign dm_WREADY[79] = M_AXIMM_79_WREADY;
            assign dm_BRESP[79] = M_AXIMM_79_BRESP;
            assign dm_BVALID[79] = M_AXIMM_79_BVALID;
            assign M_AXIMM_79_BREADY = dm_BREADY[79];
            assign M_AXIMM_79_ARADDR = dm_ARADDR[79][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_79_ARLEN = dm_ARLEN[79];
            assign M_AXIMM_79_ARSIZE = dm_ARSIZE[79];
            assign M_AXIMM_79_ARBURST = dm_ARBURST[79];
            assign M_AXIMM_79_ARLOCK = dm_ARLOCK[79];
            assign M_AXIMM_79_ARCACHE = dm_ARCACHE[79];
            assign M_AXIMM_79_ARPROT = dm_ARPROT[79];
            assign M_AXIMM_79_ARREGION = dm_ARREGION[79];
            assign M_AXIMM_79_ARQOS = dm_ARQOS[79];
            assign M_AXIMM_79_ARVALID = dm_ARVALID[79];
            assign dm_ARREADY[79] = M_AXIMM_79_ARREADY;
            assign dm_RDATA[79][M_AXIMM_79_DATA_WIDTH-1:0] = M_AXIMM_79_RDATA;
            assign dm_RRESP[79] = M_AXIMM_79_RRESP;
            assign dm_RLAST[79] = M_AXIMM_79_RLAST;
            assign dm_RVALID[79] = M_AXIMM_79_RVALID;
            assign M_AXIMM_79_RREADY = dm_RREADY[79];
        end
        if(C_NUM_AXIMMs > 80) begin
            assign ap_AWADDR[80][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_80_AWADDR;
            assign ap_AWLEN[80] = AP_AXIMM_80_AWLEN;
            assign ap_AWSIZE[80] = AP_AXIMM_80_AWSIZE;
            assign ap_AWBURST[80] = AP_AXIMM_80_AWBURST;
            assign ap_AWLOCK[80] = AP_AXIMM_80_AWLOCK;
            assign ap_AWCACHE[80] = AP_AXIMM_80_AWCACHE;
            assign ap_AWPROT[80] = AP_AXIMM_80_AWPROT;
            assign ap_AWREGION[80] = AP_AXIMM_80_AWREGION;
            assign ap_AWQOS[80] = AP_AXIMM_80_AWQOS;
            assign ap_AWVALID[80] = AP_AXIMM_80_AWVALID;
            assign AP_AXIMM_80_AWREADY = ap_AWREADY[80];
            assign ap_WDATA[80][M_AXIMM_80_DATA_WIDTH-1:0] = AP_AXIMM_80_WDATA;
            assign ap_WSTRB[80][M_AXIMM_80_DATA_WIDTH/8-1:0] = AP_AXIMM_80_WSTRB;
            assign ap_WLAST[80] = AP_AXIMM_80_WLAST;
            assign ap_WVALID[80] = AP_AXIMM_80_WVALID;
            assign AP_AXIMM_80_WREADY = ap_WREADY[80];
            assign AP_AXIMM_80_BRESP = ap_BRESP[80];
            assign AP_AXIMM_80_BVALID = ap_BVALID[80];
            assign ap_BREADY[80] = AP_AXIMM_80_BREADY;
            assign ap_ARADDR[80][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_80_ARADDR;
            assign ap_ARLEN[80] = AP_AXIMM_80_ARLEN;
            assign ap_ARSIZE[80] = AP_AXIMM_80_ARSIZE;
            assign ap_ARBURST[80] = AP_AXIMM_80_ARBURST;
            assign ap_ARLOCK[80] = AP_AXIMM_80_ARLOCK;
            assign ap_ARCACHE[80] = AP_AXIMM_80_ARCACHE;
            assign ap_ARPROT[80] = AP_AXIMM_80_ARPROT;
            assign ap_ARREGION[80] = AP_AXIMM_80_ARREGION;
            assign ap_ARQOS[80] = AP_AXIMM_80_ARQOS;
            assign ap_ARVALID[80] = AP_AXIMM_80_ARVALID;
            assign AP_AXIMM_80_ARREADY = ap_ARREADY[80];
            assign AP_AXIMM_80_RDATA = ap_RDATA[80][M_AXIMM_80_DATA_WIDTH-1:0];
            assign AP_AXIMM_80_RRESP = ap_RRESP[80];
            assign AP_AXIMM_80_RLAST = ap_RLAST[80];
            assign AP_AXIMM_80_RVALID = ap_RVALID[80];
            assign ap_RREADY[80] = AP_AXIMM_80_RREADY;
            assign M_AXIMM_80_AWADDR = dm_AWADDR[80][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_80_AWLEN = dm_AWLEN[80];
            assign M_AXIMM_80_AWSIZE = dm_AWSIZE[80];
            assign M_AXIMM_80_AWBURST = dm_AWBURST[80];
            assign M_AXIMM_80_AWLOCK = dm_AWLOCK[80];
            assign M_AXIMM_80_AWCACHE = dm_AWCACHE[80];
            assign M_AXIMM_80_AWPROT = dm_AWPROT[80];
            assign M_AXIMM_80_AWREGION = dm_AWREGION[80];
            assign M_AXIMM_80_AWQOS = dm_AWQOS[80];
            assign M_AXIMM_80_AWVALID = dm_AWVALID[80];
            assign dm_AWREADY[80] = M_AXIMM_80_AWREADY;
            assign M_AXIMM_80_WDATA = dm_WDATA[80][M_AXIMM_80_DATA_WIDTH-1:0];
            assign M_AXIMM_80_WSTRB = dm_WSTRB[80][M_AXIMM_80_DATA_WIDTH/8-1:0];
            assign M_AXIMM_80_WLAST = dm_WLAST[80];
            assign M_AXIMM_80_WVALID = dm_WVALID[80];
            assign dm_WREADY[80] = M_AXIMM_80_WREADY;
            assign dm_BRESP[80] = M_AXIMM_80_BRESP;
            assign dm_BVALID[80] = M_AXIMM_80_BVALID;
            assign M_AXIMM_80_BREADY = dm_BREADY[80];
            assign M_AXIMM_80_ARADDR = dm_ARADDR[80][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_80_ARLEN = dm_ARLEN[80];
            assign M_AXIMM_80_ARSIZE = dm_ARSIZE[80];
            assign M_AXIMM_80_ARBURST = dm_ARBURST[80];
            assign M_AXIMM_80_ARLOCK = dm_ARLOCK[80];
            assign M_AXIMM_80_ARCACHE = dm_ARCACHE[80];
            assign M_AXIMM_80_ARPROT = dm_ARPROT[80];
            assign M_AXIMM_80_ARREGION = dm_ARREGION[80];
            assign M_AXIMM_80_ARQOS = dm_ARQOS[80];
            assign M_AXIMM_80_ARVALID = dm_ARVALID[80];
            assign dm_ARREADY[80] = M_AXIMM_80_ARREADY;
            assign dm_RDATA[80][M_AXIMM_80_DATA_WIDTH-1:0] = M_AXIMM_80_RDATA;
            assign dm_RRESP[80] = M_AXIMM_80_RRESP;
            assign dm_RLAST[80] = M_AXIMM_80_RLAST;
            assign dm_RVALID[80] = M_AXIMM_80_RVALID;
            assign M_AXIMM_80_RREADY = dm_RREADY[80];
        end
        if(C_NUM_AXIMMs > 81) begin
            assign ap_AWADDR[81][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_81_AWADDR;
            assign ap_AWLEN[81] = AP_AXIMM_81_AWLEN;
            assign ap_AWSIZE[81] = AP_AXIMM_81_AWSIZE;
            assign ap_AWBURST[81] = AP_AXIMM_81_AWBURST;
            assign ap_AWLOCK[81] = AP_AXIMM_81_AWLOCK;
            assign ap_AWCACHE[81] = AP_AXIMM_81_AWCACHE;
            assign ap_AWPROT[81] = AP_AXIMM_81_AWPROT;
            assign ap_AWREGION[81] = AP_AXIMM_81_AWREGION;
            assign ap_AWQOS[81] = AP_AXIMM_81_AWQOS;
            assign ap_AWVALID[81] = AP_AXIMM_81_AWVALID;
            assign AP_AXIMM_81_AWREADY = ap_AWREADY[81];
            assign ap_WDATA[81][M_AXIMM_81_DATA_WIDTH-1:0] = AP_AXIMM_81_WDATA;
            assign ap_WSTRB[81][M_AXIMM_81_DATA_WIDTH/8-1:0] = AP_AXIMM_81_WSTRB;
            assign ap_WLAST[81] = AP_AXIMM_81_WLAST;
            assign ap_WVALID[81] = AP_AXIMM_81_WVALID;
            assign AP_AXIMM_81_WREADY = ap_WREADY[81];
            assign AP_AXIMM_81_BRESP = ap_BRESP[81];
            assign AP_AXIMM_81_BVALID = ap_BVALID[81];
            assign ap_BREADY[81] = AP_AXIMM_81_BREADY;
            assign ap_ARADDR[81][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_81_ARADDR;
            assign ap_ARLEN[81] = AP_AXIMM_81_ARLEN;
            assign ap_ARSIZE[81] = AP_AXIMM_81_ARSIZE;
            assign ap_ARBURST[81] = AP_AXIMM_81_ARBURST;
            assign ap_ARLOCK[81] = AP_AXIMM_81_ARLOCK;
            assign ap_ARCACHE[81] = AP_AXIMM_81_ARCACHE;
            assign ap_ARPROT[81] = AP_AXIMM_81_ARPROT;
            assign ap_ARREGION[81] = AP_AXIMM_81_ARREGION;
            assign ap_ARQOS[81] = AP_AXIMM_81_ARQOS;
            assign ap_ARVALID[81] = AP_AXIMM_81_ARVALID;
            assign AP_AXIMM_81_ARREADY = ap_ARREADY[81];
            assign AP_AXIMM_81_RDATA = ap_RDATA[81][M_AXIMM_81_DATA_WIDTH-1:0];
            assign AP_AXIMM_81_RRESP = ap_RRESP[81];
            assign AP_AXIMM_81_RLAST = ap_RLAST[81];
            assign AP_AXIMM_81_RVALID = ap_RVALID[81];
            assign ap_RREADY[81] = AP_AXIMM_81_RREADY;
            assign M_AXIMM_81_AWADDR = dm_AWADDR[81][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_81_AWLEN = dm_AWLEN[81];
            assign M_AXIMM_81_AWSIZE = dm_AWSIZE[81];
            assign M_AXIMM_81_AWBURST = dm_AWBURST[81];
            assign M_AXIMM_81_AWLOCK = dm_AWLOCK[81];
            assign M_AXIMM_81_AWCACHE = dm_AWCACHE[81];
            assign M_AXIMM_81_AWPROT = dm_AWPROT[81];
            assign M_AXIMM_81_AWREGION = dm_AWREGION[81];
            assign M_AXIMM_81_AWQOS = dm_AWQOS[81];
            assign M_AXIMM_81_AWVALID = dm_AWVALID[81];
            assign dm_AWREADY[81] = M_AXIMM_81_AWREADY;
            assign M_AXIMM_81_WDATA = dm_WDATA[81][M_AXIMM_81_DATA_WIDTH-1:0];
            assign M_AXIMM_81_WSTRB = dm_WSTRB[81][M_AXIMM_81_DATA_WIDTH/8-1:0];
            assign M_AXIMM_81_WLAST = dm_WLAST[81];
            assign M_AXIMM_81_WVALID = dm_WVALID[81];
            assign dm_WREADY[81] = M_AXIMM_81_WREADY;
            assign dm_BRESP[81] = M_AXIMM_81_BRESP;
            assign dm_BVALID[81] = M_AXIMM_81_BVALID;
            assign M_AXIMM_81_BREADY = dm_BREADY[81];
            assign M_AXIMM_81_ARADDR = dm_ARADDR[81][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_81_ARLEN = dm_ARLEN[81];
            assign M_AXIMM_81_ARSIZE = dm_ARSIZE[81];
            assign M_AXIMM_81_ARBURST = dm_ARBURST[81];
            assign M_AXIMM_81_ARLOCK = dm_ARLOCK[81];
            assign M_AXIMM_81_ARCACHE = dm_ARCACHE[81];
            assign M_AXIMM_81_ARPROT = dm_ARPROT[81];
            assign M_AXIMM_81_ARREGION = dm_ARREGION[81];
            assign M_AXIMM_81_ARQOS = dm_ARQOS[81];
            assign M_AXIMM_81_ARVALID = dm_ARVALID[81];
            assign dm_ARREADY[81] = M_AXIMM_81_ARREADY;
            assign dm_RDATA[81][M_AXIMM_81_DATA_WIDTH-1:0] = M_AXIMM_81_RDATA;
            assign dm_RRESP[81] = M_AXIMM_81_RRESP;
            assign dm_RLAST[81] = M_AXIMM_81_RLAST;
            assign dm_RVALID[81] = M_AXIMM_81_RVALID;
            assign M_AXIMM_81_RREADY = dm_RREADY[81];
        end
        if(C_NUM_AXIMMs > 82) begin
            assign ap_AWADDR[82][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_82_AWADDR;
            assign ap_AWLEN[82] = AP_AXIMM_82_AWLEN;
            assign ap_AWSIZE[82] = AP_AXIMM_82_AWSIZE;
            assign ap_AWBURST[82] = AP_AXIMM_82_AWBURST;
            assign ap_AWLOCK[82] = AP_AXIMM_82_AWLOCK;
            assign ap_AWCACHE[82] = AP_AXIMM_82_AWCACHE;
            assign ap_AWPROT[82] = AP_AXIMM_82_AWPROT;
            assign ap_AWREGION[82] = AP_AXIMM_82_AWREGION;
            assign ap_AWQOS[82] = AP_AXIMM_82_AWQOS;
            assign ap_AWVALID[82] = AP_AXIMM_82_AWVALID;
            assign AP_AXIMM_82_AWREADY = ap_AWREADY[82];
            assign ap_WDATA[82][M_AXIMM_82_DATA_WIDTH-1:0] = AP_AXIMM_82_WDATA;
            assign ap_WSTRB[82][M_AXIMM_82_DATA_WIDTH/8-1:0] = AP_AXIMM_82_WSTRB;
            assign ap_WLAST[82] = AP_AXIMM_82_WLAST;
            assign ap_WVALID[82] = AP_AXIMM_82_WVALID;
            assign AP_AXIMM_82_WREADY = ap_WREADY[82];
            assign AP_AXIMM_82_BRESP = ap_BRESP[82];
            assign AP_AXIMM_82_BVALID = ap_BVALID[82];
            assign ap_BREADY[82] = AP_AXIMM_82_BREADY;
            assign ap_ARADDR[82][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_82_ARADDR;
            assign ap_ARLEN[82] = AP_AXIMM_82_ARLEN;
            assign ap_ARSIZE[82] = AP_AXIMM_82_ARSIZE;
            assign ap_ARBURST[82] = AP_AXIMM_82_ARBURST;
            assign ap_ARLOCK[82] = AP_AXIMM_82_ARLOCK;
            assign ap_ARCACHE[82] = AP_AXIMM_82_ARCACHE;
            assign ap_ARPROT[82] = AP_AXIMM_82_ARPROT;
            assign ap_ARREGION[82] = AP_AXIMM_82_ARREGION;
            assign ap_ARQOS[82] = AP_AXIMM_82_ARQOS;
            assign ap_ARVALID[82] = AP_AXIMM_82_ARVALID;
            assign AP_AXIMM_82_ARREADY = ap_ARREADY[82];
            assign AP_AXIMM_82_RDATA = ap_RDATA[82][M_AXIMM_82_DATA_WIDTH-1:0];
            assign AP_AXIMM_82_RRESP = ap_RRESP[82];
            assign AP_AXIMM_82_RLAST = ap_RLAST[82];
            assign AP_AXIMM_82_RVALID = ap_RVALID[82];
            assign ap_RREADY[82] = AP_AXIMM_82_RREADY;
            assign M_AXIMM_82_AWADDR = dm_AWADDR[82][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_82_AWLEN = dm_AWLEN[82];
            assign M_AXIMM_82_AWSIZE = dm_AWSIZE[82];
            assign M_AXIMM_82_AWBURST = dm_AWBURST[82];
            assign M_AXIMM_82_AWLOCK = dm_AWLOCK[82];
            assign M_AXIMM_82_AWCACHE = dm_AWCACHE[82];
            assign M_AXIMM_82_AWPROT = dm_AWPROT[82];
            assign M_AXIMM_82_AWREGION = dm_AWREGION[82];
            assign M_AXIMM_82_AWQOS = dm_AWQOS[82];
            assign M_AXIMM_82_AWVALID = dm_AWVALID[82];
            assign dm_AWREADY[82] = M_AXIMM_82_AWREADY;
            assign M_AXIMM_82_WDATA = dm_WDATA[82][M_AXIMM_82_DATA_WIDTH-1:0];
            assign M_AXIMM_82_WSTRB = dm_WSTRB[82][M_AXIMM_82_DATA_WIDTH/8-1:0];
            assign M_AXIMM_82_WLAST = dm_WLAST[82];
            assign M_AXIMM_82_WVALID = dm_WVALID[82];
            assign dm_WREADY[82] = M_AXIMM_82_WREADY;
            assign dm_BRESP[82] = M_AXIMM_82_BRESP;
            assign dm_BVALID[82] = M_AXIMM_82_BVALID;
            assign M_AXIMM_82_BREADY = dm_BREADY[82];
            assign M_AXIMM_82_ARADDR = dm_ARADDR[82][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_82_ARLEN = dm_ARLEN[82];
            assign M_AXIMM_82_ARSIZE = dm_ARSIZE[82];
            assign M_AXIMM_82_ARBURST = dm_ARBURST[82];
            assign M_AXIMM_82_ARLOCK = dm_ARLOCK[82];
            assign M_AXIMM_82_ARCACHE = dm_ARCACHE[82];
            assign M_AXIMM_82_ARPROT = dm_ARPROT[82];
            assign M_AXIMM_82_ARREGION = dm_ARREGION[82];
            assign M_AXIMM_82_ARQOS = dm_ARQOS[82];
            assign M_AXIMM_82_ARVALID = dm_ARVALID[82];
            assign dm_ARREADY[82] = M_AXIMM_82_ARREADY;
            assign dm_RDATA[82][M_AXIMM_82_DATA_WIDTH-1:0] = M_AXIMM_82_RDATA;
            assign dm_RRESP[82] = M_AXIMM_82_RRESP;
            assign dm_RLAST[82] = M_AXIMM_82_RLAST;
            assign dm_RVALID[82] = M_AXIMM_82_RVALID;
            assign M_AXIMM_82_RREADY = dm_RREADY[82];
        end
        if(C_NUM_AXIMMs > 83) begin
            assign ap_AWADDR[83][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_83_AWADDR;
            assign ap_AWLEN[83] = AP_AXIMM_83_AWLEN;
            assign ap_AWSIZE[83] = AP_AXIMM_83_AWSIZE;
            assign ap_AWBURST[83] = AP_AXIMM_83_AWBURST;
            assign ap_AWLOCK[83] = AP_AXIMM_83_AWLOCK;
            assign ap_AWCACHE[83] = AP_AXIMM_83_AWCACHE;
            assign ap_AWPROT[83] = AP_AXIMM_83_AWPROT;
            assign ap_AWREGION[83] = AP_AXIMM_83_AWREGION;
            assign ap_AWQOS[83] = AP_AXIMM_83_AWQOS;
            assign ap_AWVALID[83] = AP_AXIMM_83_AWVALID;
            assign AP_AXIMM_83_AWREADY = ap_AWREADY[83];
            assign ap_WDATA[83][M_AXIMM_83_DATA_WIDTH-1:0] = AP_AXIMM_83_WDATA;
            assign ap_WSTRB[83][M_AXIMM_83_DATA_WIDTH/8-1:0] = AP_AXIMM_83_WSTRB;
            assign ap_WLAST[83] = AP_AXIMM_83_WLAST;
            assign ap_WVALID[83] = AP_AXIMM_83_WVALID;
            assign AP_AXIMM_83_WREADY = ap_WREADY[83];
            assign AP_AXIMM_83_BRESP = ap_BRESP[83];
            assign AP_AXIMM_83_BVALID = ap_BVALID[83];
            assign ap_BREADY[83] = AP_AXIMM_83_BREADY;
            assign ap_ARADDR[83][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_83_ARADDR;
            assign ap_ARLEN[83] = AP_AXIMM_83_ARLEN;
            assign ap_ARSIZE[83] = AP_AXIMM_83_ARSIZE;
            assign ap_ARBURST[83] = AP_AXIMM_83_ARBURST;
            assign ap_ARLOCK[83] = AP_AXIMM_83_ARLOCK;
            assign ap_ARCACHE[83] = AP_AXIMM_83_ARCACHE;
            assign ap_ARPROT[83] = AP_AXIMM_83_ARPROT;
            assign ap_ARREGION[83] = AP_AXIMM_83_ARREGION;
            assign ap_ARQOS[83] = AP_AXIMM_83_ARQOS;
            assign ap_ARVALID[83] = AP_AXIMM_83_ARVALID;
            assign AP_AXIMM_83_ARREADY = ap_ARREADY[83];
            assign AP_AXIMM_83_RDATA = ap_RDATA[83][M_AXIMM_83_DATA_WIDTH-1:0];
            assign AP_AXIMM_83_RRESP = ap_RRESP[83];
            assign AP_AXIMM_83_RLAST = ap_RLAST[83];
            assign AP_AXIMM_83_RVALID = ap_RVALID[83];
            assign ap_RREADY[83] = AP_AXIMM_83_RREADY;
            assign M_AXIMM_83_AWADDR = dm_AWADDR[83][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_83_AWLEN = dm_AWLEN[83];
            assign M_AXIMM_83_AWSIZE = dm_AWSIZE[83];
            assign M_AXIMM_83_AWBURST = dm_AWBURST[83];
            assign M_AXIMM_83_AWLOCK = dm_AWLOCK[83];
            assign M_AXIMM_83_AWCACHE = dm_AWCACHE[83];
            assign M_AXIMM_83_AWPROT = dm_AWPROT[83];
            assign M_AXIMM_83_AWREGION = dm_AWREGION[83];
            assign M_AXIMM_83_AWQOS = dm_AWQOS[83];
            assign M_AXIMM_83_AWVALID = dm_AWVALID[83];
            assign dm_AWREADY[83] = M_AXIMM_83_AWREADY;
            assign M_AXIMM_83_WDATA = dm_WDATA[83][M_AXIMM_83_DATA_WIDTH-1:0];
            assign M_AXIMM_83_WSTRB = dm_WSTRB[83][M_AXIMM_83_DATA_WIDTH/8-1:0];
            assign M_AXIMM_83_WLAST = dm_WLAST[83];
            assign M_AXIMM_83_WVALID = dm_WVALID[83];
            assign dm_WREADY[83] = M_AXIMM_83_WREADY;
            assign dm_BRESP[83] = M_AXIMM_83_BRESP;
            assign dm_BVALID[83] = M_AXIMM_83_BVALID;
            assign M_AXIMM_83_BREADY = dm_BREADY[83];
            assign M_AXIMM_83_ARADDR = dm_ARADDR[83][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_83_ARLEN = dm_ARLEN[83];
            assign M_AXIMM_83_ARSIZE = dm_ARSIZE[83];
            assign M_AXIMM_83_ARBURST = dm_ARBURST[83];
            assign M_AXIMM_83_ARLOCK = dm_ARLOCK[83];
            assign M_AXIMM_83_ARCACHE = dm_ARCACHE[83];
            assign M_AXIMM_83_ARPROT = dm_ARPROT[83];
            assign M_AXIMM_83_ARREGION = dm_ARREGION[83];
            assign M_AXIMM_83_ARQOS = dm_ARQOS[83];
            assign M_AXIMM_83_ARVALID = dm_ARVALID[83];
            assign dm_ARREADY[83] = M_AXIMM_83_ARREADY;
            assign dm_RDATA[83][M_AXIMM_83_DATA_WIDTH-1:0] = M_AXIMM_83_RDATA;
            assign dm_RRESP[83] = M_AXIMM_83_RRESP;
            assign dm_RLAST[83] = M_AXIMM_83_RLAST;
            assign dm_RVALID[83] = M_AXIMM_83_RVALID;
            assign M_AXIMM_83_RREADY = dm_RREADY[83];
        end
        if(C_NUM_AXIMMs > 84) begin
            assign ap_AWADDR[84][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_84_AWADDR;
            assign ap_AWLEN[84] = AP_AXIMM_84_AWLEN;
            assign ap_AWSIZE[84] = AP_AXIMM_84_AWSIZE;
            assign ap_AWBURST[84] = AP_AXIMM_84_AWBURST;
            assign ap_AWLOCK[84] = AP_AXIMM_84_AWLOCK;
            assign ap_AWCACHE[84] = AP_AXIMM_84_AWCACHE;
            assign ap_AWPROT[84] = AP_AXIMM_84_AWPROT;
            assign ap_AWREGION[84] = AP_AXIMM_84_AWREGION;
            assign ap_AWQOS[84] = AP_AXIMM_84_AWQOS;
            assign ap_AWVALID[84] = AP_AXIMM_84_AWVALID;
            assign AP_AXIMM_84_AWREADY = ap_AWREADY[84];
            assign ap_WDATA[84][M_AXIMM_84_DATA_WIDTH-1:0] = AP_AXIMM_84_WDATA;
            assign ap_WSTRB[84][M_AXIMM_84_DATA_WIDTH/8-1:0] = AP_AXIMM_84_WSTRB;
            assign ap_WLAST[84] = AP_AXIMM_84_WLAST;
            assign ap_WVALID[84] = AP_AXIMM_84_WVALID;
            assign AP_AXIMM_84_WREADY = ap_WREADY[84];
            assign AP_AXIMM_84_BRESP = ap_BRESP[84];
            assign AP_AXIMM_84_BVALID = ap_BVALID[84];
            assign ap_BREADY[84] = AP_AXIMM_84_BREADY;
            assign ap_ARADDR[84][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_84_ARADDR;
            assign ap_ARLEN[84] = AP_AXIMM_84_ARLEN;
            assign ap_ARSIZE[84] = AP_AXIMM_84_ARSIZE;
            assign ap_ARBURST[84] = AP_AXIMM_84_ARBURST;
            assign ap_ARLOCK[84] = AP_AXIMM_84_ARLOCK;
            assign ap_ARCACHE[84] = AP_AXIMM_84_ARCACHE;
            assign ap_ARPROT[84] = AP_AXIMM_84_ARPROT;
            assign ap_ARREGION[84] = AP_AXIMM_84_ARREGION;
            assign ap_ARQOS[84] = AP_AXIMM_84_ARQOS;
            assign ap_ARVALID[84] = AP_AXIMM_84_ARVALID;
            assign AP_AXIMM_84_ARREADY = ap_ARREADY[84];
            assign AP_AXIMM_84_RDATA = ap_RDATA[84][M_AXIMM_84_DATA_WIDTH-1:0];
            assign AP_AXIMM_84_RRESP = ap_RRESP[84];
            assign AP_AXIMM_84_RLAST = ap_RLAST[84];
            assign AP_AXIMM_84_RVALID = ap_RVALID[84];
            assign ap_RREADY[84] = AP_AXIMM_84_RREADY;
            assign M_AXIMM_84_AWADDR = dm_AWADDR[84][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_84_AWLEN = dm_AWLEN[84];
            assign M_AXIMM_84_AWSIZE = dm_AWSIZE[84];
            assign M_AXIMM_84_AWBURST = dm_AWBURST[84];
            assign M_AXIMM_84_AWLOCK = dm_AWLOCK[84];
            assign M_AXIMM_84_AWCACHE = dm_AWCACHE[84];
            assign M_AXIMM_84_AWPROT = dm_AWPROT[84];
            assign M_AXIMM_84_AWREGION = dm_AWREGION[84];
            assign M_AXIMM_84_AWQOS = dm_AWQOS[84];
            assign M_AXIMM_84_AWVALID = dm_AWVALID[84];
            assign dm_AWREADY[84] = M_AXIMM_84_AWREADY;
            assign M_AXIMM_84_WDATA = dm_WDATA[84][M_AXIMM_84_DATA_WIDTH-1:0];
            assign M_AXIMM_84_WSTRB = dm_WSTRB[84][M_AXIMM_84_DATA_WIDTH/8-1:0];
            assign M_AXIMM_84_WLAST = dm_WLAST[84];
            assign M_AXIMM_84_WVALID = dm_WVALID[84];
            assign dm_WREADY[84] = M_AXIMM_84_WREADY;
            assign dm_BRESP[84] = M_AXIMM_84_BRESP;
            assign dm_BVALID[84] = M_AXIMM_84_BVALID;
            assign M_AXIMM_84_BREADY = dm_BREADY[84];
            assign M_AXIMM_84_ARADDR = dm_ARADDR[84][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_84_ARLEN = dm_ARLEN[84];
            assign M_AXIMM_84_ARSIZE = dm_ARSIZE[84];
            assign M_AXIMM_84_ARBURST = dm_ARBURST[84];
            assign M_AXIMM_84_ARLOCK = dm_ARLOCK[84];
            assign M_AXIMM_84_ARCACHE = dm_ARCACHE[84];
            assign M_AXIMM_84_ARPROT = dm_ARPROT[84];
            assign M_AXIMM_84_ARREGION = dm_ARREGION[84];
            assign M_AXIMM_84_ARQOS = dm_ARQOS[84];
            assign M_AXIMM_84_ARVALID = dm_ARVALID[84];
            assign dm_ARREADY[84] = M_AXIMM_84_ARREADY;
            assign dm_RDATA[84][M_AXIMM_84_DATA_WIDTH-1:0] = M_AXIMM_84_RDATA;
            assign dm_RRESP[84] = M_AXIMM_84_RRESP;
            assign dm_RLAST[84] = M_AXIMM_84_RLAST;
            assign dm_RVALID[84] = M_AXIMM_84_RVALID;
            assign M_AXIMM_84_RREADY = dm_RREADY[84];
        end
        if(C_NUM_AXIMMs > 85) begin
            assign ap_AWADDR[85][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_85_AWADDR;
            assign ap_AWLEN[85] = AP_AXIMM_85_AWLEN;
            assign ap_AWSIZE[85] = AP_AXIMM_85_AWSIZE;
            assign ap_AWBURST[85] = AP_AXIMM_85_AWBURST;
            assign ap_AWLOCK[85] = AP_AXIMM_85_AWLOCK;
            assign ap_AWCACHE[85] = AP_AXIMM_85_AWCACHE;
            assign ap_AWPROT[85] = AP_AXIMM_85_AWPROT;
            assign ap_AWREGION[85] = AP_AXIMM_85_AWREGION;
            assign ap_AWQOS[85] = AP_AXIMM_85_AWQOS;
            assign ap_AWVALID[85] = AP_AXIMM_85_AWVALID;
            assign AP_AXIMM_85_AWREADY = ap_AWREADY[85];
            assign ap_WDATA[85][M_AXIMM_85_DATA_WIDTH-1:0] = AP_AXIMM_85_WDATA;
            assign ap_WSTRB[85][M_AXIMM_85_DATA_WIDTH/8-1:0] = AP_AXIMM_85_WSTRB;
            assign ap_WLAST[85] = AP_AXIMM_85_WLAST;
            assign ap_WVALID[85] = AP_AXIMM_85_WVALID;
            assign AP_AXIMM_85_WREADY = ap_WREADY[85];
            assign AP_AXIMM_85_BRESP = ap_BRESP[85];
            assign AP_AXIMM_85_BVALID = ap_BVALID[85];
            assign ap_BREADY[85] = AP_AXIMM_85_BREADY;
            assign ap_ARADDR[85][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_85_ARADDR;
            assign ap_ARLEN[85] = AP_AXIMM_85_ARLEN;
            assign ap_ARSIZE[85] = AP_AXIMM_85_ARSIZE;
            assign ap_ARBURST[85] = AP_AXIMM_85_ARBURST;
            assign ap_ARLOCK[85] = AP_AXIMM_85_ARLOCK;
            assign ap_ARCACHE[85] = AP_AXIMM_85_ARCACHE;
            assign ap_ARPROT[85] = AP_AXIMM_85_ARPROT;
            assign ap_ARREGION[85] = AP_AXIMM_85_ARREGION;
            assign ap_ARQOS[85] = AP_AXIMM_85_ARQOS;
            assign ap_ARVALID[85] = AP_AXIMM_85_ARVALID;
            assign AP_AXIMM_85_ARREADY = ap_ARREADY[85];
            assign AP_AXIMM_85_RDATA = ap_RDATA[85][M_AXIMM_85_DATA_WIDTH-1:0];
            assign AP_AXIMM_85_RRESP = ap_RRESP[85];
            assign AP_AXIMM_85_RLAST = ap_RLAST[85];
            assign AP_AXIMM_85_RVALID = ap_RVALID[85];
            assign ap_RREADY[85] = AP_AXIMM_85_RREADY;
            assign M_AXIMM_85_AWADDR = dm_AWADDR[85][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_85_AWLEN = dm_AWLEN[85];
            assign M_AXIMM_85_AWSIZE = dm_AWSIZE[85];
            assign M_AXIMM_85_AWBURST = dm_AWBURST[85];
            assign M_AXIMM_85_AWLOCK = dm_AWLOCK[85];
            assign M_AXIMM_85_AWCACHE = dm_AWCACHE[85];
            assign M_AXIMM_85_AWPROT = dm_AWPROT[85];
            assign M_AXIMM_85_AWREGION = dm_AWREGION[85];
            assign M_AXIMM_85_AWQOS = dm_AWQOS[85];
            assign M_AXIMM_85_AWVALID = dm_AWVALID[85];
            assign dm_AWREADY[85] = M_AXIMM_85_AWREADY;
            assign M_AXIMM_85_WDATA = dm_WDATA[85][M_AXIMM_85_DATA_WIDTH-1:0];
            assign M_AXIMM_85_WSTRB = dm_WSTRB[85][M_AXIMM_85_DATA_WIDTH/8-1:0];
            assign M_AXIMM_85_WLAST = dm_WLAST[85];
            assign M_AXIMM_85_WVALID = dm_WVALID[85];
            assign dm_WREADY[85] = M_AXIMM_85_WREADY;
            assign dm_BRESP[85] = M_AXIMM_85_BRESP;
            assign dm_BVALID[85] = M_AXIMM_85_BVALID;
            assign M_AXIMM_85_BREADY = dm_BREADY[85];
            assign M_AXIMM_85_ARADDR = dm_ARADDR[85][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_85_ARLEN = dm_ARLEN[85];
            assign M_AXIMM_85_ARSIZE = dm_ARSIZE[85];
            assign M_AXIMM_85_ARBURST = dm_ARBURST[85];
            assign M_AXIMM_85_ARLOCK = dm_ARLOCK[85];
            assign M_AXIMM_85_ARCACHE = dm_ARCACHE[85];
            assign M_AXIMM_85_ARPROT = dm_ARPROT[85];
            assign M_AXIMM_85_ARREGION = dm_ARREGION[85];
            assign M_AXIMM_85_ARQOS = dm_ARQOS[85];
            assign M_AXIMM_85_ARVALID = dm_ARVALID[85];
            assign dm_ARREADY[85] = M_AXIMM_85_ARREADY;
            assign dm_RDATA[85][M_AXIMM_85_DATA_WIDTH-1:0] = M_AXIMM_85_RDATA;
            assign dm_RRESP[85] = M_AXIMM_85_RRESP;
            assign dm_RLAST[85] = M_AXIMM_85_RLAST;
            assign dm_RVALID[85] = M_AXIMM_85_RVALID;
            assign M_AXIMM_85_RREADY = dm_RREADY[85];
        end
        if(C_NUM_AXIMMs > 86) begin
            assign ap_AWADDR[86][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_86_AWADDR;
            assign ap_AWLEN[86] = AP_AXIMM_86_AWLEN;
            assign ap_AWSIZE[86] = AP_AXIMM_86_AWSIZE;
            assign ap_AWBURST[86] = AP_AXIMM_86_AWBURST;
            assign ap_AWLOCK[86] = AP_AXIMM_86_AWLOCK;
            assign ap_AWCACHE[86] = AP_AXIMM_86_AWCACHE;
            assign ap_AWPROT[86] = AP_AXIMM_86_AWPROT;
            assign ap_AWREGION[86] = AP_AXIMM_86_AWREGION;
            assign ap_AWQOS[86] = AP_AXIMM_86_AWQOS;
            assign ap_AWVALID[86] = AP_AXIMM_86_AWVALID;
            assign AP_AXIMM_86_AWREADY = ap_AWREADY[86];
            assign ap_WDATA[86][M_AXIMM_86_DATA_WIDTH-1:0] = AP_AXIMM_86_WDATA;
            assign ap_WSTRB[86][M_AXIMM_86_DATA_WIDTH/8-1:0] = AP_AXIMM_86_WSTRB;
            assign ap_WLAST[86] = AP_AXIMM_86_WLAST;
            assign ap_WVALID[86] = AP_AXIMM_86_WVALID;
            assign AP_AXIMM_86_WREADY = ap_WREADY[86];
            assign AP_AXIMM_86_BRESP = ap_BRESP[86];
            assign AP_AXIMM_86_BVALID = ap_BVALID[86];
            assign ap_BREADY[86] = AP_AXIMM_86_BREADY;
            assign ap_ARADDR[86][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_86_ARADDR;
            assign ap_ARLEN[86] = AP_AXIMM_86_ARLEN;
            assign ap_ARSIZE[86] = AP_AXIMM_86_ARSIZE;
            assign ap_ARBURST[86] = AP_AXIMM_86_ARBURST;
            assign ap_ARLOCK[86] = AP_AXIMM_86_ARLOCK;
            assign ap_ARCACHE[86] = AP_AXIMM_86_ARCACHE;
            assign ap_ARPROT[86] = AP_AXIMM_86_ARPROT;
            assign ap_ARREGION[86] = AP_AXIMM_86_ARREGION;
            assign ap_ARQOS[86] = AP_AXIMM_86_ARQOS;
            assign ap_ARVALID[86] = AP_AXIMM_86_ARVALID;
            assign AP_AXIMM_86_ARREADY = ap_ARREADY[86];
            assign AP_AXIMM_86_RDATA = ap_RDATA[86][M_AXIMM_86_DATA_WIDTH-1:0];
            assign AP_AXIMM_86_RRESP = ap_RRESP[86];
            assign AP_AXIMM_86_RLAST = ap_RLAST[86];
            assign AP_AXIMM_86_RVALID = ap_RVALID[86];
            assign ap_RREADY[86] = AP_AXIMM_86_RREADY;
            assign M_AXIMM_86_AWADDR = dm_AWADDR[86][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_86_AWLEN = dm_AWLEN[86];
            assign M_AXIMM_86_AWSIZE = dm_AWSIZE[86];
            assign M_AXIMM_86_AWBURST = dm_AWBURST[86];
            assign M_AXIMM_86_AWLOCK = dm_AWLOCK[86];
            assign M_AXIMM_86_AWCACHE = dm_AWCACHE[86];
            assign M_AXIMM_86_AWPROT = dm_AWPROT[86];
            assign M_AXIMM_86_AWREGION = dm_AWREGION[86];
            assign M_AXIMM_86_AWQOS = dm_AWQOS[86];
            assign M_AXIMM_86_AWVALID = dm_AWVALID[86];
            assign dm_AWREADY[86] = M_AXIMM_86_AWREADY;
            assign M_AXIMM_86_WDATA = dm_WDATA[86][M_AXIMM_86_DATA_WIDTH-1:0];
            assign M_AXIMM_86_WSTRB = dm_WSTRB[86][M_AXIMM_86_DATA_WIDTH/8-1:0];
            assign M_AXIMM_86_WLAST = dm_WLAST[86];
            assign M_AXIMM_86_WVALID = dm_WVALID[86];
            assign dm_WREADY[86] = M_AXIMM_86_WREADY;
            assign dm_BRESP[86] = M_AXIMM_86_BRESP;
            assign dm_BVALID[86] = M_AXIMM_86_BVALID;
            assign M_AXIMM_86_BREADY = dm_BREADY[86];
            assign M_AXIMM_86_ARADDR = dm_ARADDR[86][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_86_ARLEN = dm_ARLEN[86];
            assign M_AXIMM_86_ARSIZE = dm_ARSIZE[86];
            assign M_AXIMM_86_ARBURST = dm_ARBURST[86];
            assign M_AXIMM_86_ARLOCK = dm_ARLOCK[86];
            assign M_AXIMM_86_ARCACHE = dm_ARCACHE[86];
            assign M_AXIMM_86_ARPROT = dm_ARPROT[86];
            assign M_AXIMM_86_ARREGION = dm_ARREGION[86];
            assign M_AXIMM_86_ARQOS = dm_ARQOS[86];
            assign M_AXIMM_86_ARVALID = dm_ARVALID[86];
            assign dm_ARREADY[86] = M_AXIMM_86_ARREADY;
            assign dm_RDATA[86][M_AXIMM_86_DATA_WIDTH-1:0] = M_AXIMM_86_RDATA;
            assign dm_RRESP[86] = M_AXIMM_86_RRESP;
            assign dm_RLAST[86] = M_AXIMM_86_RLAST;
            assign dm_RVALID[86] = M_AXIMM_86_RVALID;
            assign M_AXIMM_86_RREADY = dm_RREADY[86];
        end
        if(C_NUM_AXIMMs > 87) begin
            assign ap_AWADDR[87][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_87_AWADDR;
            assign ap_AWLEN[87] = AP_AXIMM_87_AWLEN;
            assign ap_AWSIZE[87] = AP_AXIMM_87_AWSIZE;
            assign ap_AWBURST[87] = AP_AXIMM_87_AWBURST;
            assign ap_AWLOCK[87] = AP_AXIMM_87_AWLOCK;
            assign ap_AWCACHE[87] = AP_AXIMM_87_AWCACHE;
            assign ap_AWPROT[87] = AP_AXIMM_87_AWPROT;
            assign ap_AWREGION[87] = AP_AXIMM_87_AWREGION;
            assign ap_AWQOS[87] = AP_AXIMM_87_AWQOS;
            assign ap_AWVALID[87] = AP_AXIMM_87_AWVALID;
            assign AP_AXIMM_87_AWREADY = ap_AWREADY[87];
            assign ap_WDATA[87][M_AXIMM_87_DATA_WIDTH-1:0] = AP_AXIMM_87_WDATA;
            assign ap_WSTRB[87][M_AXIMM_87_DATA_WIDTH/8-1:0] = AP_AXIMM_87_WSTRB;
            assign ap_WLAST[87] = AP_AXIMM_87_WLAST;
            assign ap_WVALID[87] = AP_AXIMM_87_WVALID;
            assign AP_AXIMM_87_WREADY = ap_WREADY[87];
            assign AP_AXIMM_87_BRESP = ap_BRESP[87];
            assign AP_AXIMM_87_BVALID = ap_BVALID[87];
            assign ap_BREADY[87] = AP_AXIMM_87_BREADY;
            assign ap_ARADDR[87][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_87_ARADDR;
            assign ap_ARLEN[87] = AP_AXIMM_87_ARLEN;
            assign ap_ARSIZE[87] = AP_AXIMM_87_ARSIZE;
            assign ap_ARBURST[87] = AP_AXIMM_87_ARBURST;
            assign ap_ARLOCK[87] = AP_AXIMM_87_ARLOCK;
            assign ap_ARCACHE[87] = AP_AXIMM_87_ARCACHE;
            assign ap_ARPROT[87] = AP_AXIMM_87_ARPROT;
            assign ap_ARREGION[87] = AP_AXIMM_87_ARREGION;
            assign ap_ARQOS[87] = AP_AXIMM_87_ARQOS;
            assign ap_ARVALID[87] = AP_AXIMM_87_ARVALID;
            assign AP_AXIMM_87_ARREADY = ap_ARREADY[87];
            assign AP_AXIMM_87_RDATA = ap_RDATA[87][M_AXIMM_87_DATA_WIDTH-1:0];
            assign AP_AXIMM_87_RRESP = ap_RRESP[87];
            assign AP_AXIMM_87_RLAST = ap_RLAST[87];
            assign AP_AXIMM_87_RVALID = ap_RVALID[87];
            assign ap_RREADY[87] = AP_AXIMM_87_RREADY;
            assign M_AXIMM_87_AWADDR = dm_AWADDR[87][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_87_AWLEN = dm_AWLEN[87];
            assign M_AXIMM_87_AWSIZE = dm_AWSIZE[87];
            assign M_AXIMM_87_AWBURST = dm_AWBURST[87];
            assign M_AXIMM_87_AWLOCK = dm_AWLOCK[87];
            assign M_AXIMM_87_AWCACHE = dm_AWCACHE[87];
            assign M_AXIMM_87_AWPROT = dm_AWPROT[87];
            assign M_AXIMM_87_AWREGION = dm_AWREGION[87];
            assign M_AXIMM_87_AWQOS = dm_AWQOS[87];
            assign M_AXIMM_87_AWVALID = dm_AWVALID[87];
            assign dm_AWREADY[87] = M_AXIMM_87_AWREADY;
            assign M_AXIMM_87_WDATA = dm_WDATA[87][M_AXIMM_87_DATA_WIDTH-1:0];
            assign M_AXIMM_87_WSTRB = dm_WSTRB[87][M_AXIMM_87_DATA_WIDTH/8-1:0];
            assign M_AXIMM_87_WLAST = dm_WLAST[87];
            assign M_AXIMM_87_WVALID = dm_WVALID[87];
            assign dm_WREADY[87] = M_AXIMM_87_WREADY;
            assign dm_BRESP[87] = M_AXIMM_87_BRESP;
            assign dm_BVALID[87] = M_AXIMM_87_BVALID;
            assign M_AXIMM_87_BREADY = dm_BREADY[87];
            assign M_AXIMM_87_ARADDR = dm_ARADDR[87][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_87_ARLEN = dm_ARLEN[87];
            assign M_AXIMM_87_ARSIZE = dm_ARSIZE[87];
            assign M_AXIMM_87_ARBURST = dm_ARBURST[87];
            assign M_AXIMM_87_ARLOCK = dm_ARLOCK[87];
            assign M_AXIMM_87_ARCACHE = dm_ARCACHE[87];
            assign M_AXIMM_87_ARPROT = dm_ARPROT[87];
            assign M_AXIMM_87_ARREGION = dm_ARREGION[87];
            assign M_AXIMM_87_ARQOS = dm_ARQOS[87];
            assign M_AXIMM_87_ARVALID = dm_ARVALID[87];
            assign dm_ARREADY[87] = M_AXIMM_87_ARREADY;
            assign dm_RDATA[87][M_AXIMM_87_DATA_WIDTH-1:0] = M_AXIMM_87_RDATA;
            assign dm_RRESP[87] = M_AXIMM_87_RRESP;
            assign dm_RLAST[87] = M_AXIMM_87_RLAST;
            assign dm_RVALID[87] = M_AXIMM_87_RVALID;
            assign M_AXIMM_87_RREADY = dm_RREADY[87];
        end
        if(C_NUM_AXIMMs > 88) begin
            assign ap_AWADDR[88][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_88_AWADDR;
            assign ap_AWLEN[88] = AP_AXIMM_88_AWLEN;
            assign ap_AWSIZE[88] = AP_AXIMM_88_AWSIZE;
            assign ap_AWBURST[88] = AP_AXIMM_88_AWBURST;
            assign ap_AWLOCK[88] = AP_AXIMM_88_AWLOCK;
            assign ap_AWCACHE[88] = AP_AXIMM_88_AWCACHE;
            assign ap_AWPROT[88] = AP_AXIMM_88_AWPROT;
            assign ap_AWREGION[88] = AP_AXIMM_88_AWREGION;
            assign ap_AWQOS[88] = AP_AXIMM_88_AWQOS;
            assign ap_AWVALID[88] = AP_AXIMM_88_AWVALID;
            assign AP_AXIMM_88_AWREADY = ap_AWREADY[88];
            assign ap_WDATA[88][M_AXIMM_88_DATA_WIDTH-1:0] = AP_AXIMM_88_WDATA;
            assign ap_WSTRB[88][M_AXIMM_88_DATA_WIDTH/8-1:0] = AP_AXIMM_88_WSTRB;
            assign ap_WLAST[88] = AP_AXIMM_88_WLAST;
            assign ap_WVALID[88] = AP_AXIMM_88_WVALID;
            assign AP_AXIMM_88_WREADY = ap_WREADY[88];
            assign AP_AXIMM_88_BRESP = ap_BRESP[88];
            assign AP_AXIMM_88_BVALID = ap_BVALID[88];
            assign ap_BREADY[88] = AP_AXIMM_88_BREADY;
            assign ap_ARADDR[88][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_88_ARADDR;
            assign ap_ARLEN[88] = AP_AXIMM_88_ARLEN;
            assign ap_ARSIZE[88] = AP_AXIMM_88_ARSIZE;
            assign ap_ARBURST[88] = AP_AXIMM_88_ARBURST;
            assign ap_ARLOCK[88] = AP_AXIMM_88_ARLOCK;
            assign ap_ARCACHE[88] = AP_AXIMM_88_ARCACHE;
            assign ap_ARPROT[88] = AP_AXIMM_88_ARPROT;
            assign ap_ARREGION[88] = AP_AXIMM_88_ARREGION;
            assign ap_ARQOS[88] = AP_AXIMM_88_ARQOS;
            assign ap_ARVALID[88] = AP_AXIMM_88_ARVALID;
            assign AP_AXIMM_88_ARREADY = ap_ARREADY[88];
            assign AP_AXIMM_88_RDATA = ap_RDATA[88][M_AXIMM_88_DATA_WIDTH-1:0];
            assign AP_AXIMM_88_RRESP = ap_RRESP[88];
            assign AP_AXIMM_88_RLAST = ap_RLAST[88];
            assign AP_AXIMM_88_RVALID = ap_RVALID[88];
            assign ap_RREADY[88] = AP_AXIMM_88_RREADY;
            assign M_AXIMM_88_AWADDR = dm_AWADDR[88][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_88_AWLEN = dm_AWLEN[88];
            assign M_AXIMM_88_AWSIZE = dm_AWSIZE[88];
            assign M_AXIMM_88_AWBURST = dm_AWBURST[88];
            assign M_AXIMM_88_AWLOCK = dm_AWLOCK[88];
            assign M_AXIMM_88_AWCACHE = dm_AWCACHE[88];
            assign M_AXIMM_88_AWPROT = dm_AWPROT[88];
            assign M_AXIMM_88_AWREGION = dm_AWREGION[88];
            assign M_AXIMM_88_AWQOS = dm_AWQOS[88];
            assign M_AXIMM_88_AWVALID = dm_AWVALID[88];
            assign dm_AWREADY[88] = M_AXIMM_88_AWREADY;
            assign M_AXIMM_88_WDATA = dm_WDATA[88][M_AXIMM_88_DATA_WIDTH-1:0];
            assign M_AXIMM_88_WSTRB = dm_WSTRB[88][M_AXIMM_88_DATA_WIDTH/8-1:0];
            assign M_AXIMM_88_WLAST = dm_WLAST[88];
            assign M_AXIMM_88_WVALID = dm_WVALID[88];
            assign dm_WREADY[88] = M_AXIMM_88_WREADY;
            assign dm_BRESP[88] = M_AXIMM_88_BRESP;
            assign dm_BVALID[88] = M_AXIMM_88_BVALID;
            assign M_AXIMM_88_BREADY = dm_BREADY[88];
            assign M_AXIMM_88_ARADDR = dm_ARADDR[88][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_88_ARLEN = dm_ARLEN[88];
            assign M_AXIMM_88_ARSIZE = dm_ARSIZE[88];
            assign M_AXIMM_88_ARBURST = dm_ARBURST[88];
            assign M_AXIMM_88_ARLOCK = dm_ARLOCK[88];
            assign M_AXIMM_88_ARCACHE = dm_ARCACHE[88];
            assign M_AXIMM_88_ARPROT = dm_ARPROT[88];
            assign M_AXIMM_88_ARREGION = dm_ARREGION[88];
            assign M_AXIMM_88_ARQOS = dm_ARQOS[88];
            assign M_AXIMM_88_ARVALID = dm_ARVALID[88];
            assign dm_ARREADY[88] = M_AXIMM_88_ARREADY;
            assign dm_RDATA[88][M_AXIMM_88_DATA_WIDTH-1:0] = M_AXIMM_88_RDATA;
            assign dm_RRESP[88] = M_AXIMM_88_RRESP;
            assign dm_RLAST[88] = M_AXIMM_88_RLAST;
            assign dm_RVALID[88] = M_AXIMM_88_RVALID;
            assign M_AXIMM_88_RREADY = dm_RREADY[88];
        end
        if(C_NUM_AXIMMs > 89) begin
            assign ap_AWADDR[89][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_89_AWADDR;
            assign ap_AWLEN[89] = AP_AXIMM_89_AWLEN;
            assign ap_AWSIZE[89] = AP_AXIMM_89_AWSIZE;
            assign ap_AWBURST[89] = AP_AXIMM_89_AWBURST;
            assign ap_AWLOCK[89] = AP_AXIMM_89_AWLOCK;
            assign ap_AWCACHE[89] = AP_AXIMM_89_AWCACHE;
            assign ap_AWPROT[89] = AP_AXIMM_89_AWPROT;
            assign ap_AWREGION[89] = AP_AXIMM_89_AWREGION;
            assign ap_AWQOS[89] = AP_AXIMM_89_AWQOS;
            assign ap_AWVALID[89] = AP_AXIMM_89_AWVALID;
            assign AP_AXIMM_89_AWREADY = ap_AWREADY[89];
            assign ap_WDATA[89][M_AXIMM_89_DATA_WIDTH-1:0] = AP_AXIMM_89_WDATA;
            assign ap_WSTRB[89][M_AXIMM_89_DATA_WIDTH/8-1:0] = AP_AXIMM_89_WSTRB;
            assign ap_WLAST[89] = AP_AXIMM_89_WLAST;
            assign ap_WVALID[89] = AP_AXIMM_89_WVALID;
            assign AP_AXIMM_89_WREADY = ap_WREADY[89];
            assign AP_AXIMM_89_BRESP = ap_BRESP[89];
            assign AP_AXIMM_89_BVALID = ap_BVALID[89];
            assign ap_BREADY[89] = AP_AXIMM_89_BREADY;
            assign ap_ARADDR[89][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_89_ARADDR;
            assign ap_ARLEN[89] = AP_AXIMM_89_ARLEN;
            assign ap_ARSIZE[89] = AP_AXIMM_89_ARSIZE;
            assign ap_ARBURST[89] = AP_AXIMM_89_ARBURST;
            assign ap_ARLOCK[89] = AP_AXIMM_89_ARLOCK;
            assign ap_ARCACHE[89] = AP_AXIMM_89_ARCACHE;
            assign ap_ARPROT[89] = AP_AXIMM_89_ARPROT;
            assign ap_ARREGION[89] = AP_AXIMM_89_ARREGION;
            assign ap_ARQOS[89] = AP_AXIMM_89_ARQOS;
            assign ap_ARVALID[89] = AP_AXIMM_89_ARVALID;
            assign AP_AXIMM_89_ARREADY = ap_ARREADY[89];
            assign AP_AXIMM_89_RDATA = ap_RDATA[89][M_AXIMM_89_DATA_WIDTH-1:0];
            assign AP_AXIMM_89_RRESP = ap_RRESP[89];
            assign AP_AXIMM_89_RLAST = ap_RLAST[89];
            assign AP_AXIMM_89_RVALID = ap_RVALID[89];
            assign ap_RREADY[89] = AP_AXIMM_89_RREADY;
            assign M_AXIMM_89_AWADDR = dm_AWADDR[89][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_89_AWLEN = dm_AWLEN[89];
            assign M_AXIMM_89_AWSIZE = dm_AWSIZE[89];
            assign M_AXIMM_89_AWBURST = dm_AWBURST[89];
            assign M_AXIMM_89_AWLOCK = dm_AWLOCK[89];
            assign M_AXIMM_89_AWCACHE = dm_AWCACHE[89];
            assign M_AXIMM_89_AWPROT = dm_AWPROT[89];
            assign M_AXIMM_89_AWREGION = dm_AWREGION[89];
            assign M_AXIMM_89_AWQOS = dm_AWQOS[89];
            assign M_AXIMM_89_AWVALID = dm_AWVALID[89];
            assign dm_AWREADY[89] = M_AXIMM_89_AWREADY;
            assign M_AXIMM_89_WDATA = dm_WDATA[89][M_AXIMM_89_DATA_WIDTH-1:0];
            assign M_AXIMM_89_WSTRB = dm_WSTRB[89][M_AXIMM_89_DATA_WIDTH/8-1:0];
            assign M_AXIMM_89_WLAST = dm_WLAST[89];
            assign M_AXIMM_89_WVALID = dm_WVALID[89];
            assign dm_WREADY[89] = M_AXIMM_89_WREADY;
            assign dm_BRESP[89] = M_AXIMM_89_BRESP;
            assign dm_BVALID[89] = M_AXIMM_89_BVALID;
            assign M_AXIMM_89_BREADY = dm_BREADY[89];
            assign M_AXIMM_89_ARADDR = dm_ARADDR[89][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_89_ARLEN = dm_ARLEN[89];
            assign M_AXIMM_89_ARSIZE = dm_ARSIZE[89];
            assign M_AXIMM_89_ARBURST = dm_ARBURST[89];
            assign M_AXIMM_89_ARLOCK = dm_ARLOCK[89];
            assign M_AXIMM_89_ARCACHE = dm_ARCACHE[89];
            assign M_AXIMM_89_ARPROT = dm_ARPROT[89];
            assign M_AXIMM_89_ARREGION = dm_ARREGION[89];
            assign M_AXIMM_89_ARQOS = dm_ARQOS[89];
            assign M_AXIMM_89_ARVALID = dm_ARVALID[89];
            assign dm_ARREADY[89] = M_AXIMM_89_ARREADY;
            assign dm_RDATA[89][M_AXIMM_89_DATA_WIDTH-1:0] = M_AXIMM_89_RDATA;
            assign dm_RRESP[89] = M_AXIMM_89_RRESP;
            assign dm_RLAST[89] = M_AXIMM_89_RLAST;
            assign dm_RVALID[89] = M_AXIMM_89_RVALID;
            assign M_AXIMM_89_RREADY = dm_RREADY[89];
        end
        if(C_NUM_AXIMMs > 90) begin
            assign ap_AWADDR[90][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_90_AWADDR;
            assign ap_AWLEN[90] = AP_AXIMM_90_AWLEN;
            assign ap_AWSIZE[90] = AP_AXIMM_90_AWSIZE;
            assign ap_AWBURST[90] = AP_AXIMM_90_AWBURST;
            assign ap_AWLOCK[90] = AP_AXIMM_90_AWLOCK;
            assign ap_AWCACHE[90] = AP_AXIMM_90_AWCACHE;
            assign ap_AWPROT[90] = AP_AXIMM_90_AWPROT;
            assign ap_AWREGION[90] = AP_AXIMM_90_AWREGION;
            assign ap_AWQOS[90] = AP_AXIMM_90_AWQOS;
            assign ap_AWVALID[90] = AP_AXIMM_90_AWVALID;
            assign AP_AXIMM_90_AWREADY = ap_AWREADY[90];
            assign ap_WDATA[90][M_AXIMM_90_DATA_WIDTH-1:0] = AP_AXIMM_90_WDATA;
            assign ap_WSTRB[90][M_AXIMM_90_DATA_WIDTH/8-1:0] = AP_AXIMM_90_WSTRB;
            assign ap_WLAST[90] = AP_AXIMM_90_WLAST;
            assign ap_WVALID[90] = AP_AXIMM_90_WVALID;
            assign AP_AXIMM_90_WREADY = ap_WREADY[90];
            assign AP_AXIMM_90_BRESP = ap_BRESP[90];
            assign AP_AXIMM_90_BVALID = ap_BVALID[90];
            assign ap_BREADY[90] = AP_AXIMM_90_BREADY;
            assign ap_ARADDR[90][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_90_ARADDR;
            assign ap_ARLEN[90] = AP_AXIMM_90_ARLEN;
            assign ap_ARSIZE[90] = AP_AXIMM_90_ARSIZE;
            assign ap_ARBURST[90] = AP_AXIMM_90_ARBURST;
            assign ap_ARLOCK[90] = AP_AXIMM_90_ARLOCK;
            assign ap_ARCACHE[90] = AP_AXIMM_90_ARCACHE;
            assign ap_ARPROT[90] = AP_AXIMM_90_ARPROT;
            assign ap_ARREGION[90] = AP_AXIMM_90_ARREGION;
            assign ap_ARQOS[90] = AP_AXIMM_90_ARQOS;
            assign ap_ARVALID[90] = AP_AXIMM_90_ARVALID;
            assign AP_AXIMM_90_ARREADY = ap_ARREADY[90];
            assign AP_AXIMM_90_RDATA = ap_RDATA[90][M_AXIMM_90_DATA_WIDTH-1:0];
            assign AP_AXIMM_90_RRESP = ap_RRESP[90];
            assign AP_AXIMM_90_RLAST = ap_RLAST[90];
            assign AP_AXIMM_90_RVALID = ap_RVALID[90];
            assign ap_RREADY[90] = AP_AXIMM_90_RREADY;
            assign M_AXIMM_90_AWADDR = dm_AWADDR[90][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_90_AWLEN = dm_AWLEN[90];
            assign M_AXIMM_90_AWSIZE = dm_AWSIZE[90];
            assign M_AXIMM_90_AWBURST = dm_AWBURST[90];
            assign M_AXIMM_90_AWLOCK = dm_AWLOCK[90];
            assign M_AXIMM_90_AWCACHE = dm_AWCACHE[90];
            assign M_AXIMM_90_AWPROT = dm_AWPROT[90];
            assign M_AXIMM_90_AWREGION = dm_AWREGION[90];
            assign M_AXIMM_90_AWQOS = dm_AWQOS[90];
            assign M_AXIMM_90_AWVALID = dm_AWVALID[90];
            assign dm_AWREADY[90] = M_AXIMM_90_AWREADY;
            assign M_AXIMM_90_WDATA = dm_WDATA[90][M_AXIMM_90_DATA_WIDTH-1:0];
            assign M_AXIMM_90_WSTRB = dm_WSTRB[90][M_AXIMM_90_DATA_WIDTH/8-1:0];
            assign M_AXIMM_90_WLAST = dm_WLAST[90];
            assign M_AXIMM_90_WVALID = dm_WVALID[90];
            assign dm_WREADY[90] = M_AXIMM_90_WREADY;
            assign dm_BRESP[90] = M_AXIMM_90_BRESP;
            assign dm_BVALID[90] = M_AXIMM_90_BVALID;
            assign M_AXIMM_90_BREADY = dm_BREADY[90];
            assign M_AXIMM_90_ARADDR = dm_ARADDR[90][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_90_ARLEN = dm_ARLEN[90];
            assign M_AXIMM_90_ARSIZE = dm_ARSIZE[90];
            assign M_AXIMM_90_ARBURST = dm_ARBURST[90];
            assign M_AXIMM_90_ARLOCK = dm_ARLOCK[90];
            assign M_AXIMM_90_ARCACHE = dm_ARCACHE[90];
            assign M_AXIMM_90_ARPROT = dm_ARPROT[90];
            assign M_AXIMM_90_ARREGION = dm_ARREGION[90];
            assign M_AXIMM_90_ARQOS = dm_ARQOS[90];
            assign M_AXIMM_90_ARVALID = dm_ARVALID[90];
            assign dm_ARREADY[90] = M_AXIMM_90_ARREADY;
            assign dm_RDATA[90][M_AXIMM_90_DATA_WIDTH-1:0] = M_AXIMM_90_RDATA;
            assign dm_RRESP[90] = M_AXIMM_90_RRESP;
            assign dm_RLAST[90] = M_AXIMM_90_RLAST;
            assign dm_RVALID[90] = M_AXIMM_90_RVALID;
            assign M_AXIMM_90_RREADY = dm_RREADY[90];
        end
        if(C_NUM_AXIMMs > 91) begin
            assign ap_AWADDR[91][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_91_AWADDR;
            assign ap_AWLEN[91] = AP_AXIMM_91_AWLEN;
            assign ap_AWSIZE[91] = AP_AXIMM_91_AWSIZE;
            assign ap_AWBURST[91] = AP_AXIMM_91_AWBURST;
            assign ap_AWLOCK[91] = AP_AXIMM_91_AWLOCK;
            assign ap_AWCACHE[91] = AP_AXIMM_91_AWCACHE;
            assign ap_AWPROT[91] = AP_AXIMM_91_AWPROT;
            assign ap_AWREGION[91] = AP_AXIMM_91_AWREGION;
            assign ap_AWQOS[91] = AP_AXIMM_91_AWQOS;
            assign ap_AWVALID[91] = AP_AXIMM_91_AWVALID;
            assign AP_AXIMM_91_AWREADY = ap_AWREADY[91];
            assign ap_WDATA[91][M_AXIMM_91_DATA_WIDTH-1:0] = AP_AXIMM_91_WDATA;
            assign ap_WSTRB[91][M_AXIMM_91_DATA_WIDTH/8-1:0] = AP_AXIMM_91_WSTRB;
            assign ap_WLAST[91] = AP_AXIMM_91_WLAST;
            assign ap_WVALID[91] = AP_AXIMM_91_WVALID;
            assign AP_AXIMM_91_WREADY = ap_WREADY[91];
            assign AP_AXIMM_91_BRESP = ap_BRESP[91];
            assign AP_AXIMM_91_BVALID = ap_BVALID[91];
            assign ap_BREADY[91] = AP_AXIMM_91_BREADY;
            assign ap_ARADDR[91][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_91_ARADDR;
            assign ap_ARLEN[91] = AP_AXIMM_91_ARLEN;
            assign ap_ARSIZE[91] = AP_AXIMM_91_ARSIZE;
            assign ap_ARBURST[91] = AP_AXIMM_91_ARBURST;
            assign ap_ARLOCK[91] = AP_AXIMM_91_ARLOCK;
            assign ap_ARCACHE[91] = AP_AXIMM_91_ARCACHE;
            assign ap_ARPROT[91] = AP_AXIMM_91_ARPROT;
            assign ap_ARREGION[91] = AP_AXIMM_91_ARREGION;
            assign ap_ARQOS[91] = AP_AXIMM_91_ARQOS;
            assign ap_ARVALID[91] = AP_AXIMM_91_ARVALID;
            assign AP_AXIMM_91_ARREADY = ap_ARREADY[91];
            assign AP_AXIMM_91_RDATA = ap_RDATA[91][M_AXIMM_91_DATA_WIDTH-1:0];
            assign AP_AXIMM_91_RRESP = ap_RRESP[91];
            assign AP_AXIMM_91_RLAST = ap_RLAST[91];
            assign AP_AXIMM_91_RVALID = ap_RVALID[91];
            assign ap_RREADY[91] = AP_AXIMM_91_RREADY;
            assign M_AXIMM_91_AWADDR = dm_AWADDR[91][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_91_AWLEN = dm_AWLEN[91];
            assign M_AXIMM_91_AWSIZE = dm_AWSIZE[91];
            assign M_AXIMM_91_AWBURST = dm_AWBURST[91];
            assign M_AXIMM_91_AWLOCK = dm_AWLOCK[91];
            assign M_AXIMM_91_AWCACHE = dm_AWCACHE[91];
            assign M_AXIMM_91_AWPROT = dm_AWPROT[91];
            assign M_AXIMM_91_AWREGION = dm_AWREGION[91];
            assign M_AXIMM_91_AWQOS = dm_AWQOS[91];
            assign M_AXIMM_91_AWVALID = dm_AWVALID[91];
            assign dm_AWREADY[91] = M_AXIMM_91_AWREADY;
            assign M_AXIMM_91_WDATA = dm_WDATA[91][M_AXIMM_91_DATA_WIDTH-1:0];
            assign M_AXIMM_91_WSTRB = dm_WSTRB[91][M_AXIMM_91_DATA_WIDTH/8-1:0];
            assign M_AXIMM_91_WLAST = dm_WLAST[91];
            assign M_AXIMM_91_WVALID = dm_WVALID[91];
            assign dm_WREADY[91] = M_AXIMM_91_WREADY;
            assign dm_BRESP[91] = M_AXIMM_91_BRESP;
            assign dm_BVALID[91] = M_AXIMM_91_BVALID;
            assign M_AXIMM_91_BREADY = dm_BREADY[91];
            assign M_AXIMM_91_ARADDR = dm_ARADDR[91][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_91_ARLEN = dm_ARLEN[91];
            assign M_AXIMM_91_ARSIZE = dm_ARSIZE[91];
            assign M_AXIMM_91_ARBURST = dm_ARBURST[91];
            assign M_AXIMM_91_ARLOCK = dm_ARLOCK[91];
            assign M_AXIMM_91_ARCACHE = dm_ARCACHE[91];
            assign M_AXIMM_91_ARPROT = dm_ARPROT[91];
            assign M_AXIMM_91_ARREGION = dm_ARREGION[91];
            assign M_AXIMM_91_ARQOS = dm_ARQOS[91];
            assign M_AXIMM_91_ARVALID = dm_ARVALID[91];
            assign dm_ARREADY[91] = M_AXIMM_91_ARREADY;
            assign dm_RDATA[91][M_AXIMM_91_DATA_WIDTH-1:0] = M_AXIMM_91_RDATA;
            assign dm_RRESP[91] = M_AXIMM_91_RRESP;
            assign dm_RLAST[91] = M_AXIMM_91_RLAST;
            assign dm_RVALID[91] = M_AXIMM_91_RVALID;
            assign M_AXIMM_91_RREADY = dm_RREADY[91];
        end
        if(C_NUM_AXIMMs > 92) begin
            assign ap_AWADDR[92][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_92_AWADDR;
            assign ap_AWLEN[92] = AP_AXIMM_92_AWLEN;
            assign ap_AWSIZE[92] = AP_AXIMM_92_AWSIZE;
            assign ap_AWBURST[92] = AP_AXIMM_92_AWBURST;
            assign ap_AWLOCK[92] = AP_AXIMM_92_AWLOCK;
            assign ap_AWCACHE[92] = AP_AXIMM_92_AWCACHE;
            assign ap_AWPROT[92] = AP_AXIMM_92_AWPROT;
            assign ap_AWREGION[92] = AP_AXIMM_92_AWREGION;
            assign ap_AWQOS[92] = AP_AXIMM_92_AWQOS;
            assign ap_AWVALID[92] = AP_AXIMM_92_AWVALID;
            assign AP_AXIMM_92_AWREADY = ap_AWREADY[92];
            assign ap_WDATA[92][M_AXIMM_92_DATA_WIDTH-1:0] = AP_AXIMM_92_WDATA;
            assign ap_WSTRB[92][M_AXIMM_92_DATA_WIDTH/8-1:0] = AP_AXIMM_92_WSTRB;
            assign ap_WLAST[92] = AP_AXIMM_92_WLAST;
            assign ap_WVALID[92] = AP_AXIMM_92_WVALID;
            assign AP_AXIMM_92_WREADY = ap_WREADY[92];
            assign AP_AXIMM_92_BRESP = ap_BRESP[92];
            assign AP_AXIMM_92_BVALID = ap_BVALID[92];
            assign ap_BREADY[92] = AP_AXIMM_92_BREADY;
            assign ap_ARADDR[92][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_92_ARADDR;
            assign ap_ARLEN[92] = AP_AXIMM_92_ARLEN;
            assign ap_ARSIZE[92] = AP_AXIMM_92_ARSIZE;
            assign ap_ARBURST[92] = AP_AXIMM_92_ARBURST;
            assign ap_ARLOCK[92] = AP_AXIMM_92_ARLOCK;
            assign ap_ARCACHE[92] = AP_AXIMM_92_ARCACHE;
            assign ap_ARPROT[92] = AP_AXIMM_92_ARPROT;
            assign ap_ARREGION[92] = AP_AXIMM_92_ARREGION;
            assign ap_ARQOS[92] = AP_AXIMM_92_ARQOS;
            assign ap_ARVALID[92] = AP_AXIMM_92_ARVALID;
            assign AP_AXIMM_92_ARREADY = ap_ARREADY[92];
            assign AP_AXIMM_92_RDATA = ap_RDATA[92][M_AXIMM_92_DATA_WIDTH-1:0];
            assign AP_AXIMM_92_RRESP = ap_RRESP[92];
            assign AP_AXIMM_92_RLAST = ap_RLAST[92];
            assign AP_AXIMM_92_RVALID = ap_RVALID[92];
            assign ap_RREADY[92] = AP_AXIMM_92_RREADY;
            assign M_AXIMM_92_AWADDR = dm_AWADDR[92][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_92_AWLEN = dm_AWLEN[92];
            assign M_AXIMM_92_AWSIZE = dm_AWSIZE[92];
            assign M_AXIMM_92_AWBURST = dm_AWBURST[92];
            assign M_AXIMM_92_AWLOCK = dm_AWLOCK[92];
            assign M_AXIMM_92_AWCACHE = dm_AWCACHE[92];
            assign M_AXIMM_92_AWPROT = dm_AWPROT[92];
            assign M_AXIMM_92_AWREGION = dm_AWREGION[92];
            assign M_AXIMM_92_AWQOS = dm_AWQOS[92];
            assign M_AXIMM_92_AWVALID = dm_AWVALID[92];
            assign dm_AWREADY[92] = M_AXIMM_92_AWREADY;
            assign M_AXIMM_92_WDATA = dm_WDATA[92][M_AXIMM_92_DATA_WIDTH-1:0];
            assign M_AXIMM_92_WSTRB = dm_WSTRB[92][M_AXIMM_92_DATA_WIDTH/8-1:0];
            assign M_AXIMM_92_WLAST = dm_WLAST[92];
            assign M_AXIMM_92_WVALID = dm_WVALID[92];
            assign dm_WREADY[92] = M_AXIMM_92_WREADY;
            assign dm_BRESP[92] = M_AXIMM_92_BRESP;
            assign dm_BVALID[92] = M_AXIMM_92_BVALID;
            assign M_AXIMM_92_BREADY = dm_BREADY[92];
            assign M_AXIMM_92_ARADDR = dm_ARADDR[92][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_92_ARLEN = dm_ARLEN[92];
            assign M_AXIMM_92_ARSIZE = dm_ARSIZE[92];
            assign M_AXIMM_92_ARBURST = dm_ARBURST[92];
            assign M_AXIMM_92_ARLOCK = dm_ARLOCK[92];
            assign M_AXIMM_92_ARCACHE = dm_ARCACHE[92];
            assign M_AXIMM_92_ARPROT = dm_ARPROT[92];
            assign M_AXIMM_92_ARREGION = dm_ARREGION[92];
            assign M_AXIMM_92_ARQOS = dm_ARQOS[92];
            assign M_AXIMM_92_ARVALID = dm_ARVALID[92];
            assign dm_ARREADY[92] = M_AXIMM_92_ARREADY;
            assign dm_RDATA[92][M_AXIMM_92_DATA_WIDTH-1:0] = M_AXIMM_92_RDATA;
            assign dm_RRESP[92] = M_AXIMM_92_RRESP;
            assign dm_RLAST[92] = M_AXIMM_92_RLAST;
            assign dm_RVALID[92] = M_AXIMM_92_RVALID;
            assign M_AXIMM_92_RREADY = dm_RREADY[92];
        end
        if(C_NUM_AXIMMs > 93) begin
            assign ap_AWADDR[93][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_93_AWADDR;
            assign ap_AWLEN[93] = AP_AXIMM_93_AWLEN;
            assign ap_AWSIZE[93] = AP_AXIMM_93_AWSIZE;
            assign ap_AWBURST[93] = AP_AXIMM_93_AWBURST;
            assign ap_AWLOCK[93] = AP_AXIMM_93_AWLOCK;
            assign ap_AWCACHE[93] = AP_AXIMM_93_AWCACHE;
            assign ap_AWPROT[93] = AP_AXIMM_93_AWPROT;
            assign ap_AWREGION[93] = AP_AXIMM_93_AWREGION;
            assign ap_AWQOS[93] = AP_AXIMM_93_AWQOS;
            assign ap_AWVALID[93] = AP_AXIMM_93_AWVALID;
            assign AP_AXIMM_93_AWREADY = ap_AWREADY[93];
            assign ap_WDATA[93][M_AXIMM_93_DATA_WIDTH-1:0] = AP_AXIMM_93_WDATA;
            assign ap_WSTRB[93][M_AXIMM_93_DATA_WIDTH/8-1:0] = AP_AXIMM_93_WSTRB;
            assign ap_WLAST[93] = AP_AXIMM_93_WLAST;
            assign ap_WVALID[93] = AP_AXIMM_93_WVALID;
            assign AP_AXIMM_93_WREADY = ap_WREADY[93];
            assign AP_AXIMM_93_BRESP = ap_BRESP[93];
            assign AP_AXIMM_93_BVALID = ap_BVALID[93];
            assign ap_BREADY[93] = AP_AXIMM_93_BREADY;
            assign ap_ARADDR[93][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_93_ARADDR;
            assign ap_ARLEN[93] = AP_AXIMM_93_ARLEN;
            assign ap_ARSIZE[93] = AP_AXIMM_93_ARSIZE;
            assign ap_ARBURST[93] = AP_AXIMM_93_ARBURST;
            assign ap_ARLOCK[93] = AP_AXIMM_93_ARLOCK;
            assign ap_ARCACHE[93] = AP_AXIMM_93_ARCACHE;
            assign ap_ARPROT[93] = AP_AXIMM_93_ARPROT;
            assign ap_ARREGION[93] = AP_AXIMM_93_ARREGION;
            assign ap_ARQOS[93] = AP_AXIMM_93_ARQOS;
            assign ap_ARVALID[93] = AP_AXIMM_93_ARVALID;
            assign AP_AXIMM_93_ARREADY = ap_ARREADY[93];
            assign AP_AXIMM_93_RDATA = ap_RDATA[93][M_AXIMM_93_DATA_WIDTH-1:0];
            assign AP_AXIMM_93_RRESP = ap_RRESP[93];
            assign AP_AXIMM_93_RLAST = ap_RLAST[93];
            assign AP_AXIMM_93_RVALID = ap_RVALID[93];
            assign ap_RREADY[93] = AP_AXIMM_93_RREADY;
            assign M_AXIMM_93_AWADDR = dm_AWADDR[93][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_93_AWLEN = dm_AWLEN[93];
            assign M_AXIMM_93_AWSIZE = dm_AWSIZE[93];
            assign M_AXIMM_93_AWBURST = dm_AWBURST[93];
            assign M_AXIMM_93_AWLOCK = dm_AWLOCK[93];
            assign M_AXIMM_93_AWCACHE = dm_AWCACHE[93];
            assign M_AXIMM_93_AWPROT = dm_AWPROT[93];
            assign M_AXIMM_93_AWREGION = dm_AWREGION[93];
            assign M_AXIMM_93_AWQOS = dm_AWQOS[93];
            assign M_AXIMM_93_AWVALID = dm_AWVALID[93];
            assign dm_AWREADY[93] = M_AXIMM_93_AWREADY;
            assign M_AXIMM_93_WDATA = dm_WDATA[93][M_AXIMM_93_DATA_WIDTH-1:0];
            assign M_AXIMM_93_WSTRB = dm_WSTRB[93][M_AXIMM_93_DATA_WIDTH/8-1:0];
            assign M_AXIMM_93_WLAST = dm_WLAST[93];
            assign M_AXIMM_93_WVALID = dm_WVALID[93];
            assign dm_WREADY[93] = M_AXIMM_93_WREADY;
            assign dm_BRESP[93] = M_AXIMM_93_BRESP;
            assign dm_BVALID[93] = M_AXIMM_93_BVALID;
            assign M_AXIMM_93_BREADY = dm_BREADY[93];
            assign M_AXIMM_93_ARADDR = dm_ARADDR[93][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_93_ARLEN = dm_ARLEN[93];
            assign M_AXIMM_93_ARSIZE = dm_ARSIZE[93];
            assign M_AXIMM_93_ARBURST = dm_ARBURST[93];
            assign M_AXIMM_93_ARLOCK = dm_ARLOCK[93];
            assign M_AXIMM_93_ARCACHE = dm_ARCACHE[93];
            assign M_AXIMM_93_ARPROT = dm_ARPROT[93];
            assign M_AXIMM_93_ARREGION = dm_ARREGION[93];
            assign M_AXIMM_93_ARQOS = dm_ARQOS[93];
            assign M_AXIMM_93_ARVALID = dm_ARVALID[93];
            assign dm_ARREADY[93] = M_AXIMM_93_ARREADY;
            assign dm_RDATA[93][M_AXIMM_93_DATA_WIDTH-1:0] = M_AXIMM_93_RDATA;
            assign dm_RRESP[93] = M_AXIMM_93_RRESP;
            assign dm_RLAST[93] = M_AXIMM_93_RLAST;
            assign dm_RVALID[93] = M_AXIMM_93_RVALID;
            assign M_AXIMM_93_RREADY = dm_RREADY[93];
        end
        if(C_NUM_AXIMMs > 94) begin
            assign ap_AWADDR[94][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_94_AWADDR;
            assign ap_AWLEN[94] = AP_AXIMM_94_AWLEN;
            assign ap_AWSIZE[94] = AP_AXIMM_94_AWSIZE;
            assign ap_AWBURST[94] = AP_AXIMM_94_AWBURST;
            assign ap_AWLOCK[94] = AP_AXIMM_94_AWLOCK;
            assign ap_AWCACHE[94] = AP_AXIMM_94_AWCACHE;
            assign ap_AWPROT[94] = AP_AXIMM_94_AWPROT;
            assign ap_AWREGION[94] = AP_AXIMM_94_AWREGION;
            assign ap_AWQOS[94] = AP_AXIMM_94_AWQOS;
            assign ap_AWVALID[94] = AP_AXIMM_94_AWVALID;
            assign AP_AXIMM_94_AWREADY = ap_AWREADY[94];
            assign ap_WDATA[94][M_AXIMM_94_DATA_WIDTH-1:0] = AP_AXIMM_94_WDATA;
            assign ap_WSTRB[94][M_AXIMM_94_DATA_WIDTH/8-1:0] = AP_AXIMM_94_WSTRB;
            assign ap_WLAST[94] = AP_AXIMM_94_WLAST;
            assign ap_WVALID[94] = AP_AXIMM_94_WVALID;
            assign AP_AXIMM_94_WREADY = ap_WREADY[94];
            assign AP_AXIMM_94_BRESP = ap_BRESP[94];
            assign AP_AXIMM_94_BVALID = ap_BVALID[94];
            assign ap_BREADY[94] = AP_AXIMM_94_BREADY;
            assign ap_ARADDR[94][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_94_ARADDR;
            assign ap_ARLEN[94] = AP_AXIMM_94_ARLEN;
            assign ap_ARSIZE[94] = AP_AXIMM_94_ARSIZE;
            assign ap_ARBURST[94] = AP_AXIMM_94_ARBURST;
            assign ap_ARLOCK[94] = AP_AXIMM_94_ARLOCK;
            assign ap_ARCACHE[94] = AP_AXIMM_94_ARCACHE;
            assign ap_ARPROT[94] = AP_AXIMM_94_ARPROT;
            assign ap_ARREGION[94] = AP_AXIMM_94_ARREGION;
            assign ap_ARQOS[94] = AP_AXIMM_94_ARQOS;
            assign ap_ARVALID[94] = AP_AXIMM_94_ARVALID;
            assign AP_AXIMM_94_ARREADY = ap_ARREADY[94];
            assign AP_AXIMM_94_RDATA = ap_RDATA[94][M_AXIMM_94_DATA_WIDTH-1:0];
            assign AP_AXIMM_94_RRESP = ap_RRESP[94];
            assign AP_AXIMM_94_RLAST = ap_RLAST[94];
            assign AP_AXIMM_94_RVALID = ap_RVALID[94];
            assign ap_RREADY[94] = AP_AXIMM_94_RREADY;
            assign M_AXIMM_94_AWADDR = dm_AWADDR[94][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_94_AWLEN = dm_AWLEN[94];
            assign M_AXIMM_94_AWSIZE = dm_AWSIZE[94];
            assign M_AXIMM_94_AWBURST = dm_AWBURST[94];
            assign M_AXIMM_94_AWLOCK = dm_AWLOCK[94];
            assign M_AXIMM_94_AWCACHE = dm_AWCACHE[94];
            assign M_AXIMM_94_AWPROT = dm_AWPROT[94];
            assign M_AXIMM_94_AWREGION = dm_AWREGION[94];
            assign M_AXIMM_94_AWQOS = dm_AWQOS[94];
            assign M_AXIMM_94_AWVALID = dm_AWVALID[94];
            assign dm_AWREADY[94] = M_AXIMM_94_AWREADY;
            assign M_AXIMM_94_WDATA = dm_WDATA[94][M_AXIMM_94_DATA_WIDTH-1:0];
            assign M_AXIMM_94_WSTRB = dm_WSTRB[94][M_AXIMM_94_DATA_WIDTH/8-1:0];
            assign M_AXIMM_94_WLAST = dm_WLAST[94];
            assign M_AXIMM_94_WVALID = dm_WVALID[94];
            assign dm_WREADY[94] = M_AXIMM_94_WREADY;
            assign dm_BRESP[94] = M_AXIMM_94_BRESP;
            assign dm_BVALID[94] = M_AXIMM_94_BVALID;
            assign M_AXIMM_94_BREADY = dm_BREADY[94];
            assign M_AXIMM_94_ARADDR = dm_ARADDR[94][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_94_ARLEN = dm_ARLEN[94];
            assign M_AXIMM_94_ARSIZE = dm_ARSIZE[94];
            assign M_AXIMM_94_ARBURST = dm_ARBURST[94];
            assign M_AXIMM_94_ARLOCK = dm_ARLOCK[94];
            assign M_AXIMM_94_ARCACHE = dm_ARCACHE[94];
            assign M_AXIMM_94_ARPROT = dm_ARPROT[94];
            assign M_AXIMM_94_ARREGION = dm_ARREGION[94];
            assign M_AXIMM_94_ARQOS = dm_ARQOS[94];
            assign M_AXIMM_94_ARVALID = dm_ARVALID[94];
            assign dm_ARREADY[94] = M_AXIMM_94_ARREADY;
            assign dm_RDATA[94][M_AXIMM_94_DATA_WIDTH-1:0] = M_AXIMM_94_RDATA;
            assign dm_RRESP[94] = M_AXIMM_94_RRESP;
            assign dm_RLAST[94] = M_AXIMM_94_RLAST;
            assign dm_RVALID[94] = M_AXIMM_94_RVALID;
            assign M_AXIMM_94_RREADY = dm_RREADY[94];
        end
        if(C_NUM_AXIMMs > 95) begin
            assign ap_AWADDR[95][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_95_AWADDR;
            assign ap_AWLEN[95] = AP_AXIMM_95_AWLEN;
            assign ap_AWSIZE[95] = AP_AXIMM_95_AWSIZE;
            assign ap_AWBURST[95] = AP_AXIMM_95_AWBURST;
            assign ap_AWLOCK[95] = AP_AXIMM_95_AWLOCK;
            assign ap_AWCACHE[95] = AP_AXIMM_95_AWCACHE;
            assign ap_AWPROT[95] = AP_AXIMM_95_AWPROT;
            assign ap_AWREGION[95] = AP_AXIMM_95_AWREGION;
            assign ap_AWQOS[95] = AP_AXIMM_95_AWQOS;
            assign ap_AWVALID[95] = AP_AXIMM_95_AWVALID;
            assign AP_AXIMM_95_AWREADY = ap_AWREADY[95];
            assign ap_WDATA[95][M_AXIMM_95_DATA_WIDTH-1:0] = AP_AXIMM_95_WDATA;
            assign ap_WSTRB[95][M_AXIMM_95_DATA_WIDTH/8-1:0] = AP_AXIMM_95_WSTRB;
            assign ap_WLAST[95] = AP_AXIMM_95_WLAST;
            assign ap_WVALID[95] = AP_AXIMM_95_WVALID;
            assign AP_AXIMM_95_WREADY = ap_WREADY[95];
            assign AP_AXIMM_95_BRESP = ap_BRESP[95];
            assign AP_AXIMM_95_BVALID = ap_BVALID[95];
            assign ap_BREADY[95] = AP_AXIMM_95_BREADY;
            assign ap_ARADDR[95][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_95_ARADDR;
            assign ap_ARLEN[95] = AP_AXIMM_95_ARLEN;
            assign ap_ARSIZE[95] = AP_AXIMM_95_ARSIZE;
            assign ap_ARBURST[95] = AP_AXIMM_95_ARBURST;
            assign ap_ARLOCK[95] = AP_AXIMM_95_ARLOCK;
            assign ap_ARCACHE[95] = AP_AXIMM_95_ARCACHE;
            assign ap_ARPROT[95] = AP_AXIMM_95_ARPROT;
            assign ap_ARREGION[95] = AP_AXIMM_95_ARREGION;
            assign ap_ARQOS[95] = AP_AXIMM_95_ARQOS;
            assign ap_ARVALID[95] = AP_AXIMM_95_ARVALID;
            assign AP_AXIMM_95_ARREADY = ap_ARREADY[95];
            assign AP_AXIMM_95_RDATA = ap_RDATA[95][M_AXIMM_95_DATA_WIDTH-1:0];
            assign AP_AXIMM_95_RRESP = ap_RRESP[95];
            assign AP_AXIMM_95_RLAST = ap_RLAST[95];
            assign AP_AXIMM_95_RVALID = ap_RVALID[95];
            assign ap_RREADY[95] = AP_AXIMM_95_RREADY;
            assign M_AXIMM_95_AWADDR = dm_AWADDR[95][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_95_AWLEN = dm_AWLEN[95];
            assign M_AXIMM_95_AWSIZE = dm_AWSIZE[95];
            assign M_AXIMM_95_AWBURST = dm_AWBURST[95];
            assign M_AXIMM_95_AWLOCK = dm_AWLOCK[95];
            assign M_AXIMM_95_AWCACHE = dm_AWCACHE[95];
            assign M_AXIMM_95_AWPROT = dm_AWPROT[95];
            assign M_AXIMM_95_AWREGION = dm_AWREGION[95];
            assign M_AXIMM_95_AWQOS = dm_AWQOS[95];
            assign M_AXIMM_95_AWVALID = dm_AWVALID[95];
            assign dm_AWREADY[95] = M_AXIMM_95_AWREADY;
            assign M_AXIMM_95_WDATA = dm_WDATA[95][M_AXIMM_95_DATA_WIDTH-1:0];
            assign M_AXIMM_95_WSTRB = dm_WSTRB[95][M_AXIMM_95_DATA_WIDTH/8-1:0];
            assign M_AXIMM_95_WLAST = dm_WLAST[95];
            assign M_AXIMM_95_WVALID = dm_WVALID[95];
            assign dm_WREADY[95] = M_AXIMM_95_WREADY;
            assign dm_BRESP[95] = M_AXIMM_95_BRESP;
            assign dm_BVALID[95] = M_AXIMM_95_BVALID;
            assign M_AXIMM_95_BREADY = dm_BREADY[95];
            assign M_AXIMM_95_ARADDR = dm_ARADDR[95][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_95_ARLEN = dm_ARLEN[95];
            assign M_AXIMM_95_ARSIZE = dm_ARSIZE[95];
            assign M_AXIMM_95_ARBURST = dm_ARBURST[95];
            assign M_AXIMM_95_ARLOCK = dm_ARLOCK[95];
            assign M_AXIMM_95_ARCACHE = dm_ARCACHE[95];
            assign M_AXIMM_95_ARPROT = dm_ARPROT[95];
            assign M_AXIMM_95_ARREGION = dm_ARREGION[95];
            assign M_AXIMM_95_ARQOS = dm_ARQOS[95];
            assign M_AXIMM_95_ARVALID = dm_ARVALID[95];
            assign dm_ARREADY[95] = M_AXIMM_95_ARREADY;
            assign dm_RDATA[95][M_AXIMM_95_DATA_WIDTH-1:0] = M_AXIMM_95_RDATA;
            assign dm_RRESP[95] = M_AXIMM_95_RRESP;
            assign dm_RLAST[95] = M_AXIMM_95_RLAST;
            assign dm_RVALID[95] = M_AXIMM_95_RVALID;
            assign M_AXIMM_95_RREADY = dm_RREADY[95];
        end
        if(C_NUM_AXIMMs > 96) begin
            assign ap_AWADDR[96][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_96_AWADDR;
            assign ap_AWLEN[96] = AP_AXIMM_96_AWLEN;
            assign ap_AWSIZE[96] = AP_AXIMM_96_AWSIZE;
            assign ap_AWBURST[96] = AP_AXIMM_96_AWBURST;
            assign ap_AWLOCK[96] = AP_AXIMM_96_AWLOCK;
            assign ap_AWCACHE[96] = AP_AXIMM_96_AWCACHE;
            assign ap_AWPROT[96] = AP_AXIMM_96_AWPROT;
            assign ap_AWREGION[96] = AP_AXIMM_96_AWREGION;
            assign ap_AWQOS[96] = AP_AXIMM_96_AWQOS;
            assign ap_AWVALID[96] = AP_AXIMM_96_AWVALID;
            assign AP_AXIMM_96_AWREADY = ap_AWREADY[96];
            assign ap_WDATA[96][M_AXIMM_96_DATA_WIDTH-1:0] = AP_AXIMM_96_WDATA;
            assign ap_WSTRB[96][M_AXIMM_96_DATA_WIDTH/8-1:0] = AP_AXIMM_96_WSTRB;
            assign ap_WLAST[96] = AP_AXIMM_96_WLAST;
            assign ap_WVALID[96] = AP_AXIMM_96_WVALID;
            assign AP_AXIMM_96_WREADY = ap_WREADY[96];
            assign AP_AXIMM_96_BRESP = ap_BRESP[96];
            assign AP_AXIMM_96_BVALID = ap_BVALID[96];
            assign ap_BREADY[96] = AP_AXIMM_96_BREADY;
            assign ap_ARADDR[96][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_96_ARADDR;
            assign ap_ARLEN[96] = AP_AXIMM_96_ARLEN;
            assign ap_ARSIZE[96] = AP_AXIMM_96_ARSIZE;
            assign ap_ARBURST[96] = AP_AXIMM_96_ARBURST;
            assign ap_ARLOCK[96] = AP_AXIMM_96_ARLOCK;
            assign ap_ARCACHE[96] = AP_AXIMM_96_ARCACHE;
            assign ap_ARPROT[96] = AP_AXIMM_96_ARPROT;
            assign ap_ARREGION[96] = AP_AXIMM_96_ARREGION;
            assign ap_ARQOS[96] = AP_AXIMM_96_ARQOS;
            assign ap_ARVALID[96] = AP_AXIMM_96_ARVALID;
            assign AP_AXIMM_96_ARREADY = ap_ARREADY[96];
            assign AP_AXIMM_96_RDATA = ap_RDATA[96][M_AXIMM_96_DATA_WIDTH-1:0];
            assign AP_AXIMM_96_RRESP = ap_RRESP[96];
            assign AP_AXIMM_96_RLAST = ap_RLAST[96];
            assign AP_AXIMM_96_RVALID = ap_RVALID[96];
            assign ap_RREADY[96] = AP_AXIMM_96_RREADY;
            assign M_AXIMM_96_AWADDR = dm_AWADDR[96][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_96_AWLEN = dm_AWLEN[96];
            assign M_AXIMM_96_AWSIZE = dm_AWSIZE[96];
            assign M_AXIMM_96_AWBURST = dm_AWBURST[96];
            assign M_AXIMM_96_AWLOCK = dm_AWLOCK[96];
            assign M_AXIMM_96_AWCACHE = dm_AWCACHE[96];
            assign M_AXIMM_96_AWPROT = dm_AWPROT[96];
            assign M_AXIMM_96_AWREGION = dm_AWREGION[96];
            assign M_AXIMM_96_AWQOS = dm_AWQOS[96];
            assign M_AXIMM_96_AWVALID = dm_AWVALID[96];
            assign dm_AWREADY[96] = M_AXIMM_96_AWREADY;
            assign M_AXIMM_96_WDATA = dm_WDATA[96][M_AXIMM_96_DATA_WIDTH-1:0];
            assign M_AXIMM_96_WSTRB = dm_WSTRB[96][M_AXIMM_96_DATA_WIDTH/8-1:0];
            assign M_AXIMM_96_WLAST = dm_WLAST[96];
            assign M_AXIMM_96_WVALID = dm_WVALID[96];
            assign dm_WREADY[96] = M_AXIMM_96_WREADY;
            assign dm_BRESP[96] = M_AXIMM_96_BRESP;
            assign dm_BVALID[96] = M_AXIMM_96_BVALID;
            assign M_AXIMM_96_BREADY = dm_BREADY[96];
            assign M_AXIMM_96_ARADDR = dm_ARADDR[96][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_96_ARLEN = dm_ARLEN[96];
            assign M_AXIMM_96_ARSIZE = dm_ARSIZE[96];
            assign M_AXIMM_96_ARBURST = dm_ARBURST[96];
            assign M_AXIMM_96_ARLOCK = dm_ARLOCK[96];
            assign M_AXIMM_96_ARCACHE = dm_ARCACHE[96];
            assign M_AXIMM_96_ARPROT = dm_ARPROT[96];
            assign M_AXIMM_96_ARREGION = dm_ARREGION[96];
            assign M_AXIMM_96_ARQOS = dm_ARQOS[96];
            assign M_AXIMM_96_ARVALID = dm_ARVALID[96];
            assign dm_ARREADY[96] = M_AXIMM_96_ARREADY;
            assign dm_RDATA[96][M_AXIMM_96_DATA_WIDTH-1:0] = M_AXIMM_96_RDATA;
            assign dm_RRESP[96] = M_AXIMM_96_RRESP;
            assign dm_RLAST[96] = M_AXIMM_96_RLAST;
            assign dm_RVALID[96] = M_AXIMM_96_RVALID;
            assign M_AXIMM_96_RREADY = dm_RREADY[96];
        end
        if(C_NUM_AXIMMs > 97) begin
            assign ap_AWADDR[97][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_97_AWADDR;
            assign ap_AWLEN[97] = AP_AXIMM_97_AWLEN;
            assign ap_AWSIZE[97] = AP_AXIMM_97_AWSIZE;
            assign ap_AWBURST[97] = AP_AXIMM_97_AWBURST;
            assign ap_AWLOCK[97] = AP_AXIMM_97_AWLOCK;
            assign ap_AWCACHE[97] = AP_AXIMM_97_AWCACHE;
            assign ap_AWPROT[97] = AP_AXIMM_97_AWPROT;
            assign ap_AWREGION[97] = AP_AXIMM_97_AWREGION;
            assign ap_AWQOS[97] = AP_AXIMM_97_AWQOS;
            assign ap_AWVALID[97] = AP_AXIMM_97_AWVALID;
            assign AP_AXIMM_97_AWREADY = ap_AWREADY[97];
            assign ap_WDATA[97][M_AXIMM_97_DATA_WIDTH-1:0] = AP_AXIMM_97_WDATA;
            assign ap_WSTRB[97][M_AXIMM_97_DATA_WIDTH/8-1:0] = AP_AXIMM_97_WSTRB;
            assign ap_WLAST[97] = AP_AXIMM_97_WLAST;
            assign ap_WVALID[97] = AP_AXIMM_97_WVALID;
            assign AP_AXIMM_97_WREADY = ap_WREADY[97];
            assign AP_AXIMM_97_BRESP = ap_BRESP[97];
            assign AP_AXIMM_97_BVALID = ap_BVALID[97];
            assign ap_BREADY[97] = AP_AXIMM_97_BREADY;
            assign ap_ARADDR[97][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_97_ARADDR;
            assign ap_ARLEN[97] = AP_AXIMM_97_ARLEN;
            assign ap_ARSIZE[97] = AP_AXIMM_97_ARSIZE;
            assign ap_ARBURST[97] = AP_AXIMM_97_ARBURST;
            assign ap_ARLOCK[97] = AP_AXIMM_97_ARLOCK;
            assign ap_ARCACHE[97] = AP_AXIMM_97_ARCACHE;
            assign ap_ARPROT[97] = AP_AXIMM_97_ARPROT;
            assign ap_ARREGION[97] = AP_AXIMM_97_ARREGION;
            assign ap_ARQOS[97] = AP_AXIMM_97_ARQOS;
            assign ap_ARVALID[97] = AP_AXIMM_97_ARVALID;
            assign AP_AXIMM_97_ARREADY = ap_ARREADY[97];
            assign AP_AXIMM_97_RDATA = ap_RDATA[97][M_AXIMM_97_DATA_WIDTH-1:0];
            assign AP_AXIMM_97_RRESP = ap_RRESP[97];
            assign AP_AXIMM_97_RLAST = ap_RLAST[97];
            assign AP_AXIMM_97_RVALID = ap_RVALID[97];
            assign ap_RREADY[97] = AP_AXIMM_97_RREADY;
            assign M_AXIMM_97_AWADDR = dm_AWADDR[97][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_97_AWLEN = dm_AWLEN[97];
            assign M_AXIMM_97_AWSIZE = dm_AWSIZE[97];
            assign M_AXIMM_97_AWBURST = dm_AWBURST[97];
            assign M_AXIMM_97_AWLOCK = dm_AWLOCK[97];
            assign M_AXIMM_97_AWCACHE = dm_AWCACHE[97];
            assign M_AXIMM_97_AWPROT = dm_AWPROT[97];
            assign M_AXIMM_97_AWREGION = dm_AWREGION[97];
            assign M_AXIMM_97_AWQOS = dm_AWQOS[97];
            assign M_AXIMM_97_AWVALID = dm_AWVALID[97];
            assign dm_AWREADY[97] = M_AXIMM_97_AWREADY;
            assign M_AXIMM_97_WDATA = dm_WDATA[97][M_AXIMM_97_DATA_WIDTH-1:0];
            assign M_AXIMM_97_WSTRB = dm_WSTRB[97][M_AXIMM_97_DATA_WIDTH/8-1:0];
            assign M_AXIMM_97_WLAST = dm_WLAST[97];
            assign M_AXIMM_97_WVALID = dm_WVALID[97];
            assign dm_WREADY[97] = M_AXIMM_97_WREADY;
            assign dm_BRESP[97] = M_AXIMM_97_BRESP;
            assign dm_BVALID[97] = M_AXIMM_97_BVALID;
            assign M_AXIMM_97_BREADY = dm_BREADY[97];
            assign M_AXIMM_97_ARADDR = dm_ARADDR[97][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_97_ARLEN = dm_ARLEN[97];
            assign M_AXIMM_97_ARSIZE = dm_ARSIZE[97];
            assign M_AXIMM_97_ARBURST = dm_ARBURST[97];
            assign M_AXIMM_97_ARLOCK = dm_ARLOCK[97];
            assign M_AXIMM_97_ARCACHE = dm_ARCACHE[97];
            assign M_AXIMM_97_ARPROT = dm_ARPROT[97];
            assign M_AXIMM_97_ARREGION = dm_ARREGION[97];
            assign M_AXIMM_97_ARQOS = dm_ARQOS[97];
            assign M_AXIMM_97_ARVALID = dm_ARVALID[97];
            assign dm_ARREADY[97] = M_AXIMM_97_ARREADY;
            assign dm_RDATA[97][M_AXIMM_97_DATA_WIDTH-1:0] = M_AXIMM_97_RDATA;
            assign dm_RRESP[97] = M_AXIMM_97_RRESP;
            assign dm_RLAST[97] = M_AXIMM_97_RLAST;
            assign dm_RVALID[97] = M_AXIMM_97_RVALID;
            assign M_AXIMM_97_RREADY = dm_RREADY[97];
        end
        if(C_NUM_AXIMMs > 98) begin
            assign ap_AWADDR[98][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_98_AWADDR;
            assign ap_AWLEN[98] = AP_AXIMM_98_AWLEN;
            assign ap_AWSIZE[98] = AP_AXIMM_98_AWSIZE;
            assign ap_AWBURST[98] = AP_AXIMM_98_AWBURST;
            assign ap_AWLOCK[98] = AP_AXIMM_98_AWLOCK;
            assign ap_AWCACHE[98] = AP_AXIMM_98_AWCACHE;
            assign ap_AWPROT[98] = AP_AXIMM_98_AWPROT;
            assign ap_AWREGION[98] = AP_AXIMM_98_AWREGION;
            assign ap_AWQOS[98] = AP_AXIMM_98_AWQOS;
            assign ap_AWVALID[98] = AP_AXIMM_98_AWVALID;
            assign AP_AXIMM_98_AWREADY = ap_AWREADY[98];
            assign ap_WDATA[98][M_AXIMM_98_DATA_WIDTH-1:0] = AP_AXIMM_98_WDATA;
            assign ap_WSTRB[98][M_AXIMM_98_DATA_WIDTH/8-1:0] = AP_AXIMM_98_WSTRB;
            assign ap_WLAST[98] = AP_AXIMM_98_WLAST;
            assign ap_WVALID[98] = AP_AXIMM_98_WVALID;
            assign AP_AXIMM_98_WREADY = ap_WREADY[98];
            assign AP_AXIMM_98_BRESP = ap_BRESP[98];
            assign AP_AXIMM_98_BVALID = ap_BVALID[98];
            assign ap_BREADY[98] = AP_AXIMM_98_BREADY;
            assign ap_ARADDR[98][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_98_ARADDR;
            assign ap_ARLEN[98] = AP_AXIMM_98_ARLEN;
            assign ap_ARSIZE[98] = AP_AXIMM_98_ARSIZE;
            assign ap_ARBURST[98] = AP_AXIMM_98_ARBURST;
            assign ap_ARLOCK[98] = AP_AXIMM_98_ARLOCK;
            assign ap_ARCACHE[98] = AP_AXIMM_98_ARCACHE;
            assign ap_ARPROT[98] = AP_AXIMM_98_ARPROT;
            assign ap_ARREGION[98] = AP_AXIMM_98_ARREGION;
            assign ap_ARQOS[98] = AP_AXIMM_98_ARQOS;
            assign ap_ARVALID[98] = AP_AXIMM_98_ARVALID;
            assign AP_AXIMM_98_ARREADY = ap_ARREADY[98];
            assign AP_AXIMM_98_RDATA = ap_RDATA[98][M_AXIMM_98_DATA_WIDTH-1:0];
            assign AP_AXIMM_98_RRESP = ap_RRESP[98];
            assign AP_AXIMM_98_RLAST = ap_RLAST[98];
            assign AP_AXIMM_98_RVALID = ap_RVALID[98];
            assign ap_RREADY[98] = AP_AXIMM_98_RREADY;
            assign M_AXIMM_98_AWADDR = dm_AWADDR[98][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_98_AWLEN = dm_AWLEN[98];
            assign M_AXIMM_98_AWSIZE = dm_AWSIZE[98];
            assign M_AXIMM_98_AWBURST = dm_AWBURST[98];
            assign M_AXIMM_98_AWLOCK = dm_AWLOCK[98];
            assign M_AXIMM_98_AWCACHE = dm_AWCACHE[98];
            assign M_AXIMM_98_AWPROT = dm_AWPROT[98];
            assign M_AXIMM_98_AWREGION = dm_AWREGION[98];
            assign M_AXIMM_98_AWQOS = dm_AWQOS[98];
            assign M_AXIMM_98_AWVALID = dm_AWVALID[98];
            assign dm_AWREADY[98] = M_AXIMM_98_AWREADY;
            assign M_AXIMM_98_WDATA = dm_WDATA[98][M_AXIMM_98_DATA_WIDTH-1:0];
            assign M_AXIMM_98_WSTRB = dm_WSTRB[98][M_AXIMM_98_DATA_WIDTH/8-1:0];
            assign M_AXIMM_98_WLAST = dm_WLAST[98];
            assign M_AXIMM_98_WVALID = dm_WVALID[98];
            assign dm_WREADY[98] = M_AXIMM_98_WREADY;
            assign dm_BRESP[98] = M_AXIMM_98_BRESP;
            assign dm_BVALID[98] = M_AXIMM_98_BVALID;
            assign M_AXIMM_98_BREADY = dm_BREADY[98];
            assign M_AXIMM_98_ARADDR = dm_ARADDR[98][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_98_ARLEN = dm_ARLEN[98];
            assign M_AXIMM_98_ARSIZE = dm_ARSIZE[98];
            assign M_AXIMM_98_ARBURST = dm_ARBURST[98];
            assign M_AXIMM_98_ARLOCK = dm_ARLOCK[98];
            assign M_AXIMM_98_ARCACHE = dm_ARCACHE[98];
            assign M_AXIMM_98_ARPROT = dm_ARPROT[98];
            assign M_AXIMM_98_ARREGION = dm_ARREGION[98];
            assign M_AXIMM_98_ARQOS = dm_ARQOS[98];
            assign M_AXIMM_98_ARVALID = dm_ARVALID[98];
            assign dm_ARREADY[98] = M_AXIMM_98_ARREADY;
            assign dm_RDATA[98][M_AXIMM_98_DATA_WIDTH-1:0] = M_AXIMM_98_RDATA;
            assign dm_RRESP[98] = M_AXIMM_98_RRESP;
            assign dm_RLAST[98] = M_AXIMM_98_RLAST;
            assign dm_RVALID[98] = M_AXIMM_98_RVALID;
            assign M_AXIMM_98_RREADY = dm_RREADY[98];
        end
        if(C_NUM_AXIMMs > 99) begin
            assign ap_AWADDR[99][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_99_AWADDR;
            assign ap_AWLEN[99] = AP_AXIMM_99_AWLEN;
            assign ap_AWSIZE[99] = AP_AXIMM_99_AWSIZE;
            assign ap_AWBURST[99] = AP_AXIMM_99_AWBURST;
            assign ap_AWLOCK[99] = AP_AXIMM_99_AWLOCK;
            assign ap_AWCACHE[99] = AP_AXIMM_99_AWCACHE;
            assign ap_AWPROT[99] = AP_AXIMM_99_AWPROT;
            assign ap_AWREGION[99] = AP_AXIMM_99_AWREGION;
            assign ap_AWQOS[99] = AP_AXIMM_99_AWQOS;
            assign ap_AWVALID[99] = AP_AXIMM_99_AWVALID;
            assign AP_AXIMM_99_AWREADY = ap_AWREADY[99];
            assign ap_WDATA[99][M_AXIMM_99_DATA_WIDTH-1:0] = AP_AXIMM_99_WDATA;
            assign ap_WSTRB[99][M_AXIMM_99_DATA_WIDTH/8-1:0] = AP_AXIMM_99_WSTRB;
            assign ap_WLAST[99] = AP_AXIMM_99_WLAST;
            assign ap_WVALID[99] = AP_AXIMM_99_WVALID;
            assign AP_AXIMM_99_WREADY = ap_WREADY[99];
            assign AP_AXIMM_99_BRESP = ap_BRESP[99];
            assign AP_AXIMM_99_BVALID = ap_BVALID[99];
            assign ap_BREADY[99] = AP_AXIMM_99_BREADY;
            assign ap_ARADDR[99][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_99_ARADDR;
            assign ap_ARLEN[99] = AP_AXIMM_99_ARLEN;
            assign ap_ARSIZE[99] = AP_AXIMM_99_ARSIZE;
            assign ap_ARBURST[99] = AP_AXIMM_99_ARBURST;
            assign ap_ARLOCK[99] = AP_AXIMM_99_ARLOCK;
            assign ap_ARCACHE[99] = AP_AXIMM_99_ARCACHE;
            assign ap_ARPROT[99] = AP_AXIMM_99_ARPROT;
            assign ap_ARREGION[99] = AP_AXIMM_99_ARREGION;
            assign ap_ARQOS[99] = AP_AXIMM_99_ARQOS;
            assign ap_ARVALID[99] = AP_AXIMM_99_ARVALID;
            assign AP_AXIMM_99_ARREADY = ap_ARREADY[99];
            assign AP_AXIMM_99_RDATA = ap_RDATA[99][M_AXIMM_99_DATA_WIDTH-1:0];
            assign AP_AXIMM_99_RRESP = ap_RRESP[99];
            assign AP_AXIMM_99_RLAST = ap_RLAST[99];
            assign AP_AXIMM_99_RVALID = ap_RVALID[99];
            assign ap_RREADY[99] = AP_AXIMM_99_RREADY;
            assign M_AXIMM_99_AWADDR = dm_AWADDR[99][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_99_AWLEN = dm_AWLEN[99];
            assign M_AXIMM_99_AWSIZE = dm_AWSIZE[99];
            assign M_AXIMM_99_AWBURST = dm_AWBURST[99];
            assign M_AXIMM_99_AWLOCK = dm_AWLOCK[99];
            assign M_AXIMM_99_AWCACHE = dm_AWCACHE[99];
            assign M_AXIMM_99_AWPROT = dm_AWPROT[99];
            assign M_AXIMM_99_AWREGION = dm_AWREGION[99];
            assign M_AXIMM_99_AWQOS = dm_AWQOS[99];
            assign M_AXIMM_99_AWVALID = dm_AWVALID[99];
            assign dm_AWREADY[99] = M_AXIMM_99_AWREADY;
            assign M_AXIMM_99_WDATA = dm_WDATA[99][M_AXIMM_99_DATA_WIDTH-1:0];
            assign M_AXIMM_99_WSTRB = dm_WSTRB[99][M_AXIMM_99_DATA_WIDTH/8-1:0];
            assign M_AXIMM_99_WLAST = dm_WLAST[99];
            assign M_AXIMM_99_WVALID = dm_WVALID[99];
            assign dm_WREADY[99] = M_AXIMM_99_WREADY;
            assign dm_BRESP[99] = M_AXIMM_99_BRESP;
            assign dm_BVALID[99] = M_AXIMM_99_BVALID;
            assign M_AXIMM_99_BREADY = dm_BREADY[99];
            assign M_AXIMM_99_ARADDR = dm_ARADDR[99][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_99_ARLEN = dm_ARLEN[99];
            assign M_AXIMM_99_ARSIZE = dm_ARSIZE[99];
            assign M_AXIMM_99_ARBURST = dm_ARBURST[99];
            assign M_AXIMM_99_ARLOCK = dm_ARLOCK[99];
            assign M_AXIMM_99_ARCACHE = dm_ARCACHE[99];
            assign M_AXIMM_99_ARPROT = dm_ARPROT[99];
            assign M_AXIMM_99_ARREGION = dm_ARREGION[99];
            assign M_AXIMM_99_ARQOS = dm_ARQOS[99];
            assign M_AXIMM_99_ARVALID = dm_ARVALID[99];
            assign dm_ARREADY[99] = M_AXIMM_99_ARREADY;
            assign dm_RDATA[99][M_AXIMM_99_DATA_WIDTH-1:0] = M_AXIMM_99_RDATA;
            assign dm_RRESP[99] = M_AXIMM_99_RRESP;
            assign dm_RLAST[99] = M_AXIMM_99_RLAST;
            assign dm_RVALID[99] = M_AXIMM_99_RVALID;
            assign M_AXIMM_99_RREADY = dm_RREADY[99];
        end
        if(C_NUM_AXIMMs > 100) begin
            assign ap_AWADDR[100][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_100_AWADDR;
            assign ap_AWLEN[100] = AP_AXIMM_100_AWLEN;
            assign ap_AWSIZE[100] = AP_AXIMM_100_AWSIZE;
            assign ap_AWBURST[100] = AP_AXIMM_100_AWBURST;
            assign ap_AWLOCK[100] = AP_AXIMM_100_AWLOCK;
            assign ap_AWCACHE[100] = AP_AXIMM_100_AWCACHE;
            assign ap_AWPROT[100] = AP_AXIMM_100_AWPROT;
            assign ap_AWREGION[100] = AP_AXIMM_100_AWREGION;
            assign ap_AWQOS[100] = AP_AXIMM_100_AWQOS;
            assign ap_AWVALID[100] = AP_AXIMM_100_AWVALID;
            assign AP_AXIMM_100_AWREADY = ap_AWREADY[100];
            assign ap_WDATA[100][M_AXIMM_100_DATA_WIDTH-1:0] = AP_AXIMM_100_WDATA;
            assign ap_WSTRB[100][M_AXIMM_100_DATA_WIDTH/8-1:0] = AP_AXIMM_100_WSTRB;
            assign ap_WLAST[100] = AP_AXIMM_100_WLAST;
            assign ap_WVALID[100] = AP_AXIMM_100_WVALID;
            assign AP_AXIMM_100_WREADY = ap_WREADY[100];
            assign AP_AXIMM_100_BRESP = ap_BRESP[100];
            assign AP_AXIMM_100_BVALID = ap_BVALID[100];
            assign ap_BREADY[100] = AP_AXIMM_100_BREADY;
            assign ap_ARADDR[100][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_100_ARADDR;
            assign ap_ARLEN[100] = AP_AXIMM_100_ARLEN;
            assign ap_ARSIZE[100] = AP_AXIMM_100_ARSIZE;
            assign ap_ARBURST[100] = AP_AXIMM_100_ARBURST;
            assign ap_ARLOCK[100] = AP_AXIMM_100_ARLOCK;
            assign ap_ARCACHE[100] = AP_AXIMM_100_ARCACHE;
            assign ap_ARPROT[100] = AP_AXIMM_100_ARPROT;
            assign ap_ARREGION[100] = AP_AXIMM_100_ARREGION;
            assign ap_ARQOS[100] = AP_AXIMM_100_ARQOS;
            assign ap_ARVALID[100] = AP_AXIMM_100_ARVALID;
            assign AP_AXIMM_100_ARREADY = ap_ARREADY[100];
            assign AP_AXIMM_100_RDATA = ap_RDATA[100][M_AXIMM_100_DATA_WIDTH-1:0];
            assign AP_AXIMM_100_RRESP = ap_RRESP[100];
            assign AP_AXIMM_100_RLAST = ap_RLAST[100];
            assign AP_AXIMM_100_RVALID = ap_RVALID[100];
            assign ap_RREADY[100] = AP_AXIMM_100_RREADY;
            assign M_AXIMM_100_AWADDR = dm_AWADDR[100][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_100_AWLEN = dm_AWLEN[100];
            assign M_AXIMM_100_AWSIZE = dm_AWSIZE[100];
            assign M_AXIMM_100_AWBURST = dm_AWBURST[100];
            assign M_AXIMM_100_AWLOCK = dm_AWLOCK[100];
            assign M_AXIMM_100_AWCACHE = dm_AWCACHE[100];
            assign M_AXIMM_100_AWPROT = dm_AWPROT[100];
            assign M_AXIMM_100_AWREGION = dm_AWREGION[100];
            assign M_AXIMM_100_AWQOS = dm_AWQOS[100];
            assign M_AXIMM_100_AWVALID = dm_AWVALID[100];
            assign dm_AWREADY[100] = M_AXIMM_100_AWREADY;
            assign M_AXIMM_100_WDATA = dm_WDATA[100][M_AXIMM_100_DATA_WIDTH-1:0];
            assign M_AXIMM_100_WSTRB = dm_WSTRB[100][M_AXIMM_100_DATA_WIDTH/8-1:0];
            assign M_AXIMM_100_WLAST = dm_WLAST[100];
            assign M_AXIMM_100_WVALID = dm_WVALID[100];
            assign dm_WREADY[100] = M_AXIMM_100_WREADY;
            assign dm_BRESP[100] = M_AXIMM_100_BRESP;
            assign dm_BVALID[100] = M_AXIMM_100_BVALID;
            assign M_AXIMM_100_BREADY = dm_BREADY[100];
            assign M_AXIMM_100_ARADDR = dm_ARADDR[100][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_100_ARLEN = dm_ARLEN[100];
            assign M_AXIMM_100_ARSIZE = dm_ARSIZE[100];
            assign M_AXIMM_100_ARBURST = dm_ARBURST[100];
            assign M_AXIMM_100_ARLOCK = dm_ARLOCK[100];
            assign M_AXIMM_100_ARCACHE = dm_ARCACHE[100];
            assign M_AXIMM_100_ARPROT = dm_ARPROT[100];
            assign M_AXIMM_100_ARREGION = dm_ARREGION[100];
            assign M_AXIMM_100_ARQOS = dm_ARQOS[100];
            assign M_AXIMM_100_ARVALID = dm_ARVALID[100];
            assign dm_ARREADY[100] = M_AXIMM_100_ARREADY;
            assign dm_RDATA[100][M_AXIMM_100_DATA_WIDTH-1:0] = M_AXIMM_100_RDATA;
            assign dm_RRESP[100] = M_AXIMM_100_RRESP;
            assign dm_RLAST[100] = M_AXIMM_100_RLAST;
            assign dm_RVALID[100] = M_AXIMM_100_RVALID;
            assign M_AXIMM_100_RREADY = dm_RREADY[100];
        end
        if(C_NUM_AXIMMs > 101) begin
            assign ap_AWADDR[101][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_101_AWADDR;
            assign ap_AWLEN[101] = AP_AXIMM_101_AWLEN;
            assign ap_AWSIZE[101] = AP_AXIMM_101_AWSIZE;
            assign ap_AWBURST[101] = AP_AXIMM_101_AWBURST;
            assign ap_AWLOCK[101] = AP_AXIMM_101_AWLOCK;
            assign ap_AWCACHE[101] = AP_AXIMM_101_AWCACHE;
            assign ap_AWPROT[101] = AP_AXIMM_101_AWPROT;
            assign ap_AWREGION[101] = AP_AXIMM_101_AWREGION;
            assign ap_AWQOS[101] = AP_AXIMM_101_AWQOS;
            assign ap_AWVALID[101] = AP_AXIMM_101_AWVALID;
            assign AP_AXIMM_101_AWREADY = ap_AWREADY[101];
            assign ap_WDATA[101][M_AXIMM_101_DATA_WIDTH-1:0] = AP_AXIMM_101_WDATA;
            assign ap_WSTRB[101][M_AXIMM_101_DATA_WIDTH/8-1:0] = AP_AXIMM_101_WSTRB;
            assign ap_WLAST[101] = AP_AXIMM_101_WLAST;
            assign ap_WVALID[101] = AP_AXIMM_101_WVALID;
            assign AP_AXIMM_101_WREADY = ap_WREADY[101];
            assign AP_AXIMM_101_BRESP = ap_BRESP[101];
            assign AP_AXIMM_101_BVALID = ap_BVALID[101];
            assign ap_BREADY[101] = AP_AXIMM_101_BREADY;
            assign ap_ARADDR[101][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_101_ARADDR;
            assign ap_ARLEN[101] = AP_AXIMM_101_ARLEN;
            assign ap_ARSIZE[101] = AP_AXIMM_101_ARSIZE;
            assign ap_ARBURST[101] = AP_AXIMM_101_ARBURST;
            assign ap_ARLOCK[101] = AP_AXIMM_101_ARLOCK;
            assign ap_ARCACHE[101] = AP_AXIMM_101_ARCACHE;
            assign ap_ARPROT[101] = AP_AXIMM_101_ARPROT;
            assign ap_ARREGION[101] = AP_AXIMM_101_ARREGION;
            assign ap_ARQOS[101] = AP_AXIMM_101_ARQOS;
            assign ap_ARVALID[101] = AP_AXIMM_101_ARVALID;
            assign AP_AXIMM_101_ARREADY = ap_ARREADY[101];
            assign AP_AXIMM_101_RDATA = ap_RDATA[101][M_AXIMM_101_DATA_WIDTH-1:0];
            assign AP_AXIMM_101_RRESP = ap_RRESP[101];
            assign AP_AXIMM_101_RLAST = ap_RLAST[101];
            assign AP_AXIMM_101_RVALID = ap_RVALID[101];
            assign ap_RREADY[101] = AP_AXIMM_101_RREADY;
            assign M_AXIMM_101_AWADDR = dm_AWADDR[101][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_101_AWLEN = dm_AWLEN[101];
            assign M_AXIMM_101_AWSIZE = dm_AWSIZE[101];
            assign M_AXIMM_101_AWBURST = dm_AWBURST[101];
            assign M_AXIMM_101_AWLOCK = dm_AWLOCK[101];
            assign M_AXIMM_101_AWCACHE = dm_AWCACHE[101];
            assign M_AXIMM_101_AWPROT = dm_AWPROT[101];
            assign M_AXIMM_101_AWREGION = dm_AWREGION[101];
            assign M_AXIMM_101_AWQOS = dm_AWQOS[101];
            assign M_AXIMM_101_AWVALID = dm_AWVALID[101];
            assign dm_AWREADY[101] = M_AXIMM_101_AWREADY;
            assign M_AXIMM_101_WDATA = dm_WDATA[101][M_AXIMM_101_DATA_WIDTH-1:0];
            assign M_AXIMM_101_WSTRB = dm_WSTRB[101][M_AXIMM_101_DATA_WIDTH/8-1:0];
            assign M_AXIMM_101_WLAST = dm_WLAST[101];
            assign M_AXIMM_101_WVALID = dm_WVALID[101];
            assign dm_WREADY[101] = M_AXIMM_101_WREADY;
            assign dm_BRESP[101] = M_AXIMM_101_BRESP;
            assign dm_BVALID[101] = M_AXIMM_101_BVALID;
            assign M_AXIMM_101_BREADY = dm_BREADY[101];
            assign M_AXIMM_101_ARADDR = dm_ARADDR[101][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_101_ARLEN = dm_ARLEN[101];
            assign M_AXIMM_101_ARSIZE = dm_ARSIZE[101];
            assign M_AXIMM_101_ARBURST = dm_ARBURST[101];
            assign M_AXIMM_101_ARLOCK = dm_ARLOCK[101];
            assign M_AXIMM_101_ARCACHE = dm_ARCACHE[101];
            assign M_AXIMM_101_ARPROT = dm_ARPROT[101];
            assign M_AXIMM_101_ARREGION = dm_ARREGION[101];
            assign M_AXIMM_101_ARQOS = dm_ARQOS[101];
            assign M_AXIMM_101_ARVALID = dm_ARVALID[101];
            assign dm_ARREADY[101] = M_AXIMM_101_ARREADY;
            assign dm_RDATA[101][M_AXIMM_101_DATA_WIDTH-1:0] = M_AXIMM_101_RDATA;
            assign dm_RRESP[101] = M_AXIMM_101_RRESP;
            assign dm_RLAST[101] = M_AXIMM_101_RLAST;
            assign dm_RVALID[101] = M_AXIMM_101_RVALID;
            assign M_AXIMM_101_RREADY = dm_RREADY[101];
        end
        if(C_NUM_AXIMMs > 102) begin
            assign ap_AWADDR[102][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_102_AWADDR;
            assign ap_AWLEN[102] = AP_AXIMM_102_AWLEN;
            assign ap_AWSIZE[102] = AP_AXIMM_102_AWSIZE;
            assign ap_AWBURST[102] = AP_AXIMM_102_AWBURST;
            assign ap_AWLOCK[102] = AP_AXIMM_102_AWLOCK;
            assign ap_AWCACHE[102] = AP_AXIMM_102_AWCACHE;
            assign ap_AWPROT[102] = AP_AXIMM_102_AWPROT;
            assign ap_AWREGION[102] = AP_AXIMM_102_AWREGION;
            assign ap_AWQOS[102] = AP_AXIMM_102_AWQOS;
            assign ap_AWVALID[102] = AP_AXIMM_102_AWVALID;
            assign AP_AXIMM_102_AWREADY = ap_AWREADY[102];
            assign ap_WDATA[102][M_AXIMM_102_DATA_WIDTH-1:0] = AP_AXIMM_102_WDATA;
            assign ap_WSTRB[102][M_AXIMM_102_DATA_WIDTH/8-1:0] = AP_AXIMM_102_WSTRB;
            assign ap_WLAST[102] = AP_AXIMM_102_WLAST;
            assign ap_WVALID[102] = AP_AXIMM_102_WVALID;
            assign AP_AXIMM_102_WREADY = ap_WREADY[102];
            assign AP_AXIMM_102_BRESP = ap_BRESP[102];
            assign AP_AXIMM_102_BVALID = ap_BVALID[102];
            assign ap_BREADY[102] = AP_AXIMM_102_BREADY;
            assign ap_ARADDR[102][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_102_ARADDR;
            assign ap_ARLEN[102] = AP_AXIMM_102_ARLEN;
            assign ap_ARSIZE[102] = AP_AXIMM_102_ARSIZE;
            assign ap_ARBURST[102] = AP_AXIMM_102_ARBURST;
            assign ap_ARLOCK[102] = AP_AXIMM_102_ARLOCK;
            assign ap_ARCACHE[102] = AP_AXIMM_102_ARCACHE;
            assign ap_ARPROT[102] = AP_AXIMM_102_ARPROT;
            assign ap_ARREGION[102] = AP_AXIMM_102_ARREGION;
            assign ap_ARQOS[102] = AP_AXIMM_102_ARQOS;
            assign ap_ARVALID[102] = AP_AXIMM_102_ARVALID;
            assign AP_AXIMM_102_ARREADY = ap_ARREADY[102];
            assign AP_AXIMM_102_RDATA = ap_RDATA[102][M_AXIMM_102_DATA_WIDTH-1:0];
            assign AP_AXIMM_102_RRESP = ap_RRESP[102];
            assign AP_AXIMM_102_RLAST = ap_RLAST[102];
            assign AP_AXIMM_102_RVALID = ap_RVALID[102];
            assign ap_RREADY[102] = AP_AXIMM_102_RREADY;
            assign M_AXIMM_102_AWADDR = dm_AWADDR[102][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_102_AWLEN = dm_AWLEN[102];
            assign M_AXIMM_102_AWSIZE = dm_AWSIZE[102];
            assign M_AXIMM_102_AWBURST = dm_AWBURST[102];
            assign M_AXIMM_102_AWLOCK = dm_AWLOCK[102];
            assign M_AXIMM_102_AWCACHE = dm_AWCACHE[102];
            assign M_AXIMM_102_AWPROT = dm_AWPROT[102];
            assign M_AXIMM_102_AWREGION = dm_AWREGION[102];
            assign M_AXIMM_102_AWQOS = dm_AWQOS[102];
            assign M_AXIMM_102_AWVALID = dm_AWVALID[102];
            assign dm_AWREADY[102] = M_AXIMM_102_AWREADY;
            assign M_AXIMM_102_WDATA = dm_WDATA[102][M_AXIMM_102_DATA_WIDTH-1:0];
            assign M_AXIMM_102_WSTRB = dm_WSTRB[102][M_AXIMM_102_DATA_WIDTH/8-1:0];
            assign M_AXIMM_102_WLAST = dm_WLAST[102];
            assign M_AXIMM_102_WVALID = dm_WVALID[102];
            assign dm_WREADY[102] = M_AXIMM_102_WREADY;
            assign dm_BRESP[102] = M_AXIMM_102_BRESP;
            assign dm_BVALID[102] = M_AXIMM_102_BVALID;
            assign M_AXIMM_102_BREADY = dm_BREADY[102];
            assign M_AXIMM_102_ARADDR = dm_ARADDR[102][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_102_ARLEN = dm_ARLEN[102];
            assign M_AXIMM_102_ARSIZE = dm_ARSIZE[102];
            assign M_AXIMM_102_ARBURST = dm_ARBURST[102];
            assign M_AXIMM_102_ARLOCK = dm_ARLOCK[102];
            assign M_AXIMM_102_ARCACHE = dm_ARCACHE[102];
            assign M_AXIMM_102_ARPROT = dm_ARPROT[102];
            assign M_AXIMM_102_ARREGION = dm_ARREGION[102];
            assign M_AXIMM_102_ARQOS = dm_ARQOS[102];
            assign M_AXIMM_102_ARVALID = dm_ARVALID[102];
            assign dm_ARREADY[102] = M_AXIMM_102_ARREADY;
            assign dm_RDATA[102][M_AXIMM_102_DATA_WIDTH-1:0] = M_AXIMM_102_RDATA;
            assign dm_RRESP[102] = M_AXIMM_102_RRESP;
            assign dm_RLAST[102] = M_AXIMM_102_RLAST;
            assign dm_RVALID[102] = M_AXIMM_102_RVALID;
            assign M_AXIMM_102_RREADY = dm_RREADY[102];
        end
        if(C_NUM_AXIMMs > 103) begin
            assign ap_AWADDR[103][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_103_AWADDR;
            assign ap_AWLEN[103] = AP_AXIMM_103_AWLEN;
            assign ap_AWSIZE[103] = AP_AXIMM_103_AWSIZE;
            assign ap_AWBURST[103] = AP_AXIMM_103_AWBURST;
            assign ap_AWLOCK[103] = AP_AXIMM_103_AWLOCK;
            assign ap_AWCACHE[103] = AP_AXIMM_103_AWCACHE;
            assign ap_AWPROT[103] = AP_AXIMM_103_AWPROT;
            assign ap_AWREGION[103] = AP_AXIMM_103_AWREGION;
            assign ap_AWQOS[103] = AP_AXIMM_103_AWQOS;
            assign ap_AWVALID[103] = AP_AXIMM_103_AWVALID;
            assign AP_AXIMM_103_AWREADY = ap_AWREADY[103];
            assign ap_WDATA[103][M_AXIMM_103_DATA_WIDTH-1:0] = AP_AXIMM_103_WDATA;
            assign ap_WSTRB[103][M_AXIMM_103_DATA_WIDTH/8-1:0] = AP_AXIMM_103_WSTRB;
            assign ap_WLAST[103] = AP_AXIMM_103_WLAST;
            assign ap_WVALID[103] = AP_AXIMM_103_WVALID;
            assign AP_AXIMM_103_WREADY = ap_WREADY[103];
            assign AP_AXIMM_103_BRESP = ap_BRESP[103];
            assign AP_AXIMM_103_BVALID = ap_BVALID[103];
            assign ap_BREADY[103] = AP_AXIMM_103_BREADY;
            assign ap_ARADDR[103][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_103_ARADDR;
            assign ap_ARLEN[103] = AP_AXIMM_103_ARLEN;
            assign ap_ARSIZE[103] = AP_AXIMM_103_ARSIZE;
            assign ap_ARBURST[103] = AP_AXIMM_103_ARBURST;
            assign ap_ARLOCK[103] = AP_AXIMM_103_ARLOCK;
            assign ap_ARCACHE[103] = AP_AXIMM_103_ARCACHE;
            assign ap_ARPROT[103] = AP_AXIMM_103_ARPROT;
            assign ap_ARREGION[103] = AP_AXIMM_103_ARREGION;
            assign ap_ARQOS[103] = AP_AXIMM_103_ARQOS;
            assign ap_ARVALID[103] = AP_AXIMM_103_ARVALID;
            assign AP_AXIMM_103_ARREADY = ap_ARREADY[103];
            assign AP_AXIMM_103_RDATA = ap_RDATA[103][M_AXIMM_103_DATA_WIDTH-1:0];
            assign AP_AXIMM_103_RRESP = ap_RRESP[103];
            assign AP_AXIMM_103_RLAST = ap_RLAST[103];
            assign AP_AXIMM_103_RVALID = ap_RVALID[103];
            assign ap_RREADY[103] = AP_AXIMM_103_RREADY;
            assign M_AXIMM_103_AWADDR = dm_AWADDR[103][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_103_AWLEN = dm_AWLEN[103];
            assign M_AXIMM_103_AWSIZE = dm_AWSIZE[103];
            assign M_AXIMM_103_AWBURST = dm_AWBURST[103];
            assign M_AXIMM_103_AWLOCK = dm_AWLOCK[103];
            assign M_AXIMM_103_AWCACHE = dm_AWCACHE[103];
            assign M_AXIMM_103_AWPROT = dm_AWPROT[103];
            assign M_AXIMM_103_AWREGION = dm_AWREGION[103];
            assign M_AXIMM_103_AWQOS = dm_AWQOS[103];
            assign M_AXIMM_103_AWVALID = dm_AWVALID[103];
            assign dm_AWREADY[103] = M_AXIMM_103_AWREADY;
            assign M_AXIMM_103_WDATA = dm_WDATA[103][M_AXIMM_103_DATA_WIDTH-1:0];
            assign M_AXIMM_103_WSTRB = dm_WSTRB[103][M_AXIMM_103_DATA_WIDTH/8-1:0];
            assign M_AXIMM_103_WLAST = dm_WLAST[103];
            assign M_AXIMM_103_WVALID = dm_WVALID[103];
            assign dm_WREADY[103] = M_AXIMM_103_WREADY;
            assign dm_BRESP[103] = M_AXIMM_103_BRESP;
            assign dm_BVALID[103] = M_AXIMM_103_BVALID;
            assign M_AXIMM_103_BREADY = dm_BREADY[103];
            assign M_AXIMM_103_ARADDR = dm_ARADDR[103][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_103_ARLEN = dm_ARLEN[103];
            assign M_AXIMM_103_ARSIZE = dm_ARSIZE[103];
            assign M_AXIMM_103_ARBURST = dm_ARBURST[103];
            assign M_AXIMM_103_ARLOCK = dm_ARLOCK[103];
            assign M_AXIMM_103_ARCACHE = dm_ARCACHE[103];
            assign M_AXIMM_103_ARPROT = dm_ARPROT[103];
            assign M_AXIMM_103_ARREGION = dm_ARREGION[103];
            assign M_AXIMM_103_ARQOS = dm_ARQOS[103];
            assign M_AXIMM_103_ARVALID = dm_ARVALID[103];
            assign dm_ARREADY[103] = M_AXIMM_103_ARREADY;
            assign dm_RDATA[103][M_AXIMM_103_DATA_WIDTH-1:0] = M_AXIMM_103_RDATA;
            assign dm_RRESP[103] = M_AXIMM_103_RRESP;
            assign dm_RLAST[103] = M_AXIMM_103_RLAST;
            assign dm_RVALID[103] = M_AXIMM_103_RVALID;
            assign M_AXIMM_103_RREADY = dm_RREADY[103];
        end
        if(C_NUM_AXIMMs > 104) begin
            assign ap_AWADDR[104][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_104_AWADDR;
            assign ap_AWLEN[104] = AP_AXIMM_104_AWLEN;
            assign ap_AWSIZE[104] = AP_AXIMM_104_AWSIZE;
            assign ap_AWBURST[104] = AP_AXIMM_104_AWBURST;
            assign ap_AWLOCK[104] = AP_AXIMM_104_AWLOCK;
            assign ap_AWCACHE[104] = AP_AXIMM_104_AWCACHE;
            assign ap_AWPROT[104] = AP_AXIMM_104_AWPROT;
            assign ap_AWREGION[104] = AP_AXIMM_104_AWREGION;
            assign ap_AWQOS[104] = AP_AXIMM_104_AWQOS;
            assign ap_AWVALID[104] = AP_AXIMM_104_AWVALID;
            assign AP_AXIMM_104_AWREADY = ap_AWREADY[104];
            assign ap_WDATA[104][M_AXIMM_104_DATA_WIDTH-1:0] = AP_AXIMM_104_WDATA;
            assign ap_WSTRB[104][M_AXIMM_104_DATA_WIDTH/8-1:0] = AP_AXIMM_104_WSTRB;
            assign ap_WLAST[104] = AP_AXIMM_104_WLAST;
            assign ap_WVALID[104] = AP_AXIMM_104_WVALID;
            assign AP_AXIMM_104_WREADY = ap_WREADY[104];
            assign AP_AXIMM_104_BRESP = ap_BRESP[104];
            assign AP_AXIMM_104_BVALID = ap_BVALID[104];
            assign ap_BREADY[104] = AP_AXIMM_104_BREADY;
            assign ap_ARADDR[104][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_104_ARADDR;
            assign ap_ARLEN[104] = AP_AXIMM_104_ARLEN;
            assign ap_ARSIZE[104] = AP_AXIMM_104_ARSIZE;
            assign ap_ARBURST[104] = AP_AXIMM_104_ARBURST;
            assign ap_ARLOCK[104] = AP_AXIMM_104_ARLOCK;
            assign ap_ARCACHE[104] = AP_AXIMM_104_ARCACHE;
            assign ap_ARPROT[104] = AP_AXIMM_104_ARPROT;
            assign ap_ARREGION[104] = AP_AXIMM_104_ARREGION;
            assign ap_ARQOS[104] = AP_AXIMM_104_ARQOS;
            assign ap_ARVALID[104] = AP_AXIMM_104_ARVALID;
            assign AP_AXIMM_104_ARREADY = ap_ARREADY[104];
            assign AP_AXIMM_104_RDATA = ap_RDATA[104][M_AXIMM_104_DATA_WIDTH-1:0];
            assign AP_AXIMM_104_RRESP = ap_RRESP[104];
            assign AP_AXIMM_104_RLAST = ap_RLAST[104];
            assign AP_AXIMM_104_RVALID = ap_RVALID[104];
            assign ap_RREADY[104] = AP_AXIMM_104_RREADY;
            assign M_AXIMM_104_AWADDR = dm_AWADDR[104][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_104_AWLEN = dm_AWLEN[104];
            assign M_AXIMM_104_AWSIZE = dm_AWSIZE[104];
            assign M_AXIMM_104_AWBURST = dm_AWBURST[104];
            assign M_AXIMM_104_AWLOCK = dm_AWLOCK[104];
            assign M_AXIMM_104_AWCACHE = dm_AWCACHE[104];
            assign M_AXIMM_104_AWPROT = dm_AWPROT[104];
            assign M_AXIMM_104_AWREGION = dm_AWREGION[104];
            assign M_AXIMM_104_AWQOS = dm_AWQOS[104];
            assign M_AXIMM_104_AWVALID = dm_AWVALID[104];
            assign dm_AWREADY[104] = M_AXIMM_104_AWREADY;
            assign M_AXIMM_104_WDATA = dm_WDATA[104][M_AXIMM_104_DATA_WIDTH-1:0];
            assign M_AXIMM_104_WSTRB = dm_WSTRB[104][M_AXIMM_104_DATA_WIDTH/8-1:0];
            assign M_AXIMM_104_WLAST = dm_WLAST[104];
            assign M_AXIMM_104_WVALID = dm_WVALID[104];
            assign dm_WREADY[104] = M_AXIMM_104_WREADY;
            assign dm_BRESP[104] = M_AXIMM_104_BRESP;
            assign dm_BVALID[104] = M_AXIMM_104_BVALID;
            assign M_AXIMM_104_BREADY = dm_BREADY[104];
            assign M_AXIMM_104_ARADDR = dm_ARADDR[104][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_104_ARLEN = dm_ARLEN[104];
            assign M_AXIMM_104_ARSIZE = dm_ARSIZE[104];
            assign M_AXIMM_104_ARBURST = dm_ARBURST[104];
            assign M_AXIMM_104_ARLOCK = dm_ARLOCK[104];
            assign M_AXIMM_104_ARCACHE = dm_ARCACHE[104];
            assign M_AXIMM_104_ARPROT = dm_ARPROT[104];
            assign M_AXIMM_104_ARREGION = dm_ARREGION[104];
            assign M_AXIMM_104_ARQOS = dm_ARQOS[104];
            assign M_AXIMM_104_ARVALID = dm_ARVALID[104];
            assign dm_ARREADY[104] = M_AXIMM_104_ARREADY;
            assign dm_RDATA[104][M_AXIMM_104_DATA_WIDTH-1:0] = M_AXIMM_104_RDATA;
            assign dm_RRESP[104] = M_AXIMM_104_RRESP;
            assign dm_RLAST[104] = M_AXIMM_104_RLAST;
            assign dm_RVALID[104] = M_AXIMM_104_RVALID;
            assign M_AXIMM_104_RREADY = dm_RREADY[104];
        end
        if(C_NUM_AXIMMs > 105) begin
            assign ap_AWADDR[105][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_105_AWADDR;
            assign ap_AWLEN[105] = AP_AXIMM_105_AWLEN;
            assign ap_AWSIZE[105] = AP_AXIMM_105_AWSIZE;
            assign ap_AWBURST[105] = AP_AXIMM_105_AWBURST;
            assign ap_AWLOCK[105] = AP_AXIMM_105_AWLOCK;
            assign ap_AWCACHE[105] = AP_AXIMM_105_AWCACHE;
            assign ap_AWPROT[105] = AP_AXIMM_105_AWPROT;
            assign ap_AWREGION[105] = AP_AXIMM_105_AWREGION;
            assign ap_AWQOS[105] = AP_AXIMM_105_AWQOS;
            assign ap_AWVALID[105] = AP_AXIMM_105_AWVALID;
            assign AP_AXIMM_105_AWREADY = ap_AWREADY[105];
            assign ap_WDATA[105][M_AXIMM_105_DATA_WIDTH-1:0] = AP_AXIMM_105_WDATA;
            assign ap_WSTRB[105][M_AXIMM_105_DATA_WIDTH/8-1:0] = AP_AXIMM_105_WSTRB;
            assign ap_WLAST[105] = AP_AXIMM_105_WLAST;
            assign ap_WVALID[105] = AP_AXIMM_105_WVALID;
            assign AP_AXIMM_105_WREADY = ap_WREADY[105];
            assign AP_AXIMM_105_BRESP = ap_BRESP[105];
            assign AP_AXIMM_105_BVALID = ap_BVALID[105];
            assign ap_BREADY[105] = AP_AXIMM_105_BREADY;
            assign ap_ARADDR[105][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_105_ARADDR;
            assign ap_ARLEN[105] = AP_AXIMM_105_ARLEN;
            assign ap_ARSIZE[105] = AP_AXIMM_105_ARSIZE;
            assign ap_ARBURST[105] = AP_AXIMM_105_ARBURST;
            assign ap_ARLOCK[105] = AP_AXIMM_105_ARLOCK;
            assign ap_ARCACHE[105] = AP_AXIMM_105_ARCACHE;
            assign ap_ARPROT[105] = AP_AXIMM_105_ARPROT;
            assign ap_ARREGION[105] = AP_AXIMM_105_ARREGION;
            assign ap_ARQOS[105] = AP_AXIMM_105_ARQOS;
            assign ap_ARVALID[105] = AP_AXIMM_105_ARVALID;
            assign AP_AXIMM_105_ARREADY = ap_ARREADY[105];
            assign AP_AXIMM_105_RDATA = ap_RDATA[105][M_AXIMM_105_DATA_WIDTH-1:0];
            assign AP_AXIMM_105_RRESP = ap_RRESP[105];
            assign AP_AXIMM_105_RLAST = ap_RLAST[105];
            assign AP_AXIMM_105_RVALID = ap_RVALID[105];
            assign ap_RREADY[105] = AP_AXIMM_105_RREADY;
            assign M_AXIMM_105_AWADDR = dm_AWADDR[105][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_105_AWLEN = dm_AWLEN[105];
            assign M_AXIMM_105_AWSIZE = dm_AWSIZE[105];
            assign M_AXIMM_105_AWBURST = dm_AWBURST[105];
            assign M_AXIMM_105_AWLOCK = dm_AWLOCK[105];
            assign M_AXIMM_105_AWCACHE = dm_AWCACHE[105];
            assign M_AXIMM_105_AWPROT = dm_AWPROT[105];
            assign M_AXIMM_105_AWREGION = dm_AWREGION[105];
            assign M_AXIMM_105_AWQOS = dm_AWQOS[105];
            assign M_AXIMM_105_AWVALID = dm_AWVALID[105];
            assign dm_AWREADY[105] = M_AXIMM_105_AWREADY;
            assign M_AXIMM_105_WDATA = dm_WDATA[105][M_AXIMM_105_DATA_WIDTH-1:0];
            assign M_AXIMM_105_WSTRB = dm_WSTRB[105][M_AXIMM_105_DATA_WIDTH/8-1:0];
            assign M_AXIMM_105_WLAST = dm_WLAST[105];
            assign M_AXIMM_105_WVALID = dm_WVALID[105];
            assign dm_WREADY[105] = M_AXIMM_105_WREADY;
            assign dm_BRESP[105] = M_AXIMM_105_BRESP;
            assign dm_BVALID[105] = M_AXIMM_105_BVALID;
            assign M_AXIMM_105_BREADY = dm_BREADY[105];
            assign M_AXIMM_105_ARADDR = dm_ARADDR[105][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_105_ARLEN = dm_ARLEN[105];
            assign M_AXIMM_105_ARSIZE = dm_ARSIZE[105];
            assign M_AXIMM_105_ARBURST = dm_ARBURST[105];
            assign M_AXIMM_105_ARLOCK = dm_ARLOCK[105];
            assign M_AXIMM_105_ARCACHE = dm_ARCACHE[105];
            assign M_AXIMM_105_ARPROT = dm_ARPROT[105];
            assign M_AXIMM_105_ARREGION = dm_ARREGION[105];
            assign M_AXIMM_105_ARQOS = dm_ARQOS[105];
            assign M_AXIMM_105_ARVALID = dm_ARVALID[105];
            assign dm_ARREADY[105] = M_AXIMM_105_ARREADY;
            assign dm_RDATA[105][M_AXIMM_105_DATA_WIDTH-1:0] = M_AXIMM_105_RDATA;
            assign dm_RRESP[105] = M_AXIMM_105_RRESP;
            assign dm_RLAST[105] = M_AXIMM_105_RLAST;
            assign dm_RVALID[105] = M_AXIMM_105_RVALID;
            assign M_AXIMM_105_RREADY = dm_RREADY[105];
        end
        if(C_NUM_AXIMMs > 106) begin
            assign ap_AWADDR[106][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_106_AWADDR;
            assign ap_AWLEN[106] = AP_AXIMM_106_AWLEN;
            assign ap_AWSIZE[106] = AP_AXIMM_106_AWSIZE;
            assign ap_AWBURST[106] = AP_AXIMM_106_AWBURST;
            assign ap_AWLOCK[106] = AP_AXIMM_106_AWLOCK;
            assign ap_AWCACHE[106] = AP_AXIMM_106_AWCACHE;
            assign ap_AWPROT[106] = AP_AXIMM_106_AWPROT;
            assign ap_AWREGION[106] = AP_AXIMM_106_AWREGION;
            assign ap_AWQOS[106] = AP_AXIMM_106_AWQOS;
            assign ap_AWVALID[106] = AP_AXIMM_106_AWVALID;
            assign AP_AXIMM_106_AWREADY = ap_AWREADY[106];
            assign ap_WDATA[106][M_AXIMM_106_DATA_WIDTH-1:0] = AP_AXIMM_106_WDATA;
            assign ap_WSTRB[106][M_AXIMM_106_DATA_WIDTH/8-1:0] = AP_AXIMM_106_WSTRB;
            assign ap_WLAST[106] = AP_AXIMM_106_WLAST;
            assign ap_WVALID[106] = AP_AXIMM_106_WVALID;
            assign AP_AXIMM_106_WREADY = ap_WREADY[106];
            assign AP_AXIMM_106_BRESP = ap_BRESP[106];
            assign AP_AXIMM_106_BVALID = ap_BVALID[106];
            assign ap_BREADY[106] = AP_AXIMM_106_BREADY;
            assign ap_ARADDR[106][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_106_ARADDR;
            assign ap_ARLEN[106] = AP_AXIMM_106_ARLEN;
            assign ap_ARSIZE[106] = AP_AXIMM_106_ARSIZE;
            assign ap_ARBURST[106] = AP_AXIMM_106_ARBURST;
            assign ap_ARLOCK[106] = AP_AXIMM_106_ARLOCK;
            assign ap_ARCACHE[106] = AP_AXIMM_106_ARCACHE;
            assign ap_ARPROT[106] = AP_AXIMM_106_ARPROT;
            assign ap_ARREGION[106] = AP_AXIMM_106_ARREGION;
            assign ap_ARQOS[106] = AP_AXIMM_106_ARQOS;
            assign ap_ARVALID[106] = AP_AXIMM_106_ARVALID;
            assign AP_AXIMM_106_ARREADY = ap_ARREADY[106];
            assign AP_AXIMM_106_RDATA = ap_RDATA[106][M_AXIMM_106_DATA_WIDTH-1:0];
            assign AP_AXIMM_106_RRESP = ap_RRESP[106];
            assign AP_AXIMM_106_RLAST = ap_RLAST[106];
            assign AP_AXIMM_106_RVALID = ap_RVALID[106];
            assign ap_RREADY[106] = AP_AXIMM_106_RREADY;
            assign M_AXIMM_106_AWADDR = dm_AWADDR[106][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_106_AWLEN = dm_AWLEN[106];
            assign M_AXIMM_106_AWSIZE = dm_AWSIZE[106];
            assign M_AXIMM_106_AWBURST = dm_AWBURST[106];
            assign M_AXIMM_106_AWLOCK = dm_AWLOCK[106];
            assign M_AXIMM_106_AWCACHE = dm_AWCACHE[106];
            assign M_AXIMM_106_AWPROT = dm_AWPROT[106];
            assign M_AXIMM_106_AWREGION = dm_AWREGION[106];
            assign M_AXIMM_106_AWQOS = dm_AWQOS[106];
            assign M_AXIMM_106_AWVALID = dm_AWVALID[106];
            assign dm_AWREADY[106] = M_AXIMM_106_AWREADY;
            assign M_AXIMM_106_WDATA = dm_WDATA[106][M_AXIMM_106_DATA_WIDTH-1:0];
            assign M_AXIMM_106_WSTRB = dm_WSTRB[106][M_AXIMM_106_DATA_WIDTH/8-1:0];
            assign M_AXIMM_106_WLAST = dm_WLAST[106];
            assign M_AXIMM_106_WVALID = dm_WVALID[106];
            assign dm_WREADY[106] = M_AXIMM_106_WREADY;
            assign dm_BRESP[106] = M_AXIMM_106_BRESP;
            assign dm_BVALID[106] = M_AXIMM_106_BVALID;
            assign M_AXIMM_106_BREADY = dm_BREADY[106];
            assign M_AXIMM_106_ARADDR = dm_ARADDR[106][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_106_ARLEN = dm_ARLEN[106];
            assign M_AXIMM_106_ARSIZE = dm_ARSIZE[106];
            assign M_AXIMM_106_ARBURST = dm_ARBURST[106];
            assign M_AXIMM_106_ARLOCK = dm_ARLOCK[106];
            assign M_AXIMM_106_ARCACHE = dm_ARCACHE[106];
            assign M_AXIMM_106_ARPROT = dm_ARPROT[106];
            assign M_AXIMM_106_ARREGION = dm_ARREGION[106];
            assign M_AXIMM_106_ARQOS = dm_ARQOS[106];
            assign M_AXIMM_106_ARVALID = dm_ARVALID[106];
            assign dm_ARREADY[106] = M_AXIMM_106_ARREADY;
            assign dm_RDATA[106][M_AXIMM_106_DATA_WIDTH-1:0] = M_AXIMM_106_RDATA;
            assign dm_RRESP[106] = M_AXIMM_106_RRESP;
            assign dm_RLAST[106] = M_AXIMM_106_RLAST;
            assign dm_RVALID[106] = M_AXIMM_106_RVALID;
            assign M_AXIMM_106_RREADY = dm_RREADY[106];
        end
        if(C_NUM_AXIMMs > 107) begin
            assign ap_AWADDR[107][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_107_AWADDR;
            assign ap_AWLEN[107] = AP_AXIMM_107_AWLEN;
            assign ap_AWSIZE[107] = AP_AXIMM_107_AWSIZE;
            assign ap_AWBURST[107] = AP_AXIMM_107_AWBURST;
            assign ap_AWLOCK[107] = AP_AXIMM_107_AWLOCK;
            assign ap_AWCACHE[107] = AP_AXIMM_107_AWCACHE;
            assign ap_AWPROT[107] = AP_AXIMM_107_AWPROT;
            assign ap_AWREGION[107] = AP_AXIMM_107_AWREGION;
            assign ap_AWQOS[107] = AP_AXIMM_107_AWQOS;
            assign ap_AWVALID[107] = AP_AXIMM_107_AWVALID;
            assign AP_AXIMM_107_AWREADY = ap_AWREADY[107];
            assign ap_WDATA[107][M_AXIMM_107_DATA_WIDTH-1:0] = AP_AXIMM_107_WDATA;
            assign ap_WSTRB[107][M_AXIMM_107_DATA_WIDTH/8-1:0] = AP_AXIMM_107_WSTRB;
            assign ap_WLAST[107] = AP_AXIMM_107_WLAST;
            assign ap_WVALID[107] = AP_AXIMM_107_WVALID;
            assign AP_AXIMM_107_WREADY = ap_WREADY[107];
            assign AP_AXIMM_107_BRESP = ap_BRESP[107];
            assign AP_AXIMM_107_BVALID = ap_BVALID[107];
            assign ap_BREADY[107] = AP_AXIMM_107_BREADY;
            assign ap_ARADDR[107][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_107_ARADDR;
            assign ap_ARLEN[107] = AP_AXIMM_107_ARLEN;
            assign ap_ARSIZE[107] = AP_AXIMM_107_ARSIZE;
            assign ap_ARBURST[107] = AP_AXIMM_107_ARBURST;
            assign ap_ARLOCK[107] = AP_AXIMM_107_ARLOCK;
            assign ap_ARCACHE[107] = AP_AXIMM_107_ARCACHE;
            assign ap_ARPROT[107] = AP_AXIMM_107_ARPROT;
            assign ap_ARREGION[107] = AP_AXIMM_107_ARREGION;
            assign ap_ARQOS[107] = AP_AXIMM_107_ARQOS;
            assign ap_ARVALID[107] = AP_AXIMM_107_ARVALID;
            assign AP_AXIMM_107_ARREADY = ap_ARREADY[107];
            assign AP_AXIMM_107_RDATA = ap_RDATA[107][M_AXIMM_107_DATA_WIDTH-1:0];
            assign AP_AXIMM_107_RRESP = ap_RRESP[107];
            assign AP_AXIMM_107_RLAST = ap_RLAST[107];
            assign AP_AXIMM_107_RVALID = ap_RVALID[107];
            assign ap_RREADY[107] = AP_AXIMM_107_RREADY;
            assign M_AXIMM_107_AWADDR = dm_AWADDR[107][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_107_AWLEN = dm_AWLEN[107];
            assign M_AXIMM_107_AWSIZE = dm_AWSIZE[107];
            assign M_AXIMM_107_AWBURST = dm_AWBURST[107];
            assign M_AXIMM_107_AWLOCK = dm_AWLOCK[107];
            assign M_AXIMM_107_AWCACHE = dm_AWCACHE[107];
            assign M_AXIMM_107_AWPROT = dm_AWPROT[107];
            assign M_AXIMM_107_AWREGION = dm_AWREGION[107];
            assign M_AXIMM_107_AWQOS = dm_AWQOS[107];
            assign M_AXIMM_107_AWVALID = dm_AWVALID[107];
            assign dm_AWREADY[107] = M_AXIMM_107_AWREADY;
            assign M_AXIMM_107_WDATA = dm_WDATA[107][M_AXIMM_107_DATA_WIDTH-1:0];
            assign M_AXIMM_107_WSTRB = dm_WSTRB[107][M_AXIMM_107_DATA_WIDTH/8-1:0];
            assign M_AXIMM_107_WLAST = dm_WLAST[107];
            assign M_AXIMM_107_WVALID = dm_WVALID[107];
            assign dm_WREADY[107] = M_AXIMM_107_WREADY;
            assign dm_BRESP[107] = M_AXIMM_107_BRESP;
            assign dm_BVALID[107] = M_AXIMM_107_BVALID;
            assign M_AXIMM_107_BREADY = dm_BREADY[107];
            assign M_AXIMM_107_ARADDR = dm_ARADDR[107][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_107_ARLEN = dm_ARLEN[107];
            assign M_AXIMM_107_ARSIZE = dm_ARSIZE[107];
            assign M_AXIMM_107_ARBURST = dm_ARBURST[107];
            assign M_AXIMM_107_ARLOCK = dm_ARLOCK[107];
            assign M_AXIMM_107_ARCACHE = dm_ARCACHE[107];
            assign M_AXIMM_107_ARPROT = dm_ARPROT[107];
            assign M_AXIMM_107_ARREGION = dm_ARREGION[107];
            assign M_AXIMM_107_ARQOS = dm_ARQOS[107];
            assign M_AXIMM_107_ARVALID = dm_ARVALID[107];
            assign dm_ARREADY[107] = M_AXIMM_107_ARREADY;
            assign dm_RDATA[107][M_AXIMM_107_DATA_WIDTH-1:0] = M_AXIMM_107_RDATA;
            assign dm_RRESP[107] = M_AXIMM_107_RRESP;
            assign dm_RLAST[107] = M_AXIMM_107_RLAST;
            assign dm_RVALID[107] = M_AXIMM_107_RVALID;
            assign M_AXIMM_107_RREADY = dm_RREADY[107];
        end
        if(C_NUM_AXIMMs > 108) begin
            assign ap_AWADDR[108][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_108_AWADDR;
            assign ap_AWLEN[108] = AP_AXIMM_108_AWLEN;
            assign ap_AWSIZE[108] = AP_AXIMM_108_AWSIZE;
            assign ap_AWBURST[108] = AP_AXIMM_108_AWBURST;
            assign ap_AWLOCK[108] = AP_AXIMM_108_AWLOCK;
            assign ap_AWCACHE[108] = AP_AXIMM_108_AWCACHE;
            assign ap_AWPROT[108] = AP_AXIMM_108_AWPROT;
            assign ap_AWREGION[108] = AP_AXIMM_108_AWREGION;
            assign ap_AWQOS[108] = AP_AXIMM_108_AWQOS;
            assign ap_AWVALID[108] = AP_AXIMM_108_AWVALID;
            assign AP_AXIMM_108_AWREADY = ap_AWREADY[108];
            assign ap_WDATA[108][M_AXIMM_108_DATA_WIDTH-1:0] = AP_AXIMM_108_WDATA;
            assign ap_WSTRB[108][M_AXIMM_108_DATA_WIDTH/8-1:0] = AP_AXIMM_108_WSTRB;
            assign ap_WLAST[108] = AP_AXIMM_108_WLAST;
            assign ap_WVALID[108] = AP_AXIMM_108_WVALID;
            assign AP_AXIMM_108_WREADY = ap_WREADY[108];
            assign AP_AXIMM_108_BRESP = ap_BRESP[108];
            assign AP_AXIMM_108_BVALID = ap_BVALID[108];
            assign ap_BREADY[108] = AP_AXIMM_108_BREADY;
            assign ap_ARADDR[108][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_108_ARADDR;
            assign ap_ARLEN[108] = AP_AXIMM_108_ARLEN;
            assign ap_ARSIZE[108] = AP_AXIMM_108_ARSIZE;
            assign ap_ARBURST[108] = AP_AXIMM_108_ARBURST;
            assign ap_ARLOCK[108] = AP_AXIMM_108_ARLOCK;
            assign ap_ARCACHE[108] = AP_AXIMM_108_ARCACHE;
            assign ap_ARPROT[108] = AP_AXIMM_108_ARPROT;
            assign ap_ARREGION[108] = AP_AXIMM_108_ARREGION;
            assign ap_ARQOS[108] = AP_AXIMM_108_ARQOS;
            assign ap_ARVALID[108] = AP_AXIMM_108_ARVALID;
            assign AP_AXIMM_108_ARREADY = ap_ARREADY[108];
            assign AP_AXIMM_108_RDATA = ap_RDATA[108][M_AXIMM_108_DATA_WIDTH-1:0];
            assign AP_AXIMM_108_RRESP = ap_RRESP[108];
            assign AP_AXIMM_108_RLAST = ap_RLAST[108];
            assign AP_AXIMM_108_RVALID = ap_RVALID[108];
            assign ap_RREADY[108] = AP_AXIMM_108_RREADY;
            assign M_AXIMM_108_AWADDR = dm_AWADDR[108][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_108_AWLEN = dm_AWLEN[108];
            assign M_AXIMM_108_AWSIZE = dm_AWSIZE[108];
            assign M_AXIMM_108_AWBURST = dm_AWBURST[108];
            assign M_AXIMM_108_AWLOCK = dm_AWLOCK[108];
            assign M_AXIMM_108_AWCACHE = dm_AWCACHE[108];
            assign M_AXIMM_108_AWPROT = dm_AWPROT[108];
            assign M_AXIMM_108_AWREGION = dm_AWREGION[108];
            assign M_AXIMM_108_AWQOS = dm_AWQOS[108];
            assign M_AXIMM_108_AWVALID = dm_AWVALID[108];
            assign dm_AWREADY[108] = M_AXIMM_108_AWREADY;
            assign M_AXIMM_108_WDATA = dm_WDATA[108][M_AXIMM_108_DATA_WIDTH-1:0];
            assign M_AXIMM_108_WSTRB = dm_WSTRB[108][M_AXIMM_108_DATA_WIDTH/8-1:0];
            assign M_AXIMM_108_WLAST = dm_WLAST[108];
            assign M_AXIMM_108_WVALID = dm_WVALID[108];
            assign dm_WREADY[108] = M_AXIMM_108_WREADY;
            assign dm_BRESP[108] = M_AXIMM_108_BRESP;
            assign dm_BVALID[108] = M_AXIMM_108_BVALID;
            assign M_AXIMM_108_BREADY = dm_BREADY[108];
            assign M_AXIMM_108_ARADDR = dm_ARADDR[108][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_108_ARLEN = dm_ARLEN[108];
            assign M_AXIMM_108_ARSIZE = dm_ARSIZE[108];
            assign M_AXIMM_108_ARBURST = dm_ARBURST[108];
            assign M_AXIMM_108_ARLOCK = dm_ARLOCK[108];
            assign M_AXIMM_108_ARCACHE = dm_ARCACHE[108];
            assign M_AXIMM_108_ARPROT = dm_ARPROT[108];
            assign M_AXIMM_108_ARREGION = dm_ARREGION[108];
            assign M_AXIMM_108_ARQOS = dm_ARQOS[108];
            assign M_AXIMM_108_ARVALID = dm_ARVALID[108];
            assign dm_ARREADY[108] = M_AXIMM_108_ARREADY;
            assign dm_RDATA[108][M_AXIMM_108_DATA_WIDTH-1:0] = M_AXIMM_108_RDATA;
            assign dm_RRESP[108] = M_AXIMM_108_RRESP;
            assign dm_RLAST[108] = M_AXIMM_108_RLAST;
            assign dm_RVALID[108] = M_AXIMM_108_RVALID;
            assign M_AXIMM_108_RREADY = dm_RREADY[108];
        end
        if(C_NUM_AXIMMs > 109) begin
            assign ap_AWADDR[109][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_109_AWADDR;
            assign ap_AWLEN[109] = AP_AXIMM_109_AWLEN;
            assign ap_AWSIZE[109] = AP_AXIMM_109_AWSIZE;
            assign ap_AWBURST[109] = AP_AXIMM_109_AWBURST;
            assign ap_AWLOCK[109] = AP_AXIMM_109_AWLOCK;
            assign ap_AWCACHE[109] = AP_AXIMM_109_AWCACHE;
            assign ap_AWPROT[109] = AP_AXIMM_109_AWPROT;
            assign ap_AWREGION[109] = AP_AXIMM_109_AWREGION;
            assign ap_AWQOS[109] = AP_AXIMM_109_AWQOS;
            assign ap_AWVALID[109] = AP_AXIMM_109_AWVALID;
            assign AP_AXIMM_109_AWREADY = ap_AWREADY[109];
            assign ap_WDATA[109][M_AXIMM_109_DATA_WIDTH-1:0] = AP_AXIMM_109_WDATA;
            assign ap_WSTRB[109][M_AXIMM_109_DATA_WIDTH/8-1:0] = AP_AXIMM_109_WSTRB;
            assign ap_WLAST[109] = AP_AXIMM_109_WLAST;
            assign ap_WVALID[109] = AP_AXIMM_109_WVALID;
            assign AP_AXIMM_109_WREADY = ap_WREADY[109];
            assign AP_AXIMM_109_BRESP = ap_BRESP[109];
            assign AP_AXIMM_109_BVALID = ap_BVALID[109];
            assign ap_BREADY[109] = AP_AXIMM_109_BREADY;
            assign ap_ARADDR[109][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_109_ARADDR;
            assign ap_ARLEN[109] = AP_AXIMM_109_ARLEN;
            assign ap_ARSIZE[109] = AP_AXIMM_109_ARSIZE;
            assign ap_ARBURST[109] = AP_AXIMM_109_ARBURST;
            assign ap_ARLOCK[109] = AP_AXIMM_109_ARLOCK;
            assign ap_ARCACHE[109] = AP_AXIMM_109_ARCACHE;
            assign ap_ARPROT[109] = AP_AXIMM_109_ARPROT;
            assign ap_ARREGION[109] = AP_AXIMM_109_ARREGION;
            assign ap_ARQOS[109] = AP_AXIMM_109_ARQOS;
            assign ap_ARVALID[109] = AP_AXIMM_109_ARVALID;
            assign AP_AXIMM_109_ARREADY = ap_ARREADY[109];
            assign AP_AXIMM_109_RDATA = ap_RDATA[109][M_AXIMM_109_DATA_WIDTH-1:0];
            assign AP_AXIMM_109_RRESP = ap_RRESP[109];
            assign AP_AXIMM_109_RLAST = ap_RLAST[109];
            assign AP_AXIMM_109_RVALID = ap_RVALID[109];
            assign ap_RREADY[109] = AP_AXIMM_109_RREADY;
            assign M_AXIMM_109_AWADDR = dm_AWADDR[109][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_109_AWLEN = dm_AWLEN[109];
            assign M_AXIMM_109_AWSIZE = dm_AWSIZE[109];
            assign M_AXIMM_109_AWBURST = dm_AWBURST[109];
            assign M_AXIMM_109_AWLOCK = dm_AWLOCK[109];
            assign M_AXIMM_109_AWCACHE = dm_AWCACHE[109];
            assign M_AXIMM_109_AWPROT = dm_AWPROT[109];
            assign M_AXIMM_109_AWREGION = dm_AWREGION[109];
            assign M_AXIMM_109_AWQOS = dm_AWQOS[109];
            assign M_AXIMM_109_AWVALID = dm_AWVALID[109];
            assign dm_AWREADY[109] = M_AXIMM_109_AWREADY;
            assign M_AXIMM_109_WDATA = dm_WDATA[109][M_AXIMM_109_DATA_WIDTH-1:0];
            assign M_AXIMM_109_WSTRB = dm_WSTRB[109][M_AXIMM_109_DATA_WIDTH/8-1:0];
            assign M_AXIMM_109_WLAST = dm_WLAST[109];
            assign M_AXIMM_109_WVALID = dm_WVALID[109];
            assign dm_WREADY[109] = M_AXIMM_109_WREADY;
            assign dm_BRESP[109] = M_AXIMM_109_BRESP;
            assign dm_BVALID[109] = M_AXIMM_109_BVALID;
            assign M_AXIMM_109_BREADY = dm_BREADY[109];
            assign M_AXIMM_109_ARADDR = dm_ARADDR[109][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_109_ARLEN = dm_ARLEN[109];
            assign M_AXIMM_109_ARSIZE = dm_ARSIZE[109];
            assign M_AXIMM_109_ARBURST = dm_ARBURST[109];
            assign M_AXIMM_109_ARLOCK = dm_ARLOCK[109];
            assign M_AXIMM_109_ARCACHE = dm_ARCACHE[109];
            assign M_AXIMM_109_ARPROT = dm_ARPROT[109];
            assign M_AXIMM_109_ARREGION = dm_ARREGION[109];
            assign M_AXIMM_109_ARQOS = dm_ARQOS[109];
            assign M_AXIMM_109_ARVALID = dm_ARVALID[109];
            assign dm_ARREADY[109] = M_AXIMM_109_ARREADY;
            assign dm_RDATA[109][M_AXIMM_109_DATA_WIDTH-1:0] = M_AXIMM_109_RDATA;
            assign dm_RRESP[109] = M_AXIMM_109_RRESP;
            assign dm_RLAST[109] = M_AXIMM_109_RLAST;
            assign dm_RVALID[109] = M_AXIMM_109_RVALID;
            assign M_AXIMM_109_RREADY = dm_RREADY[109];
        end
        if(C_NUM_AXIMMs > 110) begin
            assign ap_AWADDR[110][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_110_AWADDR;
            assign ap_AWLEN[110] = AP_AXIMM_110_AWLEN;
            assign ap_AWSIZE[110] = AP_AXIMM_110_AWSIZE;
            assign ap_AWBURST[110] = AP_AXIMM_110_AWBURST;
            assign ap_AWLOCK[110] = AP_AXIMM_110_AWLOCK;
            assign ap_AWCACHE[110] = AP_AXIMM_110_AWCACHE;
            assign ap_AWPROT[110] = AP_AXIMM_110_AWPROT;
            assign ap_AWREGION[110] = AP_AXIMM_110_AWREGION;
            assign ap_AWQOS[110] = AP_AXIMM_110_AWQOS;
            assign ap_AWVALID[110] = AP_AXIMM_110_AWVALID;
            assign AP_AXIMM_110_AWREADY = ap_AWREADY[110];
            assign ap_WDATA[110][M_AXIMM_110_DATA_WIDTH-1:0] = AP_AXIMM_110_WDATA;
            assign ap_WSTRB[110][M_AXIMM_110_DATA_WIDTH/8-1:0] = AP_AXIMM_110_WSTRB;
            assign ap_WLAST[110] = AP_AXIMM_110_WLAST;
            assign ap_WVALID[110] = AP_AXIMM_110_WVALID;
            assign AP_AXIMM_110_WREADY = ap_WREADY[110];
            assign AP_AXIMM_110_BRESP = ap_BRESP[110];
            assign AP_AXIMM_110_BVALID = ap_BVALID[110];
            assign ap_BREADY[110] = AP_AXIMM_110_BREADY;
            assign ap_ARADDR[110][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_110_ARADDR;
            assign ap_ARLEN[110] = AP_AXIMM_110_ARLEN;
            assign ap_ARSIZE[110] = AP_AXIMM_110_ARSIZE;
            assign ap_ARBURST[110] = AP_AXIMM_110_ARBURST;
            assign ap_ARLOCK[110] = AP_AXIMM_110_ARLOCK;
            assign ap_ARCACHE[110] = AP_AXIMM_110_ARCACHE;
            assign ap_ARPROT[110] = AP_AXIMM_110_ARPROT;
            assign ap_ARREGION[110] = AP_AXIMM_110_ARREGION;
            assign ap_ARQOS[110] = AP_AXIMM_110_ARQOS;
            assign ap_ARVALID[110] = AP_AXIMM_110_ARVALID;
            assign AP_AXIMM_110_ARREADY = ap_ARREADY[110];
            assign AP_AXIMM_110_RDATA = ap_RDATA[110][M_AXIMM_110_DATA_WIDTH-1:0];
            assign AP_AXIMM_110_RRESP = ap_RRESP[110];
            assign AP_AXIMM_110_RLAST = ap_RLAST[110];
            assign AP_AXIMM_110_RVALID = ap_RVALID[110];
            assign ap_RREADY[110] = AP_AXIMM_110_RREADY;
            assign M_AXIMM_110_AWADDR = dm_AWADDR[110][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_110_AWLEN = dm_AWLEN[110];
            assign M_AXIMM_110_AWSIZE = dm_AWSIZE[110];
            assign M_AXIMM_110_AWBURST = dm_AWBURST[110];
            assign M_AXIMM_110_AWLOCK = dm_AWLOCK[110];
            assign M_AXIMM_110_AWCACHE = dm_AWCACHE[110];
            assign M_AXIMM_110_AWPROT = dm_AWPROT[110];
            assign M_AXIMM_110_AWREGION = dm_AWREGION[110];
            assign M_AXIMM_110_AWQOS = dm_AWQOS[110];
            assign M_AXIMM_110_AWVALID = dm_AWVALID[110];
            assign dm_AWREADY[110] = M_AXIMM_110_AWREADY;
            assign M_AXIMM_110_WDATA = dm_WDATA[110][M_AXIMM_110_DATA_WIDTH-1:0];
            assign M_AXIMM_110_WSTRB = dm_WSTRB[110][M_AXIMM_110_DATA_WIDTH/8-1:0];
            assign M_AXIMM_110_WLAST = dm_WLAST[110];
            assign M_AXIMM_110_WVALID = dm_WVALID[110];
            assign dm_WREADY[110] = M_AXIMM_110_WREADY;
            assign dm_BRESP[110] = M_AXIMM_110_BRESP;
            assign dm_BVALID[110] = M_AXIMM_110_BVALID;
            assign M_AXIMM_110_BREADY = dm_BREADY[110];
            assign M_AXIMM_110_ARADDR = dm_ARADDR[110][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_110_ARLEN = dm_ARLEN[110];
            assign M_AXIMM_110_ARSIZE = dm_ARSIZE[110];
            assign M_AXIMM_110_ARBURST = dm_ARBURST[110];
            assign M_AXIMM_110_ARLOCK = dm_ARLOCK[110];
            assign M_AXIMM_110_ARCACHE = dm_ARCACHE[110];
            assign M_AXIMM_110_ARPROT = dm_ARPROT[110];
            assign M_AXIMM_110_ARREGION = dm_ARREGION[110];
            assign M_AXIMM_110_ARQOS = dm_ARQOS[110];
            assign M_AXIMM_110_ARVALID = dm_ARVALID[110];
            assign dm_ARREADY[110] = M_AXIMM_110_ARREADY;
            assign dm_RDATA[110][M_AXIMM_110_DATA_WIDTH-1:0] = M_AXIMM_110_RDATA;
            assign dm_RRESP[110] = M_AXIMM_110_RRESP;
            assign dm_RLAST[110] = M_AXIMM_110_RLAST;
            assign dm_RVALID[110] = M_AXIMM_110_RVALID;
            assign M_AXIMM_110_RREADY = dm_RREADY[110];
        end
        if(C_NUM_AXIMMs > 111) begin
            assign ap_AWADDR[111][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_111_AWADDR;
            assign ap_AWLEN[111] = AP_AXIMM_111_AWLEN;
            assign ap_AWSIZE[111] = AP_AXIMM_111_AWSIZE;
            assign ap_AWBURST[111] = AP_AXIMM_111_AWBURST;
            assign ap_AWLOCK[111] = AP_AXIMM_111_AWLOCK;
            assign ap_AWCACHE[111] = AP_AXIMM_111_AWCACHE;
            assign ap_AWPROT[111] = AP_AXIMM_111_AWPROT;
            assign ap_AWREGION[111] = AP_AXIMM_111_AWREGION;
            assign ap_AWQOS[111] = AP_AXIMM_111_AWQOS;
            assign ap_AWVALID[111] = AP_AXIMM_111_AWVALID;
            assign AP_AXIMM_111_AWREADY = ap_AWREADY[111];
            assign ap_WDATA[111][M_AXIMM_111_DATA_WIDTH-1:0] = AP_AXIMM_111_WDATA;
            assign ap_WSTRB[111][M_AXIMM_111_DATA_WIDTH/8-1:0] = AP_AXIMM_111_WSTRB;
            assign ap_WLAST[111] = AP_AXIMM_111_WLAST;
            assign ap_WVALID[111] = AP_AXIMM_111_WVALID;
            assign AP_AXIMM_111_WREADY = ap_WREADY[111];
            assign AP_AXIMM_111_BRESP = ap_BRESP[111];
            assign AP_AXIMM_111_BVALID = ap_BVALID[111];
            assign ap_BREADY[111] = AP_AXIMM_111_BREADY;
            assign ap_ARADDR[111][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_111_ARADDR;
            assign ap_ARLEN[111] = AP_AXIMM_111_ARLEN;
            assign ap_ARSIZE[111] = AP_AXIMM_111_ARSIZE;
            assign ap_ARBURST[111] = AP_AXIMM_111_ARBURST;
            assign ap_ARLOCK[111] = AP_AXIMM_111_ARLOCK;
            assign ap_ARCACHE[111] = AP_AXIMM_111_ARCACHE;
            assign ap_ARPROT[111] = AP_AXIMM_111_ARPROT;
            assign ap_ARREGION[111] = AP_AXIMM_111_ARREGION;
            assign ap_ARQOS[111] = AP_AXIMM_111_ARQOS;
            assign ap_ARVALID[111] = AP_AXIMM_111_ARVALID;
            assign AP_AXIMM_111_ARREADY = ap_ARREADY[111];
            assign AP_AXIMM_111_RDATA = ap_RDATA[111][M_AXIMM_111_DATA_WIDTH-1:0];
            assign AP_AXIMM_111_RRESP = ap_RRESP[111];
            assign AP_AXIMM_111_RLAST = ap_RLAST[111];
            assign AP_AXIMM_111_RVALID = ap_RVALID[111];
            assign ap_RREADY[111] = AP_AXIMM_111_RREADY;
            assign M_AXIMM_111_AWADDR = dm_AWADDR[111][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_111_AWLEN = dm_AWLEN[111];
            assign M_AXIMM_111_AWSIZE = dm_AWSIZE[111];
            assign M_AXIMM_111_AWBURST = dm_AWBURST[111];
            assign M_AXIMM_111_AWLOCK = dm_AWLOCK[111];
            assign M_AXIMM_111_AWCACHE = dm_AWCACHE[111];
            assign M_AXIMM_111_AWPROT = dm_AWPROT[111];
            assign M_AXIMM_111_AWREGION = dm_AWREGION[111];
            assign M_AXIMM_111_AWQOS = dm_AWQOS[111];
            assign M_AXIMM_111_AWVALID = dm_AWVALID[111];
            assign dm_AWREADY[111] = M_AXIMM_111_AWREADY;
            assign M_AXIMM_111_WDATA = dm_WDATA[111][M_AXIMM_111_DATA_WIDTH-1:0];
            assign M_AXIMM_111_WSTRB = dm_WSTRB[111][M_AXIMM_111_DATA_WIDTH/8-1:0];
            assign M_AXIMM_111_WLAST = dm_WLAST[111];
            assign M_AXIMM_111_WVALID = dm_WVALID[111];
            assign dm_WREADY[111] = M_AXIMM_111_WREADY;
            assign dm_BRESP[111] = M_AXIMM_111_BRESP;
            assign dm_BVALID[111] = M_AXIMM_111_BVALID;
            assign M_AXIMM_111_BREADY = dm_BREADY[111];
            assign M_AXIMM_111_ARADDR = dm_ARADDR[111][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_111_ARLEN = dm_ARLEN[111];
            assign M_AXIMM_111_ARSIZE = dm_ARSIZE[111];
            assign M_AXIMM_111_ARBURST = dm_ARBURST[111];
            assign M_AXIMM_111_ARLOCK = dm_ARLOCK[111];
            assign M_AXIMM_111_ARCACHE = dm_ARCACHE[111];
            assign M_AXIMM_111_ARPROT = dm_ARPROT[111];
            assign M_AXIMM_111_ARREGION = dm_ARREGION[111];
            assign M_AXIMM_111_ARQOS = dm_ARQOS[111];
            assign M_AXIMM_111_ARVALID = dm_ARVALID[111];
            assign dm_ARREADY[111] = M_AXIMM_111_ARREADY;
            assign dm_RDATA[111][M_AXIMM_111_DATA_WIDTH-1:0] = M_AXIMM_111_RDATA;
            assign dm_RRESP[111] = M_AXIMM_111_RRESP;
            assign dm_RLAST[111] = M_AXIMM_111_RLAST;
            assign dm_RVALID[111] = M_AXIMM_111_RVALID;
            assign M_AXIMM_111_RREADY = dm_RREADY[111];
        end
        if(C_NUM_AXIMMs > 112) begin
            assign ap_AWADDR[112][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_112_AWADDR;
            assign ap_AWLEN[112] = AP_AXIMM_112_AWLEN;
            assign ap_AWSIZE[112] = AP_AXIMM_112_AWSIZE;
            assign ap_AWBURST[112] = AP_AXIMM_112_AWBURST;
            assign ap_AWLOCK[112] = AP_AXIMM_112_AWLOCK;
            assign ap_AWCACHE[112] = AP_AXIMM_112_AWCACHE;
            assign ap_AWPROT[112] = AP_AXIMM_112_AWPROT;
            assign ap_AWREGION[112] = AP_AXIMM_112_AWREGION;
            assign ap_AWQOS[112] = AP_AXIMM_112_AWQOS;
            assign ap_AWVALID[112] = AP_AXIMM_112_AWVALID;
            assign AP_AXIMM_112_AWREADY = ap_AWREADY[112];
            assign ap_WDATA[112][M_AXIMM_112_DATA_WIDTH-1:0] = AP_AXIMM_112_WDATA;
            assign ap_WSTRB[112][M_AXIMM_112_DATA_WIDTH/8-1:0] = AP_AXIMM_112_WSTRB;
            assign ap_WLAST[112] = AP_AXIMM_112_WLAST;
            assign ap_WVALID[112] = AP_AXIMM_112_WVALID;
            assign AP_AXIMM_112_WREADY = ap_WREADY[112];
            assign AP_AXIMM_112_BRESP = ap_BRESP[112];
            assign AP_AXIMM_112_BVALID = ap_BVALID[112];
            assign ap_BREADY[112] = AP_AXIMM_112_BREADY;
            assign ap_ARADDR[112][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_112_ARADDR;
            assign ap_ARLEN[112] = AP_AXIMM_112_ARLEN;
            assign ap_ARSIZE[112] = AP_AXIMM_112_ARSIZE;
            assign ap_ARBURST[112] = AP_AXIMM_112_ARBURST;
            assign ap_ARLOCK[112] = AP_AXIMM_112_ARLOCK;
            assign ap_ARCACHE[112] = AP_AXIMM_112_ARCACHE;
            assign ap_ARPROT[112] = AP_AXIMM_112_ARPROT;
            assign ap_ARREGION[112] = AP_AXIMM_112_ARREGION;
            assign ap_ARQOS[112] = AP_AXIMM_112_ARQOS;
            assign ap_ARVALID[112] = AP_AXIMM_112_ARVALID;
            assign AP_AXIMM_112_ARREADY = ap_ARREADY[112];
            assign AP_AXIMM_112_RDATA = ap_RDATA[112][M_AXIMM_112_DATA_WIDTH-1:0];
            assign AP_AXIMM_112_RRESP = ap_RRESP[112];
            assign AP_AXIMM_112_RLAST = ap_RLAST[112];
            assign AP_AXIMM_112_RVALID = ap_RVALID[112];
            assign ap_RREADY[112] = AP_AXIMM_112_RREADY;
            assign M_AXIMM_112_AWADDR = dm_AWADDR[112][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_112_AWLEN = dm_AWLEN[112];
            assign M_AXIMM_112_AWSIZE = dm_AWSIZE[112];
            assign M_AXIMM_112_AWBURST = dm_AWBURST[112];
            assign M_AXIMM_112_AWLOCK = dm_AWLOCK[112];
            assign M_AXIMM_112_AWCACHE = dm_AWCACHE[112];
            assign M_AXIMM_112_AWPROT = dm_AWPROT[112];
            assign M_AXIMM_112_AWREGION = dm_AWREGION[112];
            assign M_AXIMM_112_AWQOS = dm_AWQOS[112];
            assign M_AXIMM_112_AWVALID = dm_AWVALID[112];
            assign dm_AWREADY[112] = M_AXIMM_112_AWREADY;
            assign M_AXIMM_112_WDATA = dm_WDATA[112][M_AXIMM_112_DATA_WIDTH-1:0];
            assign M_AXIMM_112_WSTRB = dm_WSTRB[112][M_AXIMM_112_DATA_WIDTH/8-1:0];
            assign M_AXIMM_112_WLAST = dm_WLAST[112];
            assign M_AXIMM_112_WVALID = dm_WVALID[112];
            assign dm_WREADY[112] = M_AXIMM_112_WREADY;
            assign dm_BRESP[112] = M_AXIMM_112_BRESP;
            assign dm_BVALID[112] = M_AXIMM_112_BVALID;
            assign M_AXIMM_112_BREADY = dm_BREADY[112];
            assign M_AXIMM_112_ARADDR = dm_ARADDR[112][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_112_ARLEN = dm_ARLEN[112];
            assign M_AXIMM_112_ARSIZE = dm_ARSIZE[112];
            assign M_AXIMM_112_ARBURST = dm_ARBURST[112];
            assign M_AXIMM_112_ARLOCK = dm_ARLOCK[112];
            assign M_AXIMM_112_ARCACHE = dm_ARCACHE[112];
            assign M_AXIMM_112_ARPROT = dm_ARPROT[112];
            assign M_AXIMM_112_ARREGION = dm_ARREGION[112];
            assign M_AXIMM_112_ARQOS = dm_ARQOS[112];
            assign M_AXIMM_112_ARVALID = dm_ARVALID[112];
            assign dm_ARREADY[112] = M_AXIMM_112_ARREADY;
            assign dm_RDATA[112][M_AXIMM_112_DATA_WIDTH-1:0] = M_AXIMM_112_RDATA;
            assign dm_RRESP[112] = M_AXIMM_112_RRESP;
            assign dm_RLAST[112] = M_AXIMM_112_RLAST;
            assign dm_RVALID[112] = M_AXIMM_112_RVALID;
            assign M_AXIMM_112_RREADY = dm_RREADY[112];
        end
        if(C_NUM_AXIMMs > 113) begin
            assign ap_AWADDR[113][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_113_AWADDR;
            assign ap_AWLEN[113] = AP_AXIMM_113_AWLEN;
            assign ap_AWSIZE[113] = AP_AXIMM_113_AWSIZE;
            assign ap_AWBURST[113] = AP_AXIMM_113_AWBURST;
            assign ap_AWLOCK[113] = AP_AXIMM_113_AWLOCK;
            assign ap_AWCACHE[113] = AP_AXIMM_113_AWCACHE;
            assign ap_AWPROT[113] = AP_AXIMM_113_AWPROT;
            assign ap_AWREGION[113] = AP_AXIMM_113_AWREGION;
            assign ap_AWQOS[113] = AP_AXIMM_113_AWQOS;
            assign ap_AWVALID[113] = AP_AXIMM_113_AWVALID;
            assign AP_AXIMM_113_AWREADY = ap_AWREADY[113];
            assign ap_WDATA[113][M_AXIMM_113_DATA_WIDTH-1:0] = AP_AXIMM_113_WDATA;
            assign ap_WSTRB[113][M_AXIMM_113_DATA_WIDTH/8-1:0] = AP_AXIMM_113_WSTRB;
            assign ap_WLAST[113] = AP_AXIMM_113_WLAST;
            assign ap_WVALID[113] = AP_AXIMM_113_WVALID;
            assign AP_AXIMM_113_WREADY = ap_WREADY[113];
            assign AP_AXIMM_113_BRESP = ap_BRESP[113];
            assign AP_AXIMM_113_BVALID = ap_BVALID[113];
            assign ap_BREADY[113] = AP_AXIMM_113_BREADY;
            assign ap_ARADDR[113][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_113_ARADDR;
            assign ap_ARLEN[113] = AP_AXIMM_113_ARLEN;
            assign ap_ARSIZE[113] = AP_AXIMM_113_ARSIZE;
            assign ap_ARBURST[113] = AP_AXIMM_113_ARBURST;
            assign ap_ARLOCK[113] = AP_AXIMM_113_ARLOCK;
            assign ap_ARCACHE[113] = AP_AXIMM_113_ARCACHE;
            assign ap_ARPROT[113] = AP_AXIMM_113_ARPROT;
            assign ap_ARREGION[113] = AP_AXIMM_113_ARREGION;
            assign ap_ARQOS[113] = AP_AXIMM_113_ARQOS;
            assign ap_ARVALID[113] = AP_AXIMM_113_ARVALID;
            assign AP_AXIMM_113_ARREADY = ap_ARREADY[113];
            assign AP_AXIMM_113_RDATA = ap_RDATA[113][M_AXIMM_113_DATA_WIDTH-1:0];
            assign AP_AXIMM_113_RRESP = ap_RRESP[113];
            assign AP_AXIMM_113_RLAST = ap_RLAST[113];
            assign AP_AXIMM_113_RVALID = ap_RVALID[113];
            assign ap_RREADY[113] = AP_AXIMM_113_RREADY;
            assign M_AXIMM_113_AWADDR = dm_AWADDR[113][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_113_AWLEN = dm_AWLEN[113];
            assign M_AXIMM_113_AWSIZE = dm_AWSIZE[113];
            assign M_AXIMM_113_AWBURST = dm_AWBURST[113];
            assign M_AXIMM_113_AWLOCK = dm_AWLOCK[113];
            assign M_AXIMM_113_AWCACHE = dm_AWCACHE[113];
            assign M_AXIMM_113_AWPROT = dm_AWPROT[113];
            assign M_AXIMM_113_AWREGION = dm_AWREGION[113];
            assign M_AXIMM_113_AWQOS = dm_AWQOS[113];
            assign M_AXIMM_113_AWVALID = dm_AWVALID[113];
            assign dm_AWREADY[113] = M_AXIMM_113_AWREADY;
            assign M_AXIMM_113_WDATA = dm_WDATA[113][M_AXIMM_113_DATA_WIDTH-1:0];
            assign M_AXIMM_113_WSTRB = dm_WSTRB[113][M_AXIMM_113_DATA_WIDTH/8-1:0];
            assign M_AXIMM_113_WLAST = dm_WLAST[113];
            assign M_AXIMM_113_WVALID = dm_WVALID[113];
            assign dm_WREADY[113] = M_AXIMM_113_WREADY;
            assign dm_BRESP[113] = M_AXIMM_113_BRESP;
            assign dm_BVALID[113] = M_AXIMM_113_BVALID;
            assign M_AXIMM_113_BREADY = dm_BREADY[113];
            assign M_AXIMM_113_ARADDR = dm_ARADDR[113][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_113_ARLEN = dm_ARLEN[113];
            assign M_AXIMM_113_ARSIZE = dm_ARSIZE[113];
            assign M_AXIMM_113_ARBURST = dm_ARBURST[113];
            assign M_AXIMM_113_ARLOCK = dm_ARLOCK[113];
            assign M_AXIMM_113_ARCACHE = dm_ARCACHE[113];
            assign M_AXIMM_113_ARPROT = dm_ARPROT[113];
            assign M_AXIMM_113_ARREGION = dm_ARREGION[113];
            assign M_AXIMM_113_ARQOS = dm_ARQOS[113];
            assign M_AXIMM_113_ARVALID = dm_ARVALID[113];
            assign dm_ARREADY[113] = M_AXIMM_113_ARREADY;
            assign dm_RDATA[113][M_AXIMM_113_DATA_WIDTH-1:0] = M_AXIMM_113_RDATA;
            assign dm_RRESP[113] = M_AXIMM_113_RRESP;
            assign dm_RLAST[113] = M_AXIMM_113_RLAST;
            assign dm_RVALID[113] = M_AXIMM_113_RVALID;
            assign M_AXIMM_113_RREADY = dm_RREADY[113];
        end
        if(C_NUM_AXIMMs > 114) begin
            assign ap_AWADDR[114][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_114_AWADDR;
            assign ap_AWLEN[114] = AP_AXIMM_114_AWLEN;
            assign ap_AWSIZE[114] = AP_AXIMM_114_AWSIZE;
            assign ap_AWBURST[114] = AP_AXIMM_114_AWBURST;
            assign ap_AWLOCK[114] = AP_AXIMM_114_AWLOCK;
            assign ap_AWCACHE[114] = AP_AXIMM_114_AWCACHE;
            assign ap_AWPROT[114] = AP_AXIMM_114_AWPROT;
            assign ap_AWREGION[114] = AP_AXIMM_114_AWREGION;
            assign ap_AWQOS[114] = AP_AXIMM_114_AWQOS;
            assign ap_AWVALID[114] = AP_AXIMM_114_AWVALID;
            assign AP_AXIMM_114_AWREADY = ap_AWREADY[114];
            assign ap_WDATA[114][M_AXIMM_114_DATA_WIDTH-1:0] = AP_AXIMM_114_WDATA;
            assign ap_WSTRB[114][M_AXIMM_114_DATA_WIDTH/8-1:0] = AP_AXIMM_114_WSTRB;
            assign ap_WLAST[114] = AP_AXIMM_114_WLAST;
            assign ap_WVALID[114] = AP_AXIMM_114_WVALID;
            assign AP_AXIMM_114_WREADY = ap_WREADY[114];
            assign AP_AXIMM_114_BRESP = ap_BRESP[114];
            assign AP_AXIMM_114_BVALID = ap_BVALID[114];
            assign ap_BREADY[114] = AP_AXIMM_114_BREADY;
            assign ap_ARADDR[114][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_114_ARADDR;
            assign ap_ARLEN[114] = AP_AXIMM_114_ARLEN;
            assign ap_ARSIZE[114] = AP_AXIMM_114_ARSIZE;
            assign ap_ARBURST[114] = AP_AXIMM_114_ARBURST;
            assign ap_ARLOCK[114] = AP_AXIMM_114_ARLOCK;
            assign ap_ARCACHE[114] = AP_AXIMM_114_ARCACHE;
            assign ap_ARPROT[114] = AP_AXIMM_114_ARPROT;
            assign ap_ARREGION[114] = AP_AXIMM_114_ARREGION;
            assign ap_ARQOS[114] = AP_AXIMM_114_ARQOS;
            assign ap_ARVALID[114] = AP_AXIMM_114_ARVALID;
            assign AP_AXIMM_114_ARREADY = ap_ARREADY[114];
            assign AP_AXIMM_114_RDATA = ap_RDATA[114][M_AXIMM_114_DATA_WIDTH-1:0];
            assign AP_AXIMM_114_RRESP = ap_RRESP[114];
            assign AP_AXIMM_114_RLAST = ap_RLAST[114];
            assign AP_AXIMM_114_RVALID = ap_RVALID[114];
            assign ap_RREADY[114] = AP_AXIMM_114_RREADY;
            assign M_AXIMM_114_AWADDR = dm_AWADDR[114][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_114_AWLEN = dm_AWLEN[114];
            assign M_AXIMM_114_AWSIZE = dm_AWSIZE[114];
            assign M_AXIMM_114_AWBURST = dm_AWBURST[114];
            assign M_AXIMM_114_AWLOCK = dm_AWLOCK[114];
            assign M_AXIMM_114_AWCACHE = dm_AWCACHE[114];
            assign M_AXIMM_114_AWPROT = dm_AWPROT[114];
            assign M_AXIMM_114_AWREGION = dm_AWREGION[114];
            assign M_AXIMM_114_AWQOS = dm_AWQOS[114];
            assign M_AXIMM_114_AWVALID = dm_AWVALID[114];
            assign dm_AWREADY[114] = M_AXIMM_114_AWREADY;
            assign M_AXIMM_114_WDATA = dm_WDATA[114][M_AXIMM_114_DATA_WIDTH-1:0];
            assign M_AXIMM_114_WSTRB = dm_WSTRB[114][M_AXIMM_114_DATA_WIDTH/8-1:0];
            assign M_AXIMM_114_WLAST = dm_WLAST[114];
            assign M_AXIMM_114_WVALID = dm_WVALID[114];
            assign dm_WREADY[114] = M_AXIMM_114_WREADY;
            assign dm_BRESP[114] = M_AXIMM_114_BRESP;
            assign dm_BVALID[114] = M_AXIMM_114_BVALID;
            assign M_AXIMM_114_BREADY = dm_BREADY[114];
            assign M_AXIMM_114_ARADDR = dm_ARADDR[114][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_114_ARLEN = dm_ARLEN[114];
            assign M_AXIMM_114_ARSIZE = dm_ARSIZE[114];
            assign M_AXIMM_114_ARBURST = dm_ARBURST[114];
            assign M_AXIMM_114_ARLOCK = dm_ARLOCK[114];
            assign M_AXIMM_114_ARCACHE = dm_ARCACHE[114];
            assign M_AXIMM_114_ARPROT = dm_ARPROT[114];
            assign M_AXIMM_114_ARREGION = dm_ARREGION[114];
            assign M_AXIMM_114_ARQOS = dm_ARQOS[114];
            assign M_AXIMM_114_ARVALID = dm_ARVALID[114];
            assign dm_ARREADY[114] = M_AXIMM_114_ARREADY;
            assign dm_RDATA[114][M_AXIMM_114_DATA_WIDTH-1:0] = M_AXIMM_114_RDATA;
            assign dm_RRESP[114] = M_AXIMM_114_RRESP;
            assign dm_RLAST[114] = M_AXIMM_114_RLAST;
            assign dm_RVALID[114] = M_AXIMM_114_RVALID;
            assign M_AXIMM_114_RREADY = dm_RREADY[114];
        end
        if(C_NUM_AXIMMs > 115) begin
            assign ap_AWADDR[115][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_115_AWADDR;
            assign ap_AWLEN[115] = AP_AXIMM_115_AWLEN;
            assign ap_AWSIZE[115] = AP_AXIMM_115_AWSIZE;
            assign ap_AWBURST[115] = AP_AXIMM_115_AWBURST;
            assign ap_AWLOCK[115] = AP_AXIMM_115_AWLOCK;
            assign ap_AWCACHE[115] = AP_AXIMM_115_AWCACHE;
            assign ap_AWPROT[115] = AP_AXIMM_115_AWPROT;
            assign ap_AWREGION[115] = AP_AXIMM_115_AWREGION;
            assign ap_AWQOS[115] = AP_AXIMM_115_AWQOS;
            assign ap_AWVALID[115] = AP_AXIMM_115_AWVALID;
            assign AP_AXIMM_115_AWREADY = ap_AWREADY[115];
            assign ap_WDATA[115][M_AXIMM_115_DATA_WIDTH-1:0] = AP_AXIMM_115_WDATA;
            assign ap_WSTRB[115][M_AXIMM_115_DATA_WIDTH/8-1:0] = AP_AXIMM_115_WSTRB;
            assign ap_WLAST[115] = AP_AXIMM_115_WLAST;
            assign ap_WVALID[115] = AP_AXIMM_115_WVALID;
            assign AP_AXIMM_115_WREADY = ap_WREADY[115];
            assign AP_AXIMM_115_BRESP = ap_BRESP[115];
            assign AP_AXIMM_115_BVALID = ap_BVALID[115];
            assign ap_BREADY[115] = AP_AXIMM_115_BREADY;
            assign ap_ARADDR[115][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_115_ARADDR;
            assign ap_ARLEN[115] = AP_AXIMM_115_ARLEN;
            assign ap_ARSIZE[115] = AP_AXIMM_115_ARSIZE;
            assign ap_ARBURST[115] = AP_AXIMM_115_ARBURST;
            assign ap_ARLOCK[115] = AP_AXIMM_115_ARLOCK;
            assign ap_ARCACHE[115] = AP_AXIMM_115_ARCACHE;
            assign ap_ARPROT[115] = AP_AXIMM_115_ARPROT;
            assign ap_ARREGION[115] = AP_AXIMM_115_ARREGION;
            assign ap_ARQOS[115] = AP_AXIMM_115_ARQOS;
            assign ap_ARVALID[115] = AP_AXIMM_115_ARVALID;
            assign AP_AXIMM_115_ARREADY = ap_ARREADY[115];
            assign AP_AXIMM_115_RDATA = ap_RDATA[115][M_AXIMM_115_DATA_WIDTH-1:0];
            assign AP_AXIMM_115_RRESP = ap_RRESP[115];
            assign AP_AXIMM_115_RLAST = ap_RLAST[115];
            assign AP_AXIMM_115_RVALID = ap_RVALID[115];
            assign ap_RREADY[115] = AP_AXIMM_115_RREADY;
            assign M_AXIMM_115_AWADDR = dm_AWADDR[115][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_115_AWLEN = dm_AWLEN[115];
            assign M_AXIMM_115_AWSIZE = dm_AWSIZE[115];
            assign M_AXIMM_115_AWBURST = dm_AWBURST[115];
            assign M_AXIMM_115_AWLOCK = dm_AWLOCK[115];
            assign M_AXIMM_115_AWCACHE = dm_AWCACHE[115];
            assign M_AXIMM_115_AWPROT = dm_AWPROT[115];
            assign M_AXIMM_115_AWREGION = dm_AWREGION[115];
            assign M_AXIMM_115_AWQOS = dm_AWQOS[115];
            assign M_AXIMM_115_AWVALID = dm_AWVALID[115];
            assign dm_AWREADY[115] = M_AXIMM_115_AWREADY;
            assign M_AXIMM_115_WDATA = dm_WDATA[115][M_AXIMM_115_DATA_WIDTH-1:0];
            assign M_AXIMM_115_WSTRB = dm_WSTRB[115][M_AXIMM_115_DATA_WIDTH/8-1:0];
            assign M_AXIMM_115_WLAST = dm_WLAST[115];
            assign M_AXIMM_115_WVALID = dm_WVALID[115];
            assign dm_WREADY[115] = M_AXIMM_115_WREADY;
            assign dm_BRESP[115] = M_AXIMM_115_BRESP;
            assign dm_BVALID[115] = M_AXIMM_115_BVALID;
            assign M_AXIMM_115_BREADY = dm_BREADY[115];
            assign M_AXIMM_115_ARADDR = dm_ARADDR[115][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_115_ARLEN = dm_ARLEN[115];
            assign M_AXIMM_115_ARSIZE = dm_ARSIZE[115];
            assign M_AXIMM_115_ARBURST = dm_ARBURST[115];
            assign M_AXIMM_115_ARLOCK = dm_ARLOCK[115];
            assign M_AXIMM_115_ARCACHE = dm_ARCACHE[115];
            assign M_AXIMM_115_ARPROT = dm_ARPROT[115];
            assign M_AXIMM_115_ARREGION = dm_ARREGION[115];
            assign M_AXIMM_115_ARQOS = dm_ARQOS[115];
            assign M_AXIMM_115_ARVALID = dm_ARVALID[115];
            assign dm_ARREADY[115] = M_AXIMM_115_ARREADY;
            assign dm_RDATA[115][M_AXIMM_115_DATA_WIDTH-1:0] = M_AXIMM_115_RDATA;
            assign dm_RRESP[115] = M_AXIMM_115_RRESP;
            assign dm_RLAST[115] = M_AXIMM_115_RLAST;
            assign dm_RVALID[115] = M_AXIMM_115_RVALID;
            assign M_AXIMM_115_RREADY = dm_RREADY[115];
        end
        if(C_NUM_AXIMMs > 116) begin
            assign ap_AWADDR[116][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_116_AWADDR;
            assign ap_AWLEN[116] = AP_AXIMM_116_AWLEN;
            assign ap_AWSIZE[116] = AP_AXIMM_116_AWSIZE;
            assign ap_AWBURST[116] = AP_AXIMM_116_AWBURST;
            assign ap_AWLOCK[116] = AP_AXIMM_116_AWLOCK;
            assign ap_AWCACHE[116] = AP_AXIMM_116_AWCACHE;
            assign ap_AWPROT[116] = AP_AXIMM_116_AWPROT;
            assign ap_AWREGION[116] = AP_AXIMM_116_AWREGION;
            assign ap_AWQOS[116] = AP_AXIMM_116_AWQOS;
            assign ap_AWVALID[116] = AP_AXIMM_116_AWVALID;
            assign AP_AXIMM_116_AWREADY = ap_AWREADY[116];
            assign ap_WDATA[116][M_AXIMM_116_DATA_WIDTH-1:0] = AP_AXIMM_116_WDATA;
            assign ap_WSTRB[116][M_AXIMM_116_DATA_WIDTH/8-1:0] = AP_AXIMM_116_WSTRB;
            assign ap_WLAST[116] = AP_AXIMM_116_WLAST;
            assign ap_WVALID[116] = AP_AXIMM_116_WVALID;
            assign AP_AXIMM_116_WREADY = ap_WREADY[116];
            assign AP_AXIMM_116_BRESP = ap_BRESP[116];
            assign AP_AXIMM_116_BVALID = ap_BVALID[116];
            assign ap_BREADY[116] = AP_AXIMM_116_BREADY;
            assign ap_ARADDR[116][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_116_ARADDR;
            assign ap_ARLEN[116] = AP_AXIMM_116_ARLEN;
            assign ap_ARSIZE[116] = AP_AXIMM_116_ARSIZE;
            assign ap_ARBURST[116] = AP_AXIMM_116_ARBURST;
            assign ap_ARLOCK[116] = AP_AXIMM_116_ARLOCK;
            assign ap_ARCACHE[116] = AP_AXIMM_116_ARCACHE;
            assign ap_ARPROT[116] = AP_AXIMM_116_ARPROT;
            assign ap_ARREGION[116] = AP_AXIMM_116_ARREGION;
            assign ap_ARQOS[116] = AP_AXIMM_116_ARQOS;
            assign ap_ARVALID[116] = AP_AXIMM_116_ARVALID;
            assign AP_AXIMM_116_ARREADY = ap_ARREADY[116];
            assign AP_AXIMM_116_RDATA = ap_RDATA[116][M_AXIMM_116_DATA_WIDTH-1:0];
            assign AP_AXIMM_116_RRESP = ap_RRESP[116];
            assign AP_AXIMM_116_RLAST = ap_RLAST[116];
            assign AP_AXIMM_116_RVALID = ap_RVALID[116];
            assign ap_RREADY[116] = AP_AXIMM_116_RREADY;
            assign M_AXIMM_116_AWADDR = dm_AWADDR[116][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_116_AWLEN = dm_AWLEN[116];
            assign M_AXIMM_116_AWSIZE = dm_AWSIZE[116];
            assign M_AXIMM_116_AWBURST = dm_AWBURST[116];
            assign M_AXIMM_116_AWLOCK = dm_AWLOCK[116];
            assign M_AXIMM_116_AWCACHE = dm_AWCACHE[116];
            assign M_AXIMM_116_AWPROT = dm_AWPROT[116];
            assign M_AXIMM_116_AWREGION = dm_AWREGION[116];
            assign M_AXIMM_116_AWQOS = dm_AWQOS[116];
            assign M_AXIMM_116_AWVALID = dm_AWVALID[116];
            assign dm_AWREADY[116] = M_AXIMM_116_AWREADY;
            assign M_AXIMM_116_WDATA = dm_WDATA[116][M_AXIMM_116_DATA_WIDTH-1:0];
            assign M_AXIMM_116_WSTRB = dm_WSTRB[116][M_AXIMM_116_DATA_WIDTH/8-1:0];
            assign M_AXIMM_116_WLAST = dm_WLAST[116];
            assign M_AXIMM_116_WVALID = dm_WVALID[116];
            assign dm_WREADY[116] = M_AXIMM_116_WREADY;
            assign dm_BRESP[116] = M_AXIMM_116_BRESP;
            assign dm_BVALID[116] = M_AXIMM_116_BVALID;
            assign M_AXIMM_116_BREADY = dm_BREADY[116];
            assign M_AXIMM_116_ARADDR = dm_ARADDR[116][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_116_ARLEN = dm_ARLEN[116];
            assign M_AXIMM_116_ARSIZE = dm_ARSIZE[116];
            assign M_AXIMM_116_ARBURST = dm_ARBURST[116];
            assign M_AXIMM_116_ARLOCK = dm_ARLOCK[116];
            assign M_AXIMM_116_ARCACHE = dm_ARCACHE[116];
            assign M_AXIMM_116_ARPROT = dm_ARPROT[116];
            assign M_AXIMM_116_ARREGION = dm_ARREGION[116];
            assign M_AXIMM_116_ARQOS = dm_ARQOS[116];
            assign M_AXIMM_116_ARVALID = dm_ARVALID[116];
            assign dm_ARREADY[116] = M_AXIMM_116_ARREADY;
            assign dm_RDATA[116][M_AXIMM_116_DATA_WIDTH-1:0] = M_AXIMM_116_RDATA;
            assign dm_RRESP[116] = M_AXIMM_116_RRESP;
            assign dm_RLAST[116] = M_AXIMM_116_RLAST;
            assign dm_RVALID[116] = M_AXIMM_116_RVALID;
            assign M_AXIMM_116_RREADY = dm_RREADY[116];
        end
        if(C_NUM_AXIMMs > 117) begin
            assign ap_AWADDR[117][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_117_AWADDR;
            assign ap_AWLEN[117] = AP_AXIMM_117_AWLEN;
            assign ap_AWSIZE[117] = AP_AXIMM_117_AWSIZE;
            assign ap_AWBURST[117] = AP_AXIMM_117_AWBURST;
            assign ap_AWLOCK[117] = AP_AXIMM_117_AWLOCK;
            assign ap_AWCACHE[117] = AP_AXIMM_117_AWCACHE;
            assign ap_AWPROT[117] = AP_AXIMM_117_AWPROT;
            assign ap_AWREGION[117] = AP_AXIMM_117_AWREGION;
            assign ap_AWQOS[117] = AP_AXIMM_117_AWQOS;
            assign ap_AWVALID[117] = AP_AXIMM_117_AWVALID;
            assign AP_AXIMM_117_AWREADY = ap_AWREADY[117];
            assign ap_WDATA[117][M_AXIMM_117_DATA_WIDTH-1:0] = AP_AXIMM_117_WDATA;
            assign ap_WSTRB[117][M_AXIMM_117_DATA_WIDTH/8-1:0] = AP_AXIMM_117_WSTRB;
            assign ap_WLAST[117] = AP_AXIMM_117_WLAST;
            assign ap_WVALID[117] = AP_AXIMM_117_WVALID;
            assign AP_AXIMM_117_WREADY = ap_WREADY[117];
            assign AP_AXIMM_117_BRESP = ap_BRESP[117];
            assign AP_AXIMM_117_BVALID = ap_BVALID[117];
            assign ap_BREADY[117] = AP_AXIMM_117_BREADY;
            assign ap_ARADDR[117][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_117_ARADDR;
            assign ap_ARLEN[117] = AP_AXIMM_117_ARLEN;
            assign ap_ARSIZE[117] = AP_AXIMM_117_ARSIZE;
            assign ap_ARBURST[117] = AP_AXIMM_117_ARBURST;
            assign ap_ARLOCK[117] = AP_AXIMM_117_ARLOCK;
            assign ap_ARCACHE[117] = AP_AXIMM_117_ARCACHE;
            assign ap_ARPROT[117] = AP_AXIMM_117_ARPROT;
            assign ap_ARREGION[117] = AP_AXIMM_117_ARREGION;
            assign ap_ARQOS[117] = AP_AXIMM_117_ARQOS;
            assign ap_ARVALID[117] = AP_AXIMM_117_ARVALID;
            assign AP_AXIMM_117_ARREADY = ap_ARREADY[117];
            assign AP_AXIMM_117_RDATA = ap_RDATA[117][M_AXIMM_117_DATA_WIDTH-1:0];
            assign AP_AXIMM_117_RRESP = ap_RRESP[117];
            assign AP_AXIMM_117_RLAST = ap_RLAST[117];
            assign AP_AXIMM_117_RVALID = ap_RVALID[117];
            assign ap_RREADY[117] = AP_AXIMM_117_RREADY;
            assign M_AXIMM_117_AWADDR = dm_AWADDR[117][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_117_AWLEN = dm_AWLEN[117];
            assign M_AXIMM_117_AWSIZE = dm_AWSIZE[117];
            assign M_AXIMM_117_AWBURST = dm_AWBURST[117];
            assign M_AXIMM_117_AWLOCK = dm_AWLOCK[117];
            assign M_AXIMM_117_AWCACHE = dm_AWCACHE[117];
            assign M_AXIMM_117_AWPROT = dm_AWPROT[117];
            assign M_AXIMM_117_AWREGION = dm_AWREGION[117];
            assign M_AXIMM_117_AWQOS = dm_AWQOS[117];
            assign M_AXIMM_117_AWVALID = dm_AWVALID[117];
            assign dm_AWREADY[117] = M_AXIMM_117_AWREADY;
            assign M_AXIMM_117_WDATA = dm_WDATA[117][M_AXIMM_117_DATA_WIDTH-1:0];
            assign M_AXIMM_117_WSTRB = dm_WSTRB[117][M_AXIMM_117_DATA_WIDTH/8-1:0];
            assign M_AXIMM_117_WLAST = dm_WLAST[117];
            assign M_AXIMM_117_WVALID = dm_WVALID[117];
            assign dm_WREADY[117] = M_AXIMM_117_WREADY;
            assign dm_BRESP[117] = M_AXIMM_117_BRESP;
            assign dm_BVALID[117] = M_AXIMM_117_BVALID;
            assign M_AXIMM_117_BREADY = dm_BREADY[117];
            assign M_AXIMM_117_ARADDR = dm_ARADDR[117][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_117_ARLEN = dm_ARLEN[117];
            assign M_AXIMM_117_ARSIZE = dm_ARSIZE[117];
            assign M_AXIMM_117_ARBURST = dm_ARBURST[117];
            assign M_AXIMM_117_ARLOCK = dm_ARLOCK[117];
            assign M_AXIMM_117_ARCACHE = dm_ARCACHE[117];
            assign M_AXIMM_117_ARPROT = dm_ARPROT[117];
            assign M_AXIMM_117_ARREGION = dm_ARREGION[117];
            assign M_AXIMM_117_ARQOS = dm_ARQOS[117];
            assign M_AXIMM_117_ARVALID = dm_ARVALID[117];
            assign dm_ARREADY[117] = M_AXIMM_117_ARREADY;
            assign dm_RDATA[117][M_AXIMM_117_DATA_WIDTH-1:0] = M_AXIMM_117_RDATA;
            assign dm_RRESP[117] = M_AXIMM_117_RRESP;
            assign dm_RLAST[117] = M_AXIMM_117_RLAST;
            assign dm_RVALID[117] = M_AXIMM_117_RVALID;
            assign M_AXIMM_117_RREADY = dm_RREADY[117];
        end
        if(C_NUM_AXIMMs > 118) begin
            assign ap_AWADDR[118][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_118_AWADDR;
            assign ap_AWLEN[118] = AP_AXIMM_118_AWLEN;
            assign ap_AWSIZE[118] = AP_AXIMM_118_AWSIZE;
            assign ap_AWBURST[118] = AP_AXIMM_118_AWBURST;
            assign ap_AWLOCK[118] = AP_AXIMM_118_AWLOCK;
            assign ap_AWCACHE[118] = AP_AXIMM_118_AWCACHE;
            assign ap_AWPROT[118] = AP_AXIMM_118_AWPROT;
            assign ap_AWREGION[118] = AP_AXIMM_118_AWREGION;
            assign ap_AWQOS[118] = AP_AXIMM_118_AWQOS;
            assign ap_AWVALID[118] = AP_AXIMM_118_AWVALID;
            assign AP_AXIMM_118_AWREADY = ap_AWREADY[118];
            assign ap_WDATA[118][M_AXIMM_118_DATA_WIDTH-1:0] = AP_AXIMM_118_WDATA;
            assign ap_WSTRB[118][M_AXIMM_118_DATA_WIDTH/8-1:0] = AP_AXIMM_118_WSTRB;
            assign ap_WLAST[118] = AP_AXIMM_118_WLAST;
            assign ap_WVALID[118] = AP_AXIMM_118_WVALID;
            assign AP_AXIMM_118_WREADY = ap_WREADY[118];
            assign AP_AXIMM_118_BRESP = ap_BRESP[118];
            assign AP_AXIMM_118_BVALID = ap_BVALID[118];
            assign ap_BREADY[118] = AP_AXIMM_118_BREADY;
            assign ap_ARADDR[118][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_118_ARADDR;
            assign ap_ARLEN[118] = AP_AXIMM_118_ARLEN;
            assign ap_ARSIZE[118] = AP_AXIMM_118_ARSIZE;
            assign ap_ARBURST[118] = AP_AXIMM_118_ARBURST;
            assign ap_ARLOCK[118] = AP_AXIMM_118_ARLOCK;
            assign ap_ARCACHE[118] = AP_AXIMM_118_ARCACHE;
            assign ap_ARPROT[118] = AP_AXIMM_118_ARPROT;
            assign ap_ARREGION[118] = AP_AXIMM_118_ARREGION;
            assign ap_ARQOS[118] = AP_AXIMM_118_ARQOS;
            assign ap_ARVALID[118] = AP_AXIMM_118_ARVALID;
            assign AP_AXIMM_118_ARREADY = ap_ARREADY[118];
            assign AP_AXIMM_118_RDATA = ap_RDATA[118][M_AXIMM_118_DATA_WIDTH-1:0];
            assign AP_AXIMM_118_RRESP = ap_RRESP[118];
            assign AP_AXIMM_118_RLAST = ap_RLAST[118];
            assign AP_AXIMM_118_RVALID = ap_RVALID[118];
            assign ap_RREADY[118] = AP_AXIMM_118_RREADY;
            assign M_AXIMM_118_AWADDR = dm_AWADDR[118][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_118_AWLEN = dm_AWLEN[118];
            assign M_AXIMM_118_AWSIZE = dm_AWSIZE[118];
            assign M_AXIMM_118_AWBURST = dm_AWBURST[118];
            assign M_AXIMM_118_AWLOCK = dm_AWLOCK[118];
            assign M_AXIMM_118_AWCACHE = dm_AWCACHE[118];
            assign M_AXIMM_118_AWPROT = dm_AWPROT[118];
            assign M_AXIMM_118_AWREGION = dm_AWREGION[118];
            assign M_AXIMM_118_AWQOS = dm_AWQOS[118];
            assign M_AXIMM_118_AWVALID = dm_AWVALID[118];
            assign dm_AWREADY[118] = M_AXIMM_118_AWREADY;
            assign M_AXIMM_118_WDATA = dm_WDATA[118][M_AXIMM_118_DATA_WIDTH-1:0];
            assign M_AXIMM_118_WSTRB = dm_WSTRB[118][M_AXIMM_118_DATA_WIDTH/8-1:0];
            assign M_AXIMM_118_WLAST = dm_WLAST[118];
            assign M_AXIMM_118_WVALID = dm_WVALID[118];
            assign dm_WREADY[118] = M_AXIMM_118_WREADY;
            assign dm_BRESP[118] = M_AXIMM_118_BRESP;
            assign dm_BVALID[118] = M_AXIMM_118_BVALID;
            assign M_AXIMM_118_BREADY = dm_BREADY[118];
            assign M_AXIMM_118_ARADDR = dm_ARADDR[118][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_118_ARLEN = dm_ARLEN[118];
            assign M_AXIMM_118_ARSIZE = dm_ARSIZE[118];
            assign M_AXIMM_118_ARBURST = dm_ARBURST[118];
            assign M_AXIMM_118_ARLOCK = dm_ARLOCK[118];
            assign M_AXIMM_118_ARCACHE = dm_ARCACHE[118];
            assign M_AXIMM_118_ARPROT = dm_ARPROT[118];
            assign M_AXIMM_118_ARREGION = dm_ARREGION[118];
            assign M_AXIMM_118_ARQOS = dm_ARQOS[118];
            assign M_AXIMM_118_ARVALID = dm_ARVALID[118];
            assign dm_ARREADY[118] = M_AXIMM_118_ARREADY;
            assign dm_RDATA[118][M_AXIMM_118_DATA_WIDTH-1:0] = M_AXIMM_118_RDATA;
            assign dm_RRESP[118] = M_AXIMM_118_RRESP;
            assign dm_RLAST[118] = M_AXIMM_118_RLAST;
            assign dm_RVALID[118] = M_AXIMM_118_RVALID;
            assign M_AXIMM_118_RREADY = dm_RREADY[118];
        end
        if(C_NUM_AXIMMs > 119) begin
            assign ap_AWADDR[119][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_119_AWADDR;
            assign ap_AWLEN[119] = AP_AXIMM_119_AWLEN;
            assign ap_AWSIZE[119] = AP_AXIMM_119_AWSIZE;
            assign ap_AWBURST[119] = AP_AXIMM_119_AWBURST;
            assign ap_AWLOCK[119] = AP_AXIMM_119_AWLOCK;
            assign ap_AWCACHE[119] = AP_AXIMM_119_AWCACHE;
            assign ap_AWPROT[119] = AP_AXIMM_119_AWPROT;
            assign ap_AWREGION[119] = AP_AXIMM_119_AWREGION;
            assign ap_AWQOS[119] = AP_AXIMM_119_AWQOS;
            assign ap_AWVALID[119] = AP_AXIMM_119_AWVALID;
            assign AP_AXIMM_119_AWREADY = ap_AWREADY[119];
            assign ap_WDATA[119][M_AXIMM_119_DATA_WIDTH-1:0] = AP_AXIMM_119_WDATA;
            assign ap_WSTRB[119][M_AXIMM_119_DATA_WIDTH/8-1:0] = AP_AXIMM_119_WSTRB;
            assign ap_WLAST[119] = AP_AXIMM_119_WLAST;
            assign ap_WVALID[119] = AP_AXIMM_119_WVALID;
            assign AP_AXIMM_119_WREADY = ap_WREADY[119];
            assign AP_AXIMM_119_BRESP = ap_BRESP[119];
            assign AP_AXIMM_119_BVALID = ap_BVALID[119];
            assign ap_BREADY[119] = AP_AXIMM_119_BREADY;
            assign ap_ARADDR[119][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_119_ARADDR;
            assign ap_ARLEN[119] = AP_AXIMM_119_ARLEN;
            assign ap_ARSIZE[119] = AP_AXIMM_119_ARSIZE;
            assign ap_ARBURST[119] = AP_AXIMM_119_ARBURST;
            assign ap_ARLOCK[119] = AP_AXIMM_119_ARLOCK;
            assign ap_ARCACHE[119] = AP_AXIMM_119_ARCACHE;
            assign ap_ARPROT[119] = AP_AXIMM_119_ARPROT;
            assign ap_ARREGION[119] = AP_AXIMM_119_ARREGION;
            assign ap_ARQOS[119] = AP_AXIMM_119_ARQOS;
            assign ap_ARVALID[119] = AP_AXIMM_119_ARVALID;
            assign AP_AXIMM_119_ARREADY = ap_ARREADY[119];
            assign AP_AXIMM_119_RDATA = ap_RDATA[119][M_AXIMM_119_DATA_WIDTH-1:0];
            assign AP_AXIMM_119_RRESP = ap_RRESP[119];
            assign AP_AXIMM_119_RLAST = ap_RLAST[119];
            assign AP_AXIMM_119_RVALID = ap_RVALID[119];
            assign ap_RREADY[119] = AP_AXIMM_119_RREADY;
            assign M_AXIMM_119_AWADDR = dm_AWADDR[119][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_119_AWLEN = dm_AWLEN[119];
            assign M_AXIMM_119_AWSIZE = dm_AWSIZE[119];
            assign M_AXIMM_119_AWBURST = dm_AWBURST[119];
            assign M_AXIMM_119_AWLOCK = dm_AWLOCK[119];
            assign M_AXIMM_119_AWCACHE = dm_AWCACHE[119];
            assign M_AXIMM_119_AWPROT = dm_AWPROT[119];
            assign M_AXIMM_119_AWREGION = dm_AWREGION[119];
            assign M_AXIMM_119_AWQOS = dm_AWQOS[119];
            assign M_AXIMM_119_AWVALID = dm_AWVALID[119];
            assign dm_AWREADY[119] = M_AXIMM_119_AWREADY;
            assign M_AXIMM_119_WDATA = dm_WDATA[119][M_AXIMM_119_DATA_WIDTH-1:0];
            assign M_AXIMM_119_WSTRB = dm_WSTRB[119][M_AXIMM_119_DATA_WIDTH/8-1:0];
            assign M_AXIMM_119_WLAST = dm_WLAST[119];
            assign M_AXIMM_119_WVALID = dm_WVALID[119];
            assign dm_WREADY[119] = M_AXIMM_119_WREADY;
            assign dm_BRESP[119] = M_AXIMM_119_BRESP;
            assign dm_BVALID[119] = M_AXIMM_119_BVALID;
            assign M_AXIMM_119_BREADY = dm_BREADY[119];
            assign M_AXIMM_119_ARADDR = dm_ARADDR[119][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_119_ARLEN = dm_ARLEN[119];
            assign M_AXIMM_119_ARSIZE = dm_ARSIZE[119];
            assign M_AXIMM_119_ARBURST = dm_ARBURST[119];
            assign M_AXIMM_119_ARLOCK = dm_ARLOCK[119];
            assign M_AXIMM_119_ARCACHE = dm_ARCACHE[119];
            assign M_AXIMM_119_ARPROT = dm_ARPROT[119];
            assign M_AXIMM_119_ARREGION = dm_ARREGION[119];
            assign M_AXIMM_119_ARQOS = dm_ARQOS[119];
            assign M_AXIMM_119_ARVALID = dm_ARVALID[119];
            assign dm_ARREADY[119] = M_AXIMM_119_ARREADY;
            assign dm_RDATA[119][M_AXIMM_119_DATA_WIDTH-1:0] = M_AXIMM_119_RDATA;
            assign dm_RRESP[119] = M_AXIMM_119_RRESP;
            assign dm_RLAST[119] = M_AXIMM_119_RLAST;
            assign dm_RVALID[119] = M_AXIMM_119_RVALID;
            assign M_AXIMM_119_RREADY = dm_RREADY[119];
        end
        if(C_NUM_AXIMMs > 120) begin
            assign ap_AWADDR[120][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_120_AWADDR;
            assign ap_AWLEN[120] = AP_AXIMM_120_AWLEN;
            assign ap_AWSIZE[120] = AP_AXIMM_120_AWSIZE;
            assign ap_AWBURST[120] = AP_AXIMM_120_AWBURST;
            assign ap_AWLOCK[120] = AP_AXIMM_120_AWLOCK;
            assign ap_AWCACHE[120] = AP_AXIMM_120_AWCACHE;
            assign ap_AWPROT[120] = AP_AXIMM_120_AWPROT;
            assign ap_AWREGION[120] = AP_AXIMM_120_AWREGION;
            assign ap_AWQOS[120] = AP_AXIMM_120_AWQOS;
            assign ap_AWVALID[120] = AP_AXIMM_120_AWVALID;
            assign AP_AXIMM_120_AWREADY = ap_AWREADY[120];
            assign ap_WDATA[120][M_AXIMM_120_DATA_WIDTH-1:0] = AP_AXIMM_120_WDATA;
            assign ap_WSTRB[120][M_AXIMM_120_DATA_WIDTH/8-1:0] = AP_AXIMM_120_WSTRB;
            assign ap_WLAST[120] = AP_AXIMM_120_WLAST;
            assign ap_WVALID[120] = AP_AXIMM_120_WVALID;
            assign AP_AXIMM_120_WREADY = ap_WREADY[120];
            assign AP_AXIMM_120_BRESP = ap_BRESP[120];
            assign AP_AXIMM_120_BVALID = ap_BVALID[120];
            assign ap_BREADY[120] = AP_AXIMM_120_BREADY;
            assign ap_ARADDR[120][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_120_ARADDR;
            assign ap_ARLEN[120] = AP_AXIMM_120_ARLEN;
            assign ap_ARSIZE[120] = AP_AXIMM_120_ARSIZE;
            assign ap_ARBURST[120] = AP_AXIMM_120_ARBURST;
            assign ap_ARLOCK[120] = AP_AXIMM_120_ARLOCK;
            assign ap_ARCACHE[120] = AP_AXIMM_120_ARCACHE;
            assign ap_ARPROT[120] = AP_AXIMM_120_ARPROT;
            assign ap_ARREGION[120] = AP_AXIMM_120_ARREGION;
            assign ap_ARQOS[120] = AP_AXIMM_120_ARQOS;
            assign ap_ARVALID[120] = AP_AXIMM_120_ARVALID;
            assign AP_AXIMM_120_ARREADY = ap_ARREADY[120];
            assign AP_AXIMM_120_RDATA = ap_RDATA[120][M_AXIMM_120_DATA_WIDTH-1:0];
            assign AP_AXIMM_120_RRESP = ap_RRESP[120];
            assign AP_AXIMM_120_RLAST = ap_RLAST[120];
            assign AP_AXIMM_120_RVALID = ap_RVALID[120];
            assign ap_RREADY[120] = AP_AXIMM_120_RREADY;
            assign M_AXIMM_120_AWADDR = dm_AWADDR[120][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_120_AWLEN = dm_AWLEN[120];
            assign M_AXIMM_120_AWSIZE = dm_AWSIZE[120];
            assign M_AXIMM_120_AWBURST = dm_AWBURST[120];
            assign M_AXIMM_120_AWLOCK = dm_AWLOCK[120];
            assign M_AXIMM_120_AWCACHE = dm_AWCACHE[120];
            assign M_AXIMM_120_AWPROT = dm_AWPROT[120];
            assign M_AXIMM_120_AWREGION = dm_AWREGION[120];
            assign M_AXIMM_120_AWQOS = dm_AWQOS[120];
            assign M_AXIMM_120_AWVALID = dm_AWVALID[120];
            assign dm_AWREADY[120] = M_AXIMM_120_AWREADY;
            assign M_AXIMM_120_WDATA = dm_WDATA[120][M_AXIMM_120_DATA_WIDTH-1:0];
            assign M_AXIMM_120_WSTRB = dm_WSTRB[120][M_AXIMM_120_DATA_WIDTH/8-1:0];
            assign M_AXIMM_120_WLAST = dm_WLAST[120];
            assign M_AXIMM_120_WVALID = dm_WVALID[120];
            assign dm_WREADY[120] = M_AXIMM_120_WREADY;
            assign dm_BRESP[120] = M_AXIMM_120_BRESP;
            assign dm_BVALID[120] = M_AXIMM_120_BVALID;
            assign M_AXIMM_120_BREADY = dm_BREADY[120];
            assign M_AXIMM_120_ARADDR = dm_ARADDR[120][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_120_ARLEN = dm_ARLEN[120];
            assign M_AXIMM_120_ARSIZE = dm_ARSIZE[120];
            assign M_AXIMM_120_ARBURST = dm_ARBURST[120];
            assign M_AXIMM_120_ARLOCK = dm_ARLOCK[120];
            assign M_AXIMM_120_ARCACHE = dm_ARCACHE[120];
            assign M_AXIMM_120_ARPROT = dm_ARPROT[120];
            assign M_AXIMM_120_ARREGION = dm_ARREGION[120];
            assign M_AXIMM_120_ARQOS = dm_ARQOS[120];
            assign M_AXIMM_120_ARVALID = dm_ARVALID[120];
            assign dm_ARREADY[120] = M_AXIMM_120_ARREADY;
            assign dm_RDATA[120][M_AXIMM_120_DATA_WIDTH-1:0] = M_AXIMM_120_RDATA;
            assign dm_RRESP[120] = M_AXIMM_120_RRESP;
            assign dm_RLAST[120] = M_AXIMM_120_RLAST;
            assign dm_RVALID[120] = M_AXIMM_120_RVALID;
            assign M_AXIMM_120_RREADY = dm_RREADY[120];
        end
        if(C_NUM_AXIMMs > 121) begin
            assign ap_AWADDR[121][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_121_AWADDR;
            assign ap_AWLEN[121] = AP_AXIMM_121_AWLEN;
            assign ap_AWSIZE[121] = AP_AXIMM_121_AWSIZE;
            assign ap_AWBURST[121] = AP_AXIMM_121_AWBURST;
            assign ap_AWLOCK[121] = AP_AXIMM_121_AWLOCK;
            assign ap_AWCACHE[121] = AP_AXIMM_121_AWCACHE;
            assign ap_AWPROT[121] = AP_AXIMM_121_AWPROT;
            assign ap_AWREGION[121] = AP_AXIMM_121_AWREGION;
            assign ap_AWQOS[121] = AP_AXIMM_121_AWQOS;
            assign ap_AWVALID[121] = AP_AXIMM_121_AWVALID;
            assign AP_AXIMM_121_AWREADY = ap_AWREADY[121];
            assign ap_WDATA[121][M_AXIMM_121_DATA_WIDTH-1:0] = AP_AXIMM_121_WDATA;
            assign ap_WSTRB[121][M_AXIMM_121_DATA_WIDTH/8-1:0] = AP_AXIMM_121_WSTRB;
            assign ap_WLAST[121] = AP_AXIMM_121_WLAST;
            assign ap_WVALID[121] = AP_AXIMM_121_WVALID;
            assign AP_AXIMM_121_WREADY = ap_WREADY[121];
            assign AP_AXIMM_121_BRESP = ap_BRESP[121];
            assign AP_AXIMM_121_BVALID = ap_BVALID[121];
            assign ap_BREADY[121] = AP_AXIMM_121_BREADY;
            assign ap_ARADDR[121][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_121_ARADDR;
            assign ap_ARLEN[121] = AP_AXIMM_121_ARLEN;
            assign ap_ARSIZE[121] = AP_AXIMM_121_ARSIZE;
            assign ap_ARBURST[121] = AP_AXIMM_121_ARBURST;
            assign ap_ARLOCK[121] = AP_AXIMM_121_ARLOCK;
            assign ap_ARCACHE[121] = AP_AXIMM_121_ARCACHE;
            assign ap_ARPROT[121] = AP_AXIMM_121_ARPROT;
            assign ap_ARREGION[121] = AP_AXIMM_121_ARREGION;
            assign ap_ARQOS[121] = AP_AXIMM_121_ARQOS;
            assign ap_ARVALID[121] = AP_AXIMM_121_ARVALID;
            assign AP_AXIMM_121_ARREADY = ap_ARREADY[121];
            assign AP_AXIMM_121_RDATA = ap_RDATA[121][M_AXIMM_121_DATA_WIDTH-1:0];
            assign AP_AXIMM_121_RRESP = ap_RRESP[121];
            assign AP_AXIMM_121_RLAST = ap_RLAST[121];
            assign AP_AXIMM_121_RVALID = ap_RVALID[121];
            assign ap_RREADY[121] = AP_AXIMM_121_RREADY;
            assign M_AXIMM_121_AWADDR = dm_AWADDR[121][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_121_AWLEN = dm_AWLEN[121];
            assign M_AXIMM_121_AWSIZE = dm_AWSIZE[121];
            assign M_AXIMM_121_AWBURST = dm_AWBURST[121];
            assign M_AXIMM_121_AWLOCK = dm_AWLOCK[121];
            assign M_AXIMM_121_AWCACHE = dm_AWCACHE[121];
            assign M_AXIMM_121_AWPROT = dm_AWPROT[121];
            assign M_AXIMM_121_AWREGION = dm_AWREGION[121];
            assign M_AXIMM_121_AWQOS = dm_AWQOS[121];
            assign M_AXIMM_121_AWVALID = dm_AWVALID[121];
            assign dm_AWREADY[121] = M_AXIMM_121_AWREADY;
            assign M_AXIMM_121_WDATA = dm_WDATA[121][M_AXIMM_121_DATA_WIDTH-1:0];
            assign M_AXIMM_121_WSTRB = dm_WSTRB[121][M_AXIMM_121_DATA_WIDTH/8-1:0];
            assign M_AXIMM_121_WLAST = dm_WLAST[121];
            assign M_AXIMM_121_WVALID = dm_WVALID[121];
            assign dm_WREADY[121] = M_AXIMM_121_WREADY;
            assign dm_BRESP[121] = M_AXIMM_121_BRESP;
            assign dm_BVALID[121] = M_AXIMM_121_BVALID;
            assign M_AXIMM_121_BREADY = dm_BREADY[121];
            assign M_AXIMM_121_ARADDR = dm_ARADDR[121][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_121_ARLEN = dm_ARLEN[121];
            assign M_AXIMM_121_ARSIZE = dm_ARSIZE[121];
            assign M_AXIMM_121_ARBURST = dm_ARBURST[121];
            assign M_AXIMM_121_ARLOCK = dm_ARLOCK[121];
            assign M_AXIMM_121_ARCACHE = dm_ARCACHE[121];
            assign M_AXIMM_121_ARPROT = dm_ARPROT[121];
            assign M_AXIMM_121_ARREGION = dm_ARREGION[121];
            assign M_AXIMM_121_ARQOS = dm_ARQOS[121];
            assign M_AXIMM_121_ARVALID = dm_ARVALID[121];
            assign dm_ARREADY[121] = M_AXIMM_121_ARREADY;
            assign dm_RDATA[121][M_AXIMM_121_DATA_WIDTH-1:0] = M_AXIMM_121_RDATA;
            assign dm_RRESP[121] = M_AXIMM_121_RRESP;
            assign dm_RLAST[121] = M_AXIMM_121_RLAST;
            assign dm_RVALID[121] = M_AXIMM_121_RVALID;
            assign M_AXIMM_121_RREADY = dm_RREADY[121];
        end
        if(C_NUM_AXIMMs > 122) begin
            assign ap_AWADDR[122][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_122_AWADDR;
            assign ap_AWLEN[122] = AP_AXIMM_122_AWLEN;
            assign ap_AWSIZE[122] = AP_AXIMM_122_AWSIZE;
            assign ap_AWBURST[122] = AP_AXIMM_122_AWBURST;
            assign ap_AWLOCK[122] = AP_AXIMM_122_AWLOCK;
            assign ap_AWCACHE[122] = AP_AXIMM_122_AWCACHE;
            assign ap_AWPROT[122] = AP_AXIMM_122_AWPROT;
            assign ap_AWREGION[122] = AP_AXIMM_122_AWREGION;
            assign ap_AWQOS[122] = AP_AXIMM_122_AWQOS;
            assign ap_AWVALID[122] = AP_AXIMM_122_AWVALID;
            assign AP_AXIMM_122_AWREADY = ap_AWREADY[122];
            assign ap_WDATA[122][M_AXIMM_122_DATA_WIDTH-1:0] = AP_AXIMM_122_WDATA;
            assign ap_WSTRB[122][M_AXIMM_122_DATA_WIDTH/8-1:0] = AP_AXIMM_122_WSTRB;
            assign ap_WLAST[122] = AP_AXIMM_122_WLAST;
            assign ap_WVALID[122] = AP_AXIMM_122_WVALID;
            assign AP_AXIMM_122_WREADY = ap_WREADY[122];
            assign AP_AXIMM_122_BRESP = ap_BRESP[122];
            assign AP_AXIMM_122_BVALID = ap_BVALID[122];
            assign ap_BREADY[122] = AP_AXIMM_122_BREADY;
            assign ap_ARADDR[122][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_122_ARADDR;
            assign ap_ARLEN[122] = AP_AXIMM_122_ARLEN;
            assign ap_ARSIZE[122] = AP_AXIMM_122_ARSIZE;
            assign ap_ARBURST[122] = AP_AXIMM_122_ARBURST;
            assign ap_ARLOCK[122] = AP_AXIMM_122_ARLOCK;
            assign ap_ARCACHE[122] = AP_AXIMM_122_ARCACHE;
            assign ap_ARPROT[122] = AP_AXIMM_122_ARPROT;
            assign ap_ARREGION[122] = AP_AXIMM_122_ARREGION;
            assign ap_ARQOS[122] = AP_AXIMM_122_ARQOS;
            assign ap_ARVALID[122] = AP_AXIMM_122_ARVALID;
            assign AP_AXIMM_122_ARREADY = ap_ARREADY[122];
            assign AP_AXIMM_122_RDATA = ap_RDATA[122][M_AXIMM_122_DATA_WIDTH-1:0];
            assign AP_AXIMM_122_RRESP = ap_RRESP[122];
            assign AP_AXIMM_122_RLAST = ap_RLAST[122];
            assign AP_AXIMM_122_RVALID = ap_RVALID[122];
            assign ap_RREADY[122] = AP_AXIMM_122_RREADY;
            assign M_AXIMM_122_AWADDR = dm_AWADDR[122][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_122_AWLEN = dm_AWLEN[122];
            assign M_AXIMM_122_AWSIZE = dm_AWSIZE[122];
            assign M_AXIMM_122_AWBURST = dm_AWBURST[122];
            assign M_AXIMM_122_AWLOCK = dm_AWLOCK[122];
            assign M_AXIMM_122_AWCACHE = dm_AWCACHE[122];
            assign M_AXIMM_122_AWPROT = dm_AWPROT[122];
            assign M_AXIMM_122_AWREGION = dm_AWREGION[122];
            assign M_AXIMM_122_AWQOS = dm_AWQOS[122];
            assign M_AXIMM_122_AWVALID = dm_AWVALID[122];
            assign dm_AWREADY[122] = M_AXIMM_122_AWREADY;
            assign M_AXIMM_122_WDATA = dm_WDATA[122][M_AXIMM_122_DATA_WIDTH-1:0];
            assign M_AXIMM_122_WSTRB = dm_WSTRB[122][M_AXIMM_122_DATA_WIDTH/8-1:0];
            assign M_AXIMM_122_WLAST = dm_WLAST[122];
            assign M_AXIMM_122_WVALID = dm_WVALID[122];
            assign dm_WREADY[122] = M_AXIMM_122_WREADY;
            assign dm_BRESP[122] = M_AXIMM_122_BRESP;
            assign dm_BVALID[122] = M_AXIMM_122_BVALID;
            assign M_AXIMM_122_BREADY = dm_BREADY[122];
            assign M_AXIMM_122_ARADDR = dm_ARADDR[122][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_122_ARLEN = dm_ARLEN[122];
            assign M_AXIMM_122_ARSIZE = dm_ARSIZE[122];
            assign M_AXIMM_122_ARBURST = dm_ARBURST[122];
            assign M_AXIMM_122_ARLOCK = dm_ARLOCK[122];
            assign M_AXIMM_122_ARCACHE = dm_ARCACHE[122];
            assign M_AXIMM_122_ARPROT = dm_ARPROT[122];
            assign M_AXIMM_122_ARREGION = dm_ARREGION[122];
            assign M_AXIMM_122_ARQOS = dm_ARQOS[122];
            assign M_AXIMM_122_ARVALID = dm_ARVALID[122];
            assign dm_ARREADY[122] = M_AXIMM_122_ARREADY;
            assign dm_RDATA[122][M_AXIMM_122_DATA_WIDTH-1:0] = M_AXIMM_122_RDATA;
            assign dm_RRESP[122] = M_AXIMM_122_RRESP;
            assign dm_RLAST[122] = M_AXIMM_122_RLAST;
            assign dm_RVALID[122] = M_AXIMM_122_RVALID;
            assign M_AXIMM_122_RREADY = dm_RREADY[122];
        end
        if(C_NUM_AXIMMs > 123) begin
            assign ap_AWADDR[123][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_123_AWADDR;
            assign ap_AWLEN[123] = AP_AXIMM_123_AWLEN;
            assign ap_AWSIZE[123] = AP_AXIMM_123_AWSIZE;
            assign ap_AWBURST[123] = AP_AXIMM_123_AWBURST;
            assign ap_AWLOCK[123] = AP_AXIMM_123_AWLOCK;
            assign ap_AWCACHE[123] = AP_AXIMM_123_AWCACHE;
            assign ap_AWPROT[123] = AP_AXIMM_123_AWPROT;
            assign ap_AWREGION[123] = AP_AXIMM_123_AWREGION;
            assign ap_AWQOS[123] = AP_AXIMM_123_AWQOS;
            assign ap_AWVALID[123] = AP_AXIMM_123_AWVALID;
            assign AP_AXIMM_123_AWREADY = ap_AWREADY[123];
            assign ap_WDATA[123][M_AXIMM_123_DATA_WIDTH-1:0] = AP_AXIMM_123_WDATA;
            assign ap_WSTRB[123][M_AXIMM_123_DATA_WIDTH/8-1:0] = AP_AXIMM_123_WSTRB;
            assign ap_WLAST[123] = AP_AXIMM_123_WLAST;
            assign ap_WVALID[123] = AP_AXIMM_123_WVALID;
            assign AP_AXIMM_123_WREADY = ap_WREADY[123];
            assign AP_AXIMM_123_BRESP = ap_BRESP[123];
            assign AP_AXIMM_123_BVALID = ap_BVALID[123];
            assign ap_BREADY[123] = AP_AXIMM_123_BREADY;
            assign ap_ARADDR[123][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_123_ARADDR;
            assign ap_ARLEN[123] = AP_AXIMM_123_ARLEN;
            assign ap_ARSIZE[123] = AP_AXIMM_123_ARSIZE;
            assign ap_ARBURST[123] = AP_AXIMM_123_ARBURST;
            assign ap_ARLOCK[123] = AP_AXIMM_123_ARLOCK;
            assign ap_ARCACHE[123] = AP_AXIMM_123_ARCACHE;
            assign ap_ARPROT[123] = AP_AXIMM_123_ARPROT;
            assign ap_ARREGION[123] = AP_AXIMM_123_ARREGION;
            assign ap_ARQOS[123] = AP_AXIMM_123_ARQOS;
            assign ap_ARVALID[123] = AP_AXIMM_123_ARVALID;
            assign AP_AXIMM_123_ARREADY = ap_ARREADY[123];
            assign AP_AXIMM_123_RDATA = ap_RDATA[123][M_AXIMM_123_DATA_WIDTH-1:0];
            assign AP_AXIMM_123_RRESP = ap_RRESP[123];
            assign AP_AXIMM_123_RLAST = ap_RLAST[123];
            assign AP_AXIMM_123_RVALID = ap_RVALID[123];
            assign ap_RREADY[123] = AP_AXIMM_123_RREADY;
            assign M_AXIMM_123_AWADDR = dm_AWADDR[123][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_123_AWLEN = dm_AWLEN[123];
            assign M_AXIMM_123_AWSIZE = dm_AWSIZE[123];
            assign M_AXIMM_123_AWBURST = dm_AWBURST[123];
            assign M_AXIMM_123_AWLOCK = dm_AWLOCK[123];
            assign M_AXIMM_123_AWCACHE = dm_AWCACHE[123];
            assign M_AXIMM_123_AWPROT = dm_AWPROT[123];
            assign M_AXIMM_123_AWREGION = dm_AWREGION[123];
            assign M_AXIMM_123_AWQOS = dm_AWQOS[123];
            assign M_AXIMM_123_AWVALID = dm_AWVALID[123];
            assign dm_AWREADY[123] = M_AXIMM_123_AWREADY;
            assign M_AXIMM_123_WDATA = dm_WDATA[123][M_AXIMM_123_DATA_WIDTH-1:0];
            assign M_AXIMM_123_WSTRB = dm_WSTRB[123][M_AXIMM_123_DATA_WIDTH/8-1:0];
            assign M_AXIMM_123_WLAST = dm_WLAST[123];
            assign M_AXIMM_123_WVALID = dm_WVALID[123];
            assign dm_WREADY[123] = M_AXIMM_123_WREADY;
            assign dm_BRESP[123] = M_AXIMM_123_BRESP;
            assign dm_BVALID[123] = M_AXIMM_123_BVALID;
            assign M_AXIMM_123_BREADY = dm_BREADY[123];
            assign M_AXIMM_123_ARADDR = dm_ARADDR[123][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_123_ARLEN = dm_ARLEN[123];
            assign M_AXIMM_123_ARSIZE = dm_ARSIZE[123];
            assign M_AXIMM_123_ARBURST = dm_ARBURST[123];
            assign M_AXIMM_123_ARLOCK = dm_ARLOCK[123];
            assign M_AXIMM_123_ARCACHE = dm_ARCACHE[123];
            assign M_AXIMM_123_ARPROT = dm_ARPROT[123];
            assign M_AXIMM_123_ARREGION = dm_ARREGION[123];
            assign M_AXIMM_123_ARQOS = dm_ARQOS[123];
            assign M_AXIMM_123_ARVALID = dm_ARVALID[123];
            assign dm_ARREADY[123] = M_AXIMM_123_ARREADY;
            assign dm_RDATA[123][M_AXIMM_123_DATA_WIDTH-1:0] = M_AXIMM_123_RDATA;
            assign dm_RRESP[123] = M_AXIMM_123_RRESP;
            assign dm_RLAST[123] = M_AXIMM_123_RLAST;
            assign dm_RVALID[123] = M_AXIMM_123_RVALID;
            assign M_AXIMM_123_RREADY = dm_RREADY[123];
        end
        if(C_NUM_AXIMMs > 124) begin
            assign ap_AWADDR[124][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_124_AWADDR;
            assign ap_AWLEN[124] = AP_AXIMM_124_AWLEN;
            assign ap_AWSIZE[124] = AP_AXIMM_124_AWSIZE;
            assign ap_AWBURST[124] = AP_AXIMM_124_AWBURST;
            assign ap_AWLOCK[124] = AP_AXIMM_124_AWLOCK;
            assign ap_AWCACHE[124] = AP_AXIMM_124_AWCACHE;
            assign ap_AWPROT[124] = AP_AXIMM_124_AWPROT;
            assign ap_AWREGION[124] = AP_AXIMM_124_AWREGION;
            assign ap_AWQOS[124] = AP_AXIMM_124_AWQOS;
            assign ap_AWVALID[124] = AP_AXIMM_124_AWVALID;
            assign AP_AXIMM_124_AWREADY = ap_AWREADY[124];
            assign ap_WDATA[124][M_AXIMM_124_DATA_WIDTH-1:0] = AP_AXIMM_124_WDATA;
            assign ap_WSTRB[124][M_AXIMM_124_DATA_WIDTH/8-1:0] = AP_AXIMM_124_WSTRB;
            assign ap_WLAST[124] = AP_AXIMM_124_WLAST;
            assign ap_WVALID[124] = AP_AXIMM_124_WVALID;
            assign AP_AXIMM_124_WREADY = ap_WREADY[124];
            assign AP_AXIMM_124_BRESP = ap_BRESP[124];
            assign AP_AXIMM_124_BVALID = ap_BVALID[124];
            assign ap_BREADY[124] = AP_AXIMM_124_BREADY;
            assign ap_ARADDR[124][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_124_ARADDR;
            assign ap_ARLEN[124] = AP_AXIMM_124_ARLEN;
            assign ap_ARSIZE[124] = AP_AXIMM_124_ARSIZE;
            assign ap_ARBURST[124] = AP_AXIMM_124_ARBURST;
            assign ap_ARLOCK[124] = AP_AXIMM_124_ARLOCK;
            assign ap_ARCACHE[124] = AP_AXIMM_124_ARCACHE;
            assign ap_ARPROT[124] = AP_AXIMM_124_ARPROT;
            assign ap_ARREGION[124] = AP_AXIMM_124_ARREGION;
            assign ap_ARQOS[124] = AP_AXIMM_124_ARQOS;
            assign ap_ARVALID[124] = AP_AXIMM_124_ARVALID;
            assign AP_AXIMM_124_ARREADY = ap_ARREADY[124];
            assign AP_AXIMM_124_RDATA = ap_RDATA[124][M_AXIMM_124_DATA_WIDTH-1:0];
            assign AP_AXIMM_124_RRESP = ap_RRESP[124];
            assign AP_AXIMM_124_RLAST = ap_RLAST[124];
            assign AP_AXIMM_124_RVALID = ap_RVALID[124];
            assign ap_RREADY[124] = AP_AXIMM_124_RREADY;
            assign M_AXIMM_124_AWADDR = dm_AWADDR[124][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_124_AWLEN = dm_AWLEN[124];
            assign M_AXIMM_124_AWSIZE = dm_AWSIZE[124];
            assign M_AXIMM_124_AWBURST = dm_AWBURST[124];
            assign M_AXIMM_124_AWLOCK = dm_AWLOCK[124];
            assign M_AXIMM_124_AWCACHE = dm_AWCACHE[124];
            assign M_AXIMM_124_AWPROT = dm_AWPROT[124];
            assign M_AXIMM_124_AWREGION = dm_AWREGION[124];
            assign M_AXIMM_124_AWQOS = dm_AWQOS[124];
            assign M_AXIMM_124_AWVALID = dm_AWVALID[124];
            assign dm_AWREADY[124] = M_AXIMM_124_AWREADY;
            assign M_AXIMM_124_WDATA = dm_WDATA[124][M_AXIMM_124_DATA_WIDTH-1:0];
            assign M_AXIMM_124_WSTRB = dm_WSTRB[124][M_AXIMM_124_DATA_WIDTH/8-1:0];
            assign M_AXIMM_124_WLAST = dm_WLAST[124];
            assign M_AXIMM_124_WVALID = dm_WVALID[124];
            assign dm_WREADY[124] = M_AXIMM_124_WREADY;
            assign dm_BRESP[124] = M_AXIMM_124_BRESP;
            assign dm_BVALID[124] = M_AXIMM_124_BVALID;
            assign M_AXIMM_124_BREADY = dm_BREADY[124];
            assign M_AXIMM_124_ARADDR = dm_ARADDR[124][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_124_ARLEN = dm_ARLEN[124];
            assign M_AXIMM_124_ARSIZE = dm_ARSIZE[124];
            assign M_AXIMM_124_ARBURST = dm_ARBURST[124];
            assign M_AXIMM_124_ARLOCK = dm_ARLOCK[124];
            assign M_AXIMM_124_ARCACHE = dm_ARCACHE[124];
            assign M_AXIMM_124_ARPROT = dm_ARPROT[124];
            assign M_AXIMM_124_ARREGION = dm_ARREGION[124];
            assign M_AXIMM_124_ARQOS = dm_ARQOS[124];
            assign M_AXIMM_124_ARVALID = dm_ARVALID[124];
            assign dm_ARREADY[124] = M_AXIMM_124_ARREADY;
            assign dm_RDATA[124][M_AXIMM_124_DATA_WIDTH-1:0] = M_AXIMM_124_RDATA;
            assign dm_RRESP[124] = M_AXIMM_124_RRESP;
            assign dm_RLAST[124] = M_AXIMM_124_RLAST;
            assign dm_RVALID[124] = M_AXIMM_124_RVALID;
            assign M_AXIMM_124_RREADY = dm_RREADY[124];
        end
        if(C_NUM_AXIMMs > 125) begin
            assign ap_AWADDR[125][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_125_AWADDR;
            assign ap_AWLEN[125] = AP_AXIMM_125_AWLEN;
            assign ap_AWSIZE[125] = AP_AXIMM_125_AWSIZE;
            assign ap_AWBURST[125] = AP_AXIMM_125_AWBURST;
            assign ap_AWLOCK[125] = AP_AXIMM_125_AWLOCK;
            assign ap_AWCACHE[125] = AP_AXIMM_125_AWCACHE;
            assign ap_AWPROT[125] = AP_AXIMM_125_AWPROT;
            assign ap_AWREGION[125] = AP_AXIMM_125_AWREGION;
            assign ap_AWQOS[125] = AP_AXIMM_125_AWQOS;
            assign ap_AWVALID[125] = AP_AXIMM_125_AWVALID;
            assign AP_AXIMM_125_AWREADY = ap_AWREADY[125];
            assign ap_WDATA[125][M_AXIMM_125_DATA_WIDTH-1:0] = AP_AXIMM_125_WDATA;
            assign ap_WSTRB[125][M_AXIMM_125_DATA_WIDTH/8-1:0] = AP_AXIMM_125_WSTRB;
            assign ap_WLAST[125] = AP_AXIMM_125_WLAST;
            assign ap_WVALID[125] = AP_AXIMM_125_WVALID;
            assign AP_AXIMM_125_WREADY = ap_WREADY[125];
            assign AP_AXIMM_125_BRESP = ap_BRESP[125];
            assign AP_AXIMM_125_BVALID = ap_BVALID[125];
            assign ap_BREADY[125] = AP_AXIMM_125_BREADY;
            assign ap_ARADDR[125][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_125_ARADDR;
            assign ap_ARLEN[125] = AP_AXIMM_125_ARLEN;
            assign ap_ARSIZE[125] = AP_AXIMM_125_ARSIZE;
            assign ap_ARBURST[125] = AP_AXIMM_125_ARBURST;
            assign ap_ARLOCK[125] = AP_AXIMM_125_ARLOCK;
            assign ap_ARCACHE[125] = AP_AXIMM_125_ARCACHE;
            assign ap_ARPROT[125] = AP_AXIMM_125_ARPROT;
            assign ap_ARREGION[125] = AP_AXIMM_125_ARREGION;
            assign ap_ARQOS[125] = AP_AXIMM_125_ARQOS;
            assign ap_ARVALID[125] = AP_AXIMM_125_ARVALID;
            assign AP_AXIMM_125_ARREADY = ap_ARREADY[125];
            assign AP_AXIMM_125_RDATA = ap_RDATA[125][M_AXIMM_125_DATA_WIDTH-1:0];
            assign AP_AXIMM_125_RRESP = ap_RRESP[125];
            assign AP_AXIMM_125_RLAST = ap_RLAST[125];
            assign AP_AXIMM_125_RVALID = ap_RVALID[125];
            assign ap_RREADY[125] = AP_AXIMM_125_RREADY;
            assign M_AXIMM_125_AWADDR = dm_AWADDR[125][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_125_AWLEN = dm_AWLEN[125];
            assign M_AXIMM_125_AWSIZE = dm_AWSIZE[125];
            assign M_AXIMM_125_AWBURST = dm_AWBURST[125];
            assign M_AXIMM_125_AWLOCK = dm_AWLOCK[125];
            assign M_AXIMM_125_AWCACHE = dm_AWCACHE[125];
            assign M_AXIMM_125_AWPROT = dm_AWPROT[125];
            assign M_AXIMM_125_AWREGION = dm_AWREGION[125];
            assign M_AXIMM_125_AWQOS = dm_AWQOS[125];
            assign M_AXIMM_125_AWVALID = dm_AWVALID[125];
            assign dm_AWREADY[125] = M_AXIMM_125_AWREADY;
            assign M_AXIMM_125_WDATA = dm_WDATA[125][M_AXIMM_125_DATA_WIDTH-1:0];
            assign M_AXIMM_125_WSTRB = dm_WSTRB[125][M_AXIMM_125_DATA_WIDTH/8-1:0];
            assign M_AXIMM_125_WLAST = dm_WLAST[125];
            assign M_AXIMM_125_WVALID = dm_WVALID[125];
            assign dm_WREADY[125] = M_AXIMM_125_WREADY;
            assign dm_BRESP[125] = M_AXIMM_125_BRESP;
            assign dm_BVALID[125] = M_AXIMM_125_BVALID;
            assign M_AXIMM_125_BREADY = dm_BREADY[125];
            assign M_AXIMM_125_ARADDR = dm_ARADDR[125][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_125_ARLEN = dm_ARLEN[125];
            assign M_AXIMM_125_ARSIZE = dm_ARSIZE[125];
            assign M_AXIMM_125_ARBURST = dm_ARBURST[125];
            assign M_AXIMM_125_ARLOCK = dm_ARLOCK[125];
            assign M_AXIMM_125_ARCACHE = dm_ARCACHE[125];
            assign M_AXIMM_125_ARPROT = dm_ARPROT[125];
            assign M_AXIMM_125_ARREGION = dm_ARREGION[125];
            assign M_AXIMM_125_ARQOS = dm_ARQOS[125];
            assign M_AXIMM_125_ARVALID = dm_ARVALID[125];
            assign dm_ARREADY[125] = M_AXIMM_125_ARREADY;
            assign dm_RDATA[125][M_AXIMM_125_DATA_WIDTH-1:0] = M_AXIMM_125_RDATA;
            assign dm_RRESP[125] = M_AXIMM_125_RRESP;
            assign dm_RLAST[125] = M_AXIMM_125_RLAST;
            assign dm_RVALID[125] = M_AXIMM_125_RVALID;
            assign M_AXIMM_125_RREADY = dm_RREADY[125];
        end
        if(C_NUM_AXIMMs > 126) begin
            assign ap_AWADDR[126][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_126_AWADDR;
            assign ap_AWLEN[126] = AP_AXIMM_126_AWLEN;
            assign ap_AWSIZE[126] = AP_AXIMM_126_AWSIZE;
            assign ap_AWBURST[126] = AP_AXIMM_126_AWBURST;
            assign ap_AWLOCK[126] = AP_AXIMM_126_AWLOCK;
            assign ap_AWCACHE[126] = AP_AXIMM_126_AWCACHE;
            assign ap_AWPROT[126] = AP_AXIMM_126_AWPROT;
            assign ap_AWREGION[126] = AP_AXIMM_126_AWREGION;
            assign ap_AWQOS[126] = AP_AXIMM_126_AWQOS;
            assign ap_AWVALID[126] = AP_AXIMM_126_AWVALID;
            assign AP_AXIMM_126_AWREADY = ap_AWREADY[126];
            assign ap_WDATA[126][M_AXIMM_126_DATA_WIDTH-1:0] = AP_AXIMM_126_WDATA;
            assign ap_WSTRB[126][M_AXIMM_126_DATA_WIDTH/8-1:0] = AP_AXIMM_126_WSTRB;
            assign ap_WLAST[126] = AP_AXIMM_126_WLAST;
            assign ap_WVALID[126] = AP_AXIMM_126_WVALID;
            assign AP_AXIMM_126_WREADY = ap_WREADY[126];
            assign AP_AXIMM_126_BRESP = ap_BRESP[126];
            assign AP_AXIMM_126_BVALID = ap_BVALID[126];
            assign ap_BREADY[126] = AP_AXIMM_126_BREADY;
            assign ap_ARADDR[126][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_126_ARADDR;
            assign ap_ARLEN[126] = AP_AXIMM_126_ARLEN;
            assign ap_ARSIZE[126] = AP_AXIMM_126_ARSIZE;
            assign ap_ARBURST[126] = AP_AXIMM_126_ARBURST;
            assign ap_ARLOCK[126] = AP_AXIMM_126_ARLOCK;
            assign ap_ARCACHE[126] = AP_AXIMM_126_ARCACHE;
            assign ap_ARPROT[126] = AP_AXIMM_126_ARPROT;
            assign ap_ARREGION[126] = AP_AXIMM_126_ARREGION;
            assign ap_ARQOS[126] = AP_AXIMM_126_ARQOS;
            assign ap_ARVALID[126] = AP_AXIMM_126_ARVALID;
            assign AP_AXIMM_126_ARREADY = ap_ARREADY[126];
            assign AP_AXIMM_126_RDATA = ap_RDATA[126][M_AXIMM_126_DATA_WIDTH-1:0];
            assign AP_AXIMM_126_RRESP = ap_RRESP[126];
            assign AP_AXIMM_126_RLAST = ap_RLAST[126];
            assign AP_AXIMM_126_RVALID = ap_RVALID[126];
            assign ap_RREADY[126] = AP_AXIMM_126_RREADY;
            assign M_AXIMM_126_AWADDR = dm_AWADDR[126][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_126_AWLEN = dm_AWLEN[126];
            assign M_AXIMM_126_AWSIZE = dm_AWSIZE[126];
            assign M_AXIMM_126_AWBURST = dm_AWBURST[126];
            assign M_AXIMM_126_AWLOCK = dm_AWLOCK[126];
            assign M_AXIMM_126_AWCACHE = dm_AWCACHE[126];
            assign M_AXIMM_126_AWPROT = dm_AWPROT[126];
            assign M_AXIMM_126_AWREGION = dm_AWREGION[126];
            assign M_AXIMM_126_AWQOS = dm_AWQOS[126];
            assign M_AXIMM_126_AWVALID = dm_AWVALID[126];
            assign dm_AWREADY[126] = M_AXIMM_126_AWREADY;
            assign M_AXIMM_126_WDATA = dm_WDATA[126][M_AXIMM_126_DATA_WIDTH-1:0];
            assign M_AXIMM_126_WSTRB = dm_WSTRB[126][M_AXIMM_126_DATA_WIDTH/8-1:0];
            assign M_AXIMM_126_WLAST = dm_WLAST[126];
            assign M_AXIMM_126_WVALID = dm_WVALID[126];
            assign dm_WREADY[126] = M_AXIMM_126_WREADY;
            assign dm_BRESP[126] = M_AXIMM_126_BRESP;
            assign dm_BVALID[126] = M_AXIMM_126_BVALID;
            assign M_AXIMM_126_BREADY = dm_BREADY[126];
            assign M_AXIMM_126_ARADDR = dm_ARADDR[126][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_126_ARLEN = dm_ARLEN[126];
            assign M_AXIMM_126_ARSIZE = dm_ARSIZE[126];
            assign M_AXIMM_126_ARBURST = dm_ARBURST[126];
            assign M_AXIMM_126_ARLOCK = dm_ARLOCK[126];
            assign M_AXIMM_126_ARCACHE = dm_ARCACHE[126];
            assign M_AXIMM_126_ARPROT = dm_ARPROT[126];
            assign M_AXIMM_126_ARREGION = dm_ARREGION[126];
            assign M_AXIMM_126_ARQOS = dm_ARQOS[126];
            assign M_AXIMM_126_ARVALID = dm_ARVALID[126];
            assign dm_ARREADY[126] = M_AXIMM_126_ARREADY;
            assign dm_RDATA[126][M_AXIMM_126_DATA_WIDTH-1:0] = M_AXIMM_126_RDATA;
            assign dm_RRESP[126] = M_AXIMM_126_RRESP;
            assign dm_RLAST[126] = M_AXIMM_126_RLAST;
            assign dm_RVALID[126] = M_AXIMM_126_RVALID;
            assign M_AXIMM_126_RREADY = dm_RREADY[126];
        end
        if(C_NUM_AXIMMs > 127) begin
            assign ap_AWADDR[127][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_127_AWADDR;
            assign ap_AWLEN[127] = AP_AXIMM_127_AWLEN;
            assign ap_AWSIZE[127] = AP_AXIMM_127_AWSIZE;
            assign ap_AWBURST[127] = AP_AXIMM_127_AWBURST;
            assign ap_AWLOCK[127] = AP_AXIMM_127_AWLOCK;
            assign ap_AWCACHE[127] = AP_AXIMM_127_AWCACHE;
            assign ap_AWPROT[127] = AP_AXIMM_127_AWPROT;
            assign ap_AWREGION[127] = AP_AXIMM_127_AWREGION;
            assign ap_AWQOS[127] = AP_AXIMM_127_AWQOS;
            assign ap_AWVALID[127] = AP_AXIMM_127_AWVALID;
            assign AP_AXIMM_127_AWREADY = ap_AWREADY[127];
            assign ap_WDATA[127][M_AXIMM_127_DATA_WIDTH-1:0] = AP_AXIMM_127_WDATA;
            assign ap_WSTRB[127][M_AXIMM_127_DATA_WIDTH/8-1:0] = AP_AXIMM_127_WSTRB;
            assign ap_WLAST[127] = AP_AXIMM_127_WLAST;
            assign ap_WVALID[127] = AP_AXIMM_127_WVALID;
            assign AP_AXIMM_127_WREADY = ap_WREADY[127];
            assign AP_AXIMM_127_BRESP = ap_BRESP[127];
            assign AP_AXIMM_127_BVALID = ap_BVALID[127];
            assign ap_BREADY[127] = AP_AXIMM_127_BREADY;
            assign ap_ARADDR[127][M_AXIMM_ADDR_WIDTH-1:0] = AP_AXIMM_127_ARADDR;
            assign ap_ARLEN[127] = AP_AXIMM_127_ARLEN;
            assign ap_ARSIZE[127] = AP_AXIMM_127_ARSIZE;
            assign ap_ARBURST[127] = AP_AXIMM_127_ARBURST;
            assign ap_ARLOCK[127] = AP_AXIMM_127_ARLOCK;
            assign ap_ARCACHE[127] = AP_AXIMM_127_ARCACHE;
            assign ap_ARPROT[127] = AP_AXIMM_127_ARPROT;
            assign ap_ARREGION[127] = AP_AXIMM_127_ARREGION;
            assign ap_ARQOS[127] = AP_AXIMM_127_ARQOS;
            assign ap_ARVALID[127] = AP_AXIMM_127_ARVALID;
            assign AP_AXIMM_127_ARREADY = ap_ARREADY[127];
            assign AP_AXIMM_127_RDATA = ap_RDATA[127][M_AXIMM_127_DATA_WIDTH-1:0];
            assign AP_AXIMM_127_RRESP = ap_RRESP[127];
            assign AP_AXIMM_127_RLAST = ap_RLAST[127];
            assign AP_AXIMM_127_RVALID = ap_RVALID[127];
            assign ap_RREADY[127] = AP_AXIMM_127_RREADY;
            assign M_AXIMM_127_AWADDR = dm_AWADDR[127][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_127_AWLEN = dm_AWLEN[127];
            assign M_AXIMM_127_AWSIZE = dm_AWSIZE[127];
            assign M_AXIMM_127_AWBURST = dm_AWBURST[127];
            assign M_AXIMM_127_AWLOCK = dm_AWLOCK[127];
            assign M_AXIMM_127_AWCACHE = dm_AWCACHE[127];
            assign M_AXIMM_127_AWPROT = dm_AWPROT[127];
            assign M_AXIMM_127_AWREGION = dm_AWREGION[127];
            assign M_AXIMM_127_AWQOS = dm_AWQOS[127];
            assign M_AXIMM_127_AWVALID = dm_AWVALID[127];
            assign dm_AWREADY[127] = M_AXIMM_127_AWREADY;
            assign M_AXIMM_127_WDATA = dm_WDATA[127][M_AXIMM_127_DATA_WIDTH-1:0];
            assign M_AXIMM_127_WSTRB = dm_WSTRB[127][M_AXIMM_127_DATA_WIDTH/8-1:0];
            assign M_AXIMM_127_WLAST = dm_WLAST[127];
            assign M_AXIMM_127_WVALID = dm_WVALID[127];
            assign dm_WREADY[127] = M_AXIMM_127_WREADY;
            assign dm_BRESP[127] = M_AXIMM_127_BRESP;
            assign dm_BVALID[127] = M_AXIMM_127_BVALID;
            assign M_AXIMM_127_BREADY = dm_BREADY[127];
            assign M_AXIMM_127_ARADDR = dm_ARADDR[127][M_AXIMM_ADDR_WIDTH-1:0];
            assign M_AXIMM_127_ARLEN = dm_ARLEN[127];
            assign M_AXIMM_127_ARSIZE = dm_ARSIZE[127];
            assign M_AXIMM_127_ARBURST = dm_ARBURST[127];
            assign M_AXIMM_127_ARLOCK = dm_ARLOCK[127];
            assign M_AXIMM_127_ARCACHE = dm_ARCACHE[127];
            assign M_AXIMM_127_ARPROT = dm_ARPROT[127];
            assign M_AXIMM_127_ARREGION = dm_ARREGION[127];
            assign M_AXIMM_127_ARQOS = dm_ARQOS[127];
            assign M_AXIMM_127_ARVALID = dm_ARVALID[127];
            assign dm_ARREADY[127] = M_AXIMM_127_ARREADY;
            assign dm_RDATA[127][M_AXIMM_127_DATA_WIDTH-1:0] = M_AXIMM_127_RDATA;
            assign dm_RRESP[127] = M_AXIMM_127_RRESP;
            assign dm_RLAST[127] = M_AXIMM_127_RLAST;
            assign dm_RVALID[127] = M_AXIMM_127_RVALID;
            assign M_AXIMM_127_RREADY = dm_RREADY[127];
        end
    endgenerate    
    
    //wire up
    genvar idx;
    generate
        for(idx=0; idx<C_NUM_AXIMMs; idx=idx+1) begin: AXIMM_GEN
            //just wire signals straight through
            assign dm_AWADDR[idx][M_AXIMM_ADDR_WIDTH-1:0] = ap_AWADDR[idx][M_AXIMM_ADDR_WIDTH-1:0];
            assign dm_AWLEN[idx] = ap_AWLEN[idx];
            assign dm_AWSIZE[idx] = ap_AWSIZE[idx];
            assign dm_AWBURST[idx] = ap_AWBURST[idx];
            assign dm_AWLOCK[idx] = ap_AWLOCK[idx];
            assign dm_AWCACHE[idx] = ap_AWCACHE[idx];
            assign dm_AWPROT[idx] = ap_AWPROT[idx];
            assign dm_AWREGION[idx] = ap_AWREGION[idx];
            assign dm_AWQOS[idx] = ap_AWQOS[idx];
            assign dm_AWVALID[idx] = ap_AWVALID[idx];
            assign ap_AWREADY[idx] = dm_AWREADY[idx];
            assign dm_WDATA[idx][M_AXIMM_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = ap_WDATA[idx][M_AXIMM_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            assign dm_WSTRB[idx][M_AXIMM_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0] = ap_WSTRB[idx][M_AXIMM_BIT_ARRAY[32*(idx+1)-1:32*idx]/8-1:0];
            assign dm_WLAST[idx] = ap_WLAST[idx];
            assign dm_WVALID[idx] = ap_WVALID[idx];
            assign ap_WREADY[idx] = dm_WREADY[idx];
            assign ap_BRESP[idx] = dm_BRESP[idx];
            assign ap_BVALID[idx] = dm_BVALID[idx];
            assign dm_BREADY[idx] = ap_BREADY[idx];
            assign dm_ARADDR[idx][M_AXIMM_ADDR_WIDTH-1:0] = ap_ARADDR[idx][M_AXIMM_ADDR_WIDTH-1:0];
            assign dm_ARLEN[idx] = ap_ARLEN[idx];
            assign dm_ARSIZE[idx] = ap_ARSIZE[idx];
            assign dm_ARBURST[idx] = ap_ARBURST[idx];
            assign dm_ARLOCK[idx] = ap_ARLOCK[idx];
            assign dm_ARCACHE[idx] = ap_ARCACHE[idx];
            assign dm_ARPROT[idx] = ap_ARPROT[idx];
            assign dm_ARREGION[idx] = ap_ARREGION[idx];
            assign dm_ARQOS[idx] = ap_ARQOS[idx];
            assign dm_ARVALID[idx] = ap_ARVALID[idx];
            assign ap_ARREADY[idx] = dm_ARREADY[idx];
            assign ap_RDATA[idx][M_AXIMM_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0] = dm_RDATA[idx][M_AXIMM_BIT_ARRAY[32*(idx+1)-1:32*idx]-1:0];
            assign ap_RRESP[idx] = dm_RRESP[idx];
            assign ap_RLAST[idx] = dm_RLAST[idx];
            assign ap_RVALID[idx] = dm_RVALID[idx];
            assign dm_RREADY[idx] = ap_RREADY[idx];
        end
    endgenerate
endmodule
